module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate1527(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate1528(.a(gate9inter0), .b(s_140), .O(gate9inter1));
  and2  gate1529(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate1530(.a(s_140), .O(gate9inter3));
  inv1  gate1531(.a(s_141), .O(gate9inter4));
  nand2 gate1532(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate1533(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate1534(.a(G1), .O(gate9inter7));
  inv1  gate1535(.a(G2), .O(gate9inter8));
  nand2 gate1536(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate1537(.a(s_141), .b(gate9inter3), .O(gate9inter10));
  nor2  gate1538(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate1539(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate1540(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate687(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate688(.a(gate20inter0), .b(s_20), .O(gate20inter1));
  and2  gate689(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate690(.a(s_20), .O(gate20inter3));
  inv1  gate691(.a(s_21), .O(gate20inter4));
  nand2 gate692(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate693(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate694(.a(G23), .O(gate20inter7));
  inv1  gate695(.a(G24), .O(gate20inter8));
  nand2 gate696(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate697(.a(s_21), .b(gate20inter3), .O(gate20inter10));
  nor2  gate698(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate699(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate700(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );

  xor2  gate841(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate842(.a(gate32inter0), .b(s_42), .O(gate32inter1));
  and2  gate843(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate844(.a(s_42), .O(gate32inter3));
  inv1  gate845(.a(s_43), .O(gate32inter4));
  nand2 gate846(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate847(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate848(.a(G12), .O(gate32inter7));
  inv1  gate849(.a(G16), .O(gate32inter8));
  nand2 gate850(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate851(.a(s_43), .b(gate32inter3), .O(gate32inter10));
  nor2  gate852(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate853(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate854(.a(gate32inter12), .b(gate32inter1), .O(G335));
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate1513(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate1514(.a(gate38inter0), .b(s_138), .O(gate38inter1));
  and2  gate1515(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate1516(.a(s_138), .O(gate38inter3));
  inv1  gate1517(.a(s_139), .O(gate38inter4));
  nand2 gate1518(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate1519(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate1520(.a(G27), .O(gate38inter7));
  inv1  gate1521(.a(G31), .O(gate38inter8));
  nand2 gate1522(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate1523(.a(s_139), .b(gate38inter3), .O(gate38inter10));
  nor2  gate1524(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate1525(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate1526(.a(gate38inter12), .b(gate38inter1), .O(G353));
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate771(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate772(.a(gate51inter0), .b(s_32), .O(gate51inter1));
  and2  gate773(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate774(.a(s_32), .O(gate51inter3));
  inv1  gate775(.a(s_33), .O(gate51inter4));
  nand2 gate776(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate777(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate778(.a(G11), .O(gate51inter7));
  inv1  gate779(.a(G281), .O(gate51inter8));
  nand2 gate780(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate781(.a(s_33), .b(gate51inter3), .O(gate51inter10));
  nor2  gate782(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate783(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate784(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate1401(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate1402(.a(gate54inter0), .b(s_122), .O(gate54inter1));
  and2  gate1403(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate1404(.a(s_122), .O(gate54inter3));
  inv1  gate1405(.a(s_123), .O(gate54inter4));
  nand2 gate1406(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate1407(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate1408(.a(G14), .O(gate54inter7));
  inv1  gate1409(.a(G284), .O(gate54inter8));
  nand2 gate1410(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate1411(.a(s_123), .b(gate54inter3), .O(gate54inter10));
  nor2  gate1412(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate1413(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate1414(.a(gate54inter12), .b(gate54inter1), .O(G375));

  xor2  gate925(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate926(.a(gate55inter0), .b(s_54), .O(gate55inter1));
  and2  gate927(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate928(.a(s_54), .O(gate55inter3));
  inv1  gate929(.a(s_55), .O(gate55inter4));
  nand2 gate930(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate931(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate932(.a(G15), .O(gate55inter7));
  inv1  gate933(.a(G287), .O(gate55inter8));
  nand2 gate934(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate935(.a(s_55), .b(gate55inter3), .O(gate55inter10));
  nor2  gate936(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate937(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate938(.a(gate55inter12), .b(gate55inter1), .O(G376));

  xor2  gate1247(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate1248(.a(gate56inter0), .b(s_100), .O(gate56inter1));
  and2  gate1249(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate1250(.a(s_100), .O(gate56inter3));
  inv1  gate1251(.a(s_101), .O(gate56inter4));
  nand2 gate1252(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate1253(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate1254(.a(G16), .O(gate56inter7));
  inv1  gate1255(.a(G287), .O(gate56inter8));
  nand2 gate1256(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate1257(.a(s_101), .b(gate56inter3), .O(gate56inter10));
  nor2  gate1258(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate1259(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate1260(.a(gate56inter12), .b(gate56inter1), .O(G377));

  xor2  gate1009(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate1010(.a(gate57inter0), .b(s_66), .O(gate57inter1));
  and2  gate1011(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate1012(.a(s_66), .O(gate57inter3));
  inv1  gate1013(.a(s_67), .O(gate57inter4));
  nand2 gate1014(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate1015(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate1016(.a(G17), .O(gate57inter7));
  inv1  gate1017(.a(G290), .O(gate57inter8));
  nand2 gate1018(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate1019(.a(s_67), .b(gate57inter3), .O(gate57inter10));
  nor2  gate1020(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate1021(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate1022(.a(gate57inter12), .b(gate57inter1), .O(G378));
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );

  xor2  gate1499(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate1500(.a(gate61inter0), .b(s_136), .O(gate61inter1));
  and2  gate1501(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate1502(.a(s_136), .O(gate61inter3));
  inv1  gate1503(.a(s_137), .O(gate61inter4));
  nand2 gate1504(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate1505(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate1506(.a(G21), .O(gate61inter7));
  inv1  gate1507(.a(G296), .O(gate61inter8));
  nand2 gate1508(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate1509(.a(s_137), .b(gate61inter3), .O(gate61inter10));
  nor2  gate1510(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate1511(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate1512(.a(gate61inter12), .b(gate61inter1), .O(G382));
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate967(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate968(.a(gate65inter0), .b(s_60), .O(gate65inter1));
  and2  gate969(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate970(.a(s_60), .O(gate65inter3));
  inv1  gate971(.a(s_61), .O(gate65inter4));
  nand2 gate972(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate973(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate974(.a(G25), .O(gate65inter7));
  inv1  gate975(.a(G302), .O(gate65inter8));
  nand2 gate976(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate977(.a(s_61), .b(gate65inter3), .O(gate65inter10));
  nor2  gate978(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate979(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate980(.a(gate65inter12), .b(gate65inter1), .O(G386));

  xor2  gate1555(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate1556(.a(gate66inter0), .b(s_144), .O(gate66inter1));
  and2  gate1557(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate1558(.a(s_144), .O(gate66inter3));
  inv1  gate1559(.a(s_145), .O(gate66inter4));
  nand2 gate1560(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate1561(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate1562(.a(G26), .O(gate66inter7));
  inv1  gate1563(.a(G302), .O(gate66inter8));
  nand2 gate1564(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate1565(.a(s_145), .b(gate66inter3), .O(gate66inter10));
  nor2  gate1566(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate1567(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate1568(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );

  xor2  gate939(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate940(.a(gate68inter0), .b(s_56), .O(gate68inter1));
  and2  gate941(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate942(.a(s_56), .O(gate68inter3));
  inv1  gate943(.a(s_57), .O(gate68inter4));
  nand2 gate944(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate945(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate946(.a(G28), .O(gate68inter7));
  inv1  gate947(.a(G305), .O(gate68inter8));
  nand2 gate948(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate949(.a(s_57), .b(gate68inter3), .O(gate68inter10));
  nor2  gate950(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate951(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate952(.a(gate68inter12), .b(gate68inter1), .O(G389));

  xor2  gate1219(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate1220(.a(gate69inter0), .b(s_96), .O(gate69inter1));
  and2  gate1221(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate1222(.a(s_96), .O(gate69inter3));
  inv1  gate1223(.a(s_97), .O(gate69inter4));
  nand2 gate1224(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate1225(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate1226(.a(G29), .O(gate69inter7));
  inv1  gate1227(.a(G308), .O(gate69inter8));
  nand2 gate1228(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate1229(.a(s_97), .b(gate69inter3), .O(gate69inter10));
  nor2  gate1230(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate1231(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate1232(.a(gate69inter12), .b(gate69inter1), .O(G390));
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );

  xor2  gate1317(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate1318(.a(gate73inter0), .b(s_110), .O(gate73inter1));
  and2  gate1319(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate1320(.a(s_110), .O(gate73inter3));
  inv1  gate1321(.a(s_111), .O(gate73inter4));
  nand2 gate1322(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate1323(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate1324(.a(G1), .O(gate73inter7));
  inv1  gate1325(.a(G314), .O(gate73inter8));
  nand2 gate1326(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate1327(.a(s_111), .b(gate73inter3), .O(gate73inter10));
  nor2  gate1328(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate1329(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate1330(.a(gate73inter12), .b(gate73inter1), .O(G394));
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate1541(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate1542(.a(gate85inter0), .b(s_142), .O(gate85inter1));
  and2  gate1543(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate1544(.a(s_142), .O(gate85inter3));
  inv1  gate1545(.a(s_143), .O(gate85inter4));
  nand2 gate1546(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate1547(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate1548(.a(G4), .O(gate85inter7));
  inv1  gate1549(.a(G332), .O(gate85inter8));
  nand2 gate1550(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate1551(.a(s_143), .b(gate85inter3), .O(gate85inter10));
  nor2  gate1552(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate1553(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate1554(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate869(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate870(.a(gate88inter0), .b(s_46), .O(gate88inter1));
  and2  gate871(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate872(.a(s_46), .O(gate88inter3));
  inv1  gate873(.a(s_47), .O(gate88inter4));
  nand2 gate874(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate875(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate876(.a(G16), .O(gate88inter7));
  inv1  gate877(.a(G335), .O(gate88inter8));
  nand2 gate878(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate879(.a(s_47), .b(gate88inter3), .O(gate88inter10));
  nor2  gate880(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate881(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate882(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate1261(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate1262(.a(gate90inter0), .b(s_102), .O(gate90inter1));
  and2  gate1263(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate1264(.a(s_102), .O(gate90inter3));
  inv1  gate1265(.a(s_103), .O(gate90inter4));
  nand2 gate1266(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate1267(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate1268(.a(G21), .O(gate90inter7));
  inv1  gate1269(.a(G338), .O(gate90inter8));
  nand2 gate1270(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate1271(.a(s_103), .b(gate90inter3), .O(gate90inter10));
  nor2  gate1272(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate1273(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate1274(.a(gate90inter12), .b(gate90inter1), .O(G411));
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate1569(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate1570(.a(gate95inter0), .b(s_146), .O(gate95inter1));
  and2  gate1571(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate1572(.a(s_146), .O(gate95inter3));
  inv1  gate1573(.a(s_147), .O(gate95inter4));
  nand2 gate1574(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate1575(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate1576(.a(G26), .O(gate95inter7));
  inv1  gate1577(.a(G347), .O(gate95inter8));
  nand2 gate1578(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate1579(.a(s_147), .b(gate95inter3), .O(gate95inter10));
  nor2  gate1580(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate1581(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate1582(.a(gate95inter12), .b(gate95inter1), .O(G416));

  xor2  gate715(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate716(.a(gate96inter0), .b(s_24), .O(gate96inter1));
  and2  gate717(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate718(.a(s_24), .O(gate96inter3));
  inv1  gate719(.a(s_25), .O(gate96inter4));
  nand2 gate720(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate721(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate722(.a(G30), .O(gate96inter7));
  inv1  gate723(.a(G347), .O(gate96inter8));
  nand2 gate724(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate725(.a(s_25), .b(gate96inter3), .O(gate96inter10));
  nor2  gate726(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate727(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate728(.a(gate96inter12), .b(gate96inter1), .O(G417));
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate981(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate982(.a(gate98inter0), .b(s_62), .O(gate98inter1));
  and2  gate983(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate984(.a(s_62), .O(gate98inter3));
  inv1  gate985(.a(s_63), .O(gate98inter4));
  nand2 gate986(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate987(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate988(.a(G23), .O(gate98inter7));
  inv1  gate989(.a(G350), .O(gate98inter8));
  nand2 gate990(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate991(.a(s_63), .b(gate98inter3), .O(gate98inter10));
  nor2  gate992(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate993(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate994(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate813(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate814(.a(gate102inter0), .b(s_38), .O(gate102inter1));
  and2  gate815(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate816(.a(s_38), .O(gate102inter3));
  inv1  gate817(.a(s_39), .O(gate102inter4));
  nand2 gate818(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate819(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate820(.a(G24), .O(gate102inter7));
  inv1  gate821(.a(G356), .O(gate102inter8));
  nand2 gate822(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate823(.a(s_39), .b(gate102inter3), .O(gate102inter10));
  nor2  gate824(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate825(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate826(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate645(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate646(.a(gate106inter0), .b(s_14), .O(gate106inter1));
  and2  gate647(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate648(.a(s_14), .O(gate106inter3));
  inv1  gate649(.a(s_15), .O(gate106inter4));
  nand2 gate650(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate651(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate652(.a(G364), .O(gate106inter7));
  inv1  gate653(.a(G365), .O(gate106inter8));
  nand2 gate654(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate655(.a(s_15), .b(gate106inter3), .O(gate106inter10));
  nor2  gate656(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate657(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate658(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate1205(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate1206(.a(gate109inter0), .b(s_94), .O(gate109inter1));
  and2  gate1207(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate1208(.a(s_94), .O(gate109inter3));
  inv1  gate1209(.a(s_95), .O(gate109inter4));
  nand2 gate1210(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate1211(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate1212(.a(G370), .O(gate109inter7));
  inv1  gate1213(.a(G371), .O(gate109inter8));
  nand2 gate1214(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate1215(.a(s_95), .b(gate109inter3), .O(gate109inter10));
  nor2  gate1216(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate1217(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate1218(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate1429(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate1430(.a(gate121inter0), .b(s_126), .O(gate121inter1));
  and2  gate1431(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate1432(.a(s_126), .O(gate121inter3));
  inv1  gate1433(.a(s_127), .O(gate121inter4));
  nand2 gate1434(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate1435(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate1436(.a(G394), .O(gate121inter7));
  inv1  gate1437(.a(G395), .O(gate121inter8));
  nand2 gate1438(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate1439(.a(s_127), .b(gate121inter3), .O(gate121inter10));
  nor2  gate1440(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate1441(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate1442(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate1191(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate1192(.a(gate123inter0), .b(s_92), .O(gate123inter1));
  and2  gate1193(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate1194(.a(s_92), .O(gate123inter3));
  inv1  gate1195(.a(s_93), .O(gate123inter4));
  nand2 gate1196(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate1197(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate1198(.a(G398), .O(gate123inter7));
  inv1  gate1199(.a(G399), .O(gate123inter8));
  nand2 gate1200(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate1201(.a(s_93), .b(gate123inter3), .O(gate123inter10));
  nor2  gate1202(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate1203(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate1204(.a(gate123inter12), .b(gate123inter1), .O(G480));

  xor2  gate617(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate618(.a(gate124inter0), .b(s_10), .O(gate124inter1));
  and2  gate619(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate620(.a(s_10), .O(gate124inter3));
  inv1  gate621(.a(s_11), .O(gate124inter4));
  nand2 gate622(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate623(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate624(.a(G400), .O(gate124inter7));
  inv1  gate625(.a(G401), .O(gate124inter8));
  nand2 gate626(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate627(.a(s_11), .b(gate124inter3), .O(gate124inter10));
  nor2  gate628(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate629(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate630(.a(gate124inter12), .b(gate124inter1), .O(G483));

  xor2  gate1625(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate1626(.a(gate125inter0), .b(s_154), .O(gate125inter1));
  and2  gate1627(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate1628(.a(s_154), .O(gate125inter3));
  inv1  gate1629(.a(s_155), .O(gate125inter4));
  nand2 gate1630(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate1631(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate1632(.a(G402), .O(gate125inter7));
  inv1  gate1633(.a(G403), .O(gate125inter8));
  nand2 gate1634(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate1635(.a(s_155), .b(gate125inter3), .O(gate125inter10));
  nor2  gate1636(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate1637(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate1638(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate1653(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate1654(.a(gate135inter0), .b(s_158), .O(gate135inter1));
  and2  gate1655(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate1656(.a(s_158), .O(gate135inter3));
  inv1  gate1657(.a(s_159), .O(gate135inter4));
  nand2 gate1658(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate1659(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate1660(.a(G422), .O(gate135inter7));
  inv1  gate1661(.a(G423), .O(gate135inter8));
  nand2 gate1662(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate1663(.a(s_159), .b(gate135inter3), .O(gate135inter10));
  nor2  gate1664(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate1665(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate1666(.a(gate135inter12), .b(gate135inter1), .O(G516));

  xor2  gate1177(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate1178(.a(gate136inter0), .b(s_90), .O(gate136inter1));
  and2  gate1179(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate1180(.a(s_90), .O(gate136inter3));
  inv1  gate1181(.a(s_91), .O(gate136inter4));
  nand2 gate1182(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate1183(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate1184(.a(G424), .O(gate136inter7));
  inv1  gate1185(.a(G425), .O(gate136inter8));
  nand2 gate1186(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate1187(.a(s_91), .b(gate136inter3), .O(gate136inter10));
  nor2  gate1188(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate1189(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate1190(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );

  xor2  gate953(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate954(.a(gate140inter0), .b(s_58), .O(gate140inter1));
  and2  gate955(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate956(.a(s_58), .O(gate140inter3));
  inv1  gate957(.a(s_59), .O(gate140inter4));
  nand2 gate958(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate959(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate960(.a(G444), .O(gate140inter7));
  inv1  gate961(.a(G447), .O(gate140inter8));
  nand2 gate962(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate963(.a(s_59), .b(gate140inter3), .O(gate140inter10));
  nor2  gate964(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate965(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate966(.a(gate140inter12), .b(gate140inter1), .O(G531));
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate1107(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate1108(.a(gate144inter0), .b(s_80), .O(gate144inter1));
  and2  gate1109(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate1110(.a(s_80), .O(gate144inter3));
  inv1  gate1111(.a(s_81), .O(gate144inter4));
  nand2 gate1112(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate1113(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate1114(.a(G468), .O(gate144inter7));
  inv1  gate1115(.a(G471), .O(gate144inter8));
  nand2 gate1116(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate1117(.a(s_81), .b(gate144inter3), .O(gate144inter10));
  nor2  gate1118(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate1119(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate1120(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate1289(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate1290(.a(gate157inter0), .b(s_106), .O(gate157inter1));
  and2  gate1291(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate1292(.a(s_106), .O(gate157inter3));
  inv1  gate1293(.a(s_107), .O(gate157inter4));
  nand2 gate1294(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate1295(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate1296(.a(G438), .O(gate157inter7));
  inv1  gate1297(.a(G528), .O(gate157inter8));
  nand2 gate1298(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate1299(.a(s_107), .b(gate157inter3), .O(gate157inter10));
  nor2  gate1300(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate1301(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate1302(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );

  xor2  gate1065(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate1066(.a(gate167inter0), .b(s_74), .O(gate167inter1));
  and2  gate1067(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate1068(.a(s_74), .O(gate167inter3));
  inv1  gate1069(.a(s_75), .O(gate167inter4));
  nand2 gate1070(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate1071(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate1072(.a(G468), .O(gate167inter7));
  inv1  gate1073(.a(G543), .O(gate167inter8));
  nand2 gate1074(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate1075(.a(s_75), .b(gate167inter3), .O(gate167inter10));
  nor2  gate1076(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate1077(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate1078(.a(gate167inter12), .b(gate167inter1), .O(G584));
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );

  xor2  gate1149(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate1150(.a(gate177inter0), .b(s_86), .O(gate177inter1));
  and2  gate1151(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate1152(.a(s_86), .O(gate177inter3));
  inv1  gate1153(.a(s_87), .O(gate177inter4));
  nand2 gate1154(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate1155(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate1156(.a(G498), .O(gate177inter7));
  inv1  gate1157(.a(G558), .O(gate177inter8));
  nand2 gate1158(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate1159(.a(s_87), .b(gate177inter3), .O(gate177inter10));
  nor2  gate1160(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate1161(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate1162(.a(gate177inter12), .b(gate177inter1), .O(G594));
nand2 gate178( .a(G501), .b(G558), .O(G595) );

  xor2  gate1359(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate1360(.a(gate179inter0), .b(s_116), .O(gate179inter1));
  and2  gate1361(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate1362(.a(s_116), .O(gate179inter3));
  inv1  gate1363(.a(s_117), .O(gate179inter4));
  nand2 gate1364(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate1365(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate1366(.a(G504), .O(gate179inter7));
  inv1  gate1367(.a(G561), .O(gate179inter8));
  nand2 gate1368(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate1369(.a(s_117), .b(gate179inter3), .O(gate179inter10));
  nor2  gate1370(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate1371(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate1372(.a(gate179inter12), .b(gate179inter1), .O(G596));

  xor2  gate1093(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate1094(.a(gate180inter0), .b(s_78), .O(gate180inter1));
  and2  gate1095(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate1096(.a(s_78), .O(gate180inter3));
  inv1  gate1097(.a(s_79), .O(gate180inter4));
  nand2 gate1098(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate1099(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate1100(.a(G507), .O(gate180inter7));
  inv1  gate1101(.a(G561), .O(gate180inter8));
  nand2 gate1102(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate1103(.a(s_79), .b(gate180inter3), .O(gate180inter10));
  nor2  gate1104(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate1105(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate1106(.a(gate180inter12), .b(gate180inter1), .O(G597));
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate659(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate660(.a(gate186inter0), .b(s_16), .O(gate186inter1));
  and2  gate661(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate662(.a(s_16), .O(gate186inter3));
  inv1  gate663(.a(s_17), .O(gate186inter4));
  nand2 gate664(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate665(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate666(.a(G572), .O(gate186inter7));
  inv1  gate667(.a(G573), .O(gate186inter8));
  nand2 gate668(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate669(.a(s_17), .b(gate186inter3), .O(gate186inter10));
  nor2  gate670(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate671(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate672(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate1737(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate1738(.a(gate195inter0), .b(s_170), .O(gate195inter1));
  and2  gate1739(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate1740(.a(s_170), .O(gate195inter3));
  inv1  gate1741(.a(s_171), .O(gate195inter4));
  nand2 gate1742(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate1743(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate1744(.a(G590), .O(gate195inter7));
  inv1  gate1745(.a(G591), .O(gate195inter8));
  nand2 gate1746(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate1747(.a(s_171), .b(gate195inter3), .O(gate195inter10));
  nor2  gate1748(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate1749(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate1750(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate911(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate912(.a(gate198inter0), .b(s_52), .O(gate198inter1));
  and2  gate913(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate914(.a(s_52), .O(gate198inter3));
  inv1  gate915(.a(s_53), .O(gate198inter4));
  nand2 gate916(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate917(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate918(.a(G596), .O(gate198inter7));
  inv1  gate919(.a(G597), .O(gate198inter8));
  nand2 gate920(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate921(.a(s_53), .b(gate198inter3), .O(gate198inter10));
  nor2  gate922(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate923(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate924(.a(gate198inter12), .b(gate198inter1), .O(G657));

  xor2  gate575(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate576(.a(gate199inter0), .b(s_4), .O(gate199inter1));
  and2  gate577(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate578(.a(s_4), .O(gate199inter3));
  inv1  gate579(.a(s_5), .O(gate199inter4));
  nand2 gate580(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate581(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate582(.a(G598), .O(gate199inter7));
  inv1  gate583(.a(G599), .O(gate199inter8));
  nand2 gate584(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate585(.a(s_5), .b(gate199inter3), .O(gate199inter10));
  nor2  gate586(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate587(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate588(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );

  xor2  gate1443(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate1444(.a(gate204inter0), .b(s_128), .O(gate204inter1));
  and2  gate1445(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate1446(.a(s_128), .O(gate204inter3));
  inv1  gate1447(.a(s_129), .O(gate204inter4));
  nand2 gate1448(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate1449(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate1450(.a(G607), .O(gate204inter7));
  inv1  gate1451(.a(G617), .O(gate204inter8));
  nand2 gate1452(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate1453(.a(s_129), .b(gate204inter3), .O(gate204inter10));
  nor2  gate1454(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate1455(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate1456(.a(gate204inter12), .b(gate204inter1), .O(G675));
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate1639(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate1640(.a(gate214inter0), .b(s_156), .O(gate214inter1));
  and2  gate1641(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate1642(.a(s_156), .O(gate214inter3));
  inv1  gate1643(.a(s_157), .O(gate214inter4));
  nand2 gate1644(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate1645(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate1646(.a(G612), .O(gate214inter7));
  inv1  gate1647(.a(G672), .O(gate214inter8));
  nand2 gate1648(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate1649(.a(s_157), .b(gate214inter3), .O(gate214inter10));
  nor2  gate1650(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate1651(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate1652(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate547(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate548(.a(gate226inter0), .b(s_0), .O(gate226inter1));
  and2  gate549(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate550(.a(s_0), .O(gate226inter3));
  inv1  gate551(.a(s_1), .O(gate226inter4));
  nand2 gate552(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate553(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate554(.a(G692), .O(gate226inter7));
  inv1  gate555(.a(G693), .O(gate226inter8));
  nand2 gate556(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate557(.a(s_1), .b(gate226inter3), .O(gate226inter10));
  nor2  gate558(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate559(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate560(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );

  xor2  gate1597(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate1598(.a(gate230inter0), .b(s_150), .O(gate230inter1));
  and2  gate1599(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate1600(.a(s_150), .O(gate230inter3));
  inv1  gate1601(.a(s_151), .O(gate230inter4));
  nand2 gate1602(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate1603(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate1604(.a(G700), .O(gate230inter7));
  inv1  gate1605(.a(G701), .O(gate230inter8));
  nand2 gate1606(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate1607(.a(s_151), .b(gate230inter3), .O(gate230inter10));
  nor2  gate1608(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate1609(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate1610(.a(gate230inter12), .b(gate230inter1), .O(G721));
nand2 gate231( .a(G702), .b(G703), .O(G724) );

  xor2  gate785(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate786(.a(gate232inter0), .b(s_34), .O(gate232inter1));
  and2  gate787(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate788(.a(s_34), .O(gate232inter3));
  inv1  gate789(.a(s_35), .O(gate232inter4));
  nand2 gate790(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate791(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate792(.a(G704), .O(gate232inter7));
  inv1  gate793(.a(G705), .O(gate232inter8));
  nand2 gate794(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate795(.a(s_35), .b(gate232inter3), .O(gate232inter10));
  nor2  gate796(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate797(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate798(.a(gate232inter12), .b(gate232inter1), .O(G727));
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );

  xor2  gate1471(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate1472(.a(gate235inter0), .b(s_132), .O(gate235inter1));
  and2  gate1473(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate1474(.a(s_132), .O(gate235inter3));
  inv1  gate1475(.a(s_133), .O(gate235inter4));
  nand2 gate1476(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate1477(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate1478(.a(G248), .O(gate235inter7));
  inv1  gate1479(.a(G724), .O(gate235inter8));
  nand2 gate1480(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate1481(.a(s_133), .b(gate235inter3), .O(gate235inter10));
  nor2  gate1482(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate1483(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate1484(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate603(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate604(.a(gate240inter0), .b(s_8), .O(gate240inter1));
  and2  gate605(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate606(.a(s_8), .O(gate240inter3));
  inv1  gate607(.a(s_9), .O(gate240inter4));
  nand2 gate608(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate609(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate610(.a(G263), .O(gate240inter7));
  inv1  gate611(.a(G715), .O(gate240inter8));
  nand2 gate612(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate613(.a(s_9), .b(gate240inter3), .O(gate240inter10));
  nor2  gate614(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate615(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate616(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );

  xor2  gate1345(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate1346(.a(gate242inter0), .b(s_114), .O(gate242inter1));
  and2  gate1347(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate1348(.a(s_114), .O(gate242inter3));
  inv1  gate1349(.a(s_115), .O(gate242inter4));
  nand2 gate1350(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate1351(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate1352(.a(G718), .O(gate242inter7));
  inv1  gate1353(.a(G730), .O(gate242inter8));
  nand2 gate1354(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate1355(.a(s_115), .b(gate242inter3), .O(gate242inter10));
  nor2  gate1356(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate1357(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate1358(.a(gate242inter12), .b(gate242inter1), .O(G755));
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate1373(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate1374(.a(gate249inter0), .b(s_118), .O(gate249inter1));
  and2  gate1375(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate1376(.a(s_118), .O(gate249inter3));
  inv1  gate1377(.a(s_119), .O(gate249inter4));
  nand2 gate1378(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate1379(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate1380(.a(G254), .O(gate249inter7));
  inv1  gate1381(.a(G742), .O(gate249inter8));
  nand2 gate1382(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate1383(.a(s_119), .b(gate249inter3), .O(gate249inter10));
  nor2  gate1384(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate1385(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate1386(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );

  xor2  gate631(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate632(.a(gate254inter0), .b(s_12), .O(gate254inter1));
  and2  gate633(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate634(.a(s_12), .O(gate254inter3));
  inv1  gate635(.a(s_13), .O(gate254inter4));
  nand2 gate636(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate637(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate638(.a(G712), .O(gate254inter7));
  inv1  gate639(.a(G748), .O(gate254inter8));
  nand2 gate640(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate641(.a(s_13), .b(gate254inter3), .O(gate254inter10));
  nor2  gate642(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate643(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate644(.a(gate254inter12), .b(gate254inter1), .O(G767));
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate1583(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate1584(.a(gate267inter0), .b(s_148), .O(gate267inter1));
  and2  gate1585(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate1586(.a(s_148), .O(gate267inter3));
  inv1  gate1587(.a(s_149), .O(gate267inter4));
  nand2 gate1588(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate1589(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate1590(.a(G648), .O(gate267inter7));
  inv1  gate1591(.a(G776), .O(gate267inter8));
  nand2 gate1592(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate1593(.a(s_149), .b(gate267inter3), .O(gate267inter10));
  nor2  gate1594(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate1595(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate1596(.a(gate267inter12), .b(gate267inter1), .O(G800));

  xor2  gate1485(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate1486(.a(gate268inter0), .b(s_134), .O(gate268inter1));
  and2  gate1487(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate1488(.a(s_134), .O(gate268inter3));
  inv1  gate1489(.a(s_135), .O(gate268inter4));
  nand2 gate1490(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1491(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1492(.a(G651), .O(gate268inter7));
  inv1  gate1493(.a(G779), .O(gate268inter8));
  nand2 gate1494(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1495(.a(s_135), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1496(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1497(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1498(.a(gate268inter12), .b(gate268inter1), .O(G803));

  xor2  gate1611(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate1612(.a(gate269inter0), .b(s_152), .O(gate269inter1));
  and2  gate1613(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate1614(.a(s_152), .O(gate269inter3));
  inv1  gate1615(.a(s_153), .O(gate269inter4));
  nand2 gate1616(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate1617(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate1618(.a(G654), .O(gate269inter7));
  inv1  gate1619(.a(G782), .O(gate269inter8));
  nand2 gate1620(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate1621(.a(s_153), .b(gate269inter3), .O(gate269inter10));
  nor2  gate1622(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate1623(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate1624(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );

  xor2  gate1163(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate1164(.a(gate273inter0), .b(s_88), .O(gate273inter1));
  and2  gate1165(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate1166(.a(s_88), .O(gate273inter3));
  inv1  gate1167(.a(s_89), .O(gate273inter4));
  nand2 gate1168(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate1169(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate1170(.a(G642), .O(gate273inter7));
  inv1  gate1171(.a(G794), .O(gate273inter8));
  nand2 gate1172(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate1173(.a(s_89), .b(gate273inter3), .O(gate273inter10));
  nor2  gate1174(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate1175(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate1176(.a(gate273inter12), .b(gate273inter1), .O(G818));
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate1051(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate1052(.a(gate276inter0), .b(s_72), .O(gate276inter1));
  and2  gate1053(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate1054(.a(s_72), .O(gate276inter3));
  inv1  gate1055(.a(s_73), .O(gate276inter4));
  nand2 gate1056(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate1057(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate1058(.a(G773), .O(gate276inter7));
  inv1  gate1059(.a(G797), .O(gate276inter8));
  nand2 gate1060(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate1061(.a(s_73), .b(gate276inter3), .O(gate276inter10));
  nor2  gate1062(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate1063(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate1064(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate1387(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate1388(.a(gate278inter0), .b(s_120), .O(gate278inter1));
  and2  gate1389(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate1390(.a(s_120), .O(gate278inter3));
  inv1  gate1391(.a(s_121), .O(gate278inter4));
  nand2 gate1392(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate1393(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate1394(.a(G776), .O(gate278inter7));
  inv1  gate1395(.a(G800), .O(gate278inter8));
  nand2 gate1396(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate1397(.a(s_121), .b(gate278inter3), .O(gate278inter10));
  nor2  gate1398(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate1399(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate1400(.a(gate278inter12), .b(gate278inter1), .O(G823));

  xor2  gate729(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate730(.a(gate279inter0), .b(s_26), .O(gate279inter1));
  and2  gate731(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate732(.a(s_26), .O(gate279inter3));
  inv1  gate733(.a(s_27), .O(gate279inter4));
  nand2 gate734(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate735(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate736(.a(G651), .O(gate279inter7));
  inv1  gate737(.a(G803), .O(gate279inter8));
  nand2 gate738(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate739(.a(s_27), .b(gate279inter3), .O(gate279inter10));
  nor2  gate740(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate741(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate742(.a(gate279inter12), .b(gate279inter1), .O(G824));

  xor2  gate1135(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate1136(.a(gate280inter0), .b(s_84), .O(gate280inter1));
  and2  gate1137(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate1138(.a(s_84), .O(gate280inter3));
  inv1  gate1139(.a(s_85), .O(gate280inter4));
  nand2 gate1140(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate1141(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate1142(.a(G779), .O(gate280inter7));
  inv1  gate1143(.a(G803), .O(gate280inter8));
  nand2 gate1144(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate1145(.a(s_85), .b(gate280inter3), .O(gate280inter10));
  nor2  gate1146(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate1147(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate1148(.a(gate280inter12), .b(gate280inter1), .O(G825));

  xor2  gate799(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate800(.a(gate281inter0), .b(s_36), .O(gate281inter1));
  and2  gate801(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate802(.a(s_36), .O(gate281inter3));
  inv1  gate803(.a(s_37), .O(gate281inter4));
  nand2 gate804(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate805(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate806(.a(G654), .O(gate281inter7));
  inv1  gate807(.a(G806), .O(gate281inter8));
  nand2 gate808(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate809(.a(s_37), .b(gate281inter3), .O(gate281inter10));
  nor2  gate810(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate811(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate812(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate855(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate856(.a(gate288inter0), .b(s_44), .O(gate288inter1));
  and2  gate857(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate858(.a(s_44), .O(gate288inter3));
  inv1  gate859(.a(s_45), .O(gate288inter4));
  nand2 gate860(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate861(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate862(.a(G791), .O(gate288inter7));
  inv1  gate863(.a(G815), .O(gate288inter8));
  nand2 gate864(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate865(.a(s_45), .b(gate288inter3), .O(gate288inter10));
  nor2  gate866(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate867(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate868(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate561(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate562(.a(gate291inter0), .b(s_2), .O(gate291inter1));
  and2  gate563(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate564(.a(s_2), .O(gate291inter3));
  inv1  gate565(.a(s_3), .O(gate291inter4));
  nand2 gate566(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate567(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate568(.a(G822), .O(gate291inter7));
  inv1  gate569(.a(G823), .O(gate291inter8));
  nand2 gate570(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate571(.a(s_3), .b(gate291inter3), .O(gate291inter10));
  nor2  gate572(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate573(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate574(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate1457(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate1458(.a(gate293inter0), .b(s_130), .O(gate293inter1));
  and2  gate1459(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate1460(.a(s_130), .O(gate293inter3));
  inv1  gate1461(.a(s_131), .O(gate293inter4));
  nand2 gate1462(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate1463(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate1464(.a(G828), .O(gate293inter7));
  inv1  gate1465(.a(G829), .O(gate293inter8));
  nand2 gate1466(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate1467(.a(s_131), .b(gate293inter3), .O(gate293inter10));
  nor2  gate1468(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate1469(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate1470(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate883(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate884(.a(gate394inter0), .b(s_48), .O(gate394inter1));
  and2  gate885(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate886(.a(s_48), .O(gate394inter3));
  inv1  gate887(.a(s_49), .O(gate394inter4));
  nand2 gate888(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate889(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate890(.a(G8), .O(gate394inter7));
  inv1  gate891(.a(G1057), .O(gate394inter8));
  nand2 gate892(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate893(.a(s_49), .b(gate394inter3), .O(gate394inter10));
  nor2  gate894(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate895(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate896(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate673(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate674(.a(gate397inter0), .b(s_18), .O(gate397inter1));
  and2  gate675(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate676(.a(s_18), .O(gate397inter3));
  inv1  gate677(.a(s_19), .O(gate397inter4));
  nand2 gate678(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate679(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate680(.a(G11), .O(gate397inter7));
  inv1  gate681(.a(G1066), .O(gate397inter8));
  nand2 gate682(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate683(.a(s_19), .b(gate397inter3), .O(gate397inter10));
  nor2  gate684(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate685(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate686(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate1275(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate1276(.a(gate411inter0), .b(s_104), .O(gate411inter1));
  and2  gate1277(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate1278(.a(s_104), .O(gate411inter3));
  inv1  gate1279(.a(s_105), .O(gate411inter4));
  nand2 gate1280(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate1281(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate1282(.a(G25), .O(gate411inter7));
  inv1  gate1283(.a(G1108), .O(gate411inter8));
  nand2 gate1284(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate1285(.a(s_105), .b(gate411inter3), .O(gate411inter10));
  nor2  gate1286(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate1287(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate1288(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate1681(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate1682(.a(gate415inter0), .b(s_162), .O(gate415inter1));
  and2  gate1683(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate1684(.a(s_162), .O(gate415inter3));
  inv1  gate1685(.a(s_163), .O(gate415inter4));
  nand2 gate1686(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate1687(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate1688(.a(G29), .O(gate415inter7));
  inv1  gate1689(.a(G1120), .O(gate415inter8));
  nand2 gate1690(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate1691(.a(s_163), .b(gate415inter3), .O(gate415inter10));
  nor2  gate1692(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate1693(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate1694(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate1079(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate1080(.a(gate435inter0), .b(s_76), .O(gate435inter1));
  and2  gate1081(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate1082(.a(s_76), .O(gate435inter3));
  inv1  gate1083(.a(s_77), .O(gate435inter4));
  nand2 gate1084(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate1085(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate1086(.a(G9), .O(gate435inter7));
  inv1  gate1087(.a(G1156), .O(gate435inter8));
  nand2 gate1088(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate1089(.a(s_77), .b(gate435inter3), .O(gate435inter10));
  nor2  gate1090(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate1091(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate1092(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );

  xor2  gate995(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate996(.a(gate440inter0), .b(s_64), .O(gate440inter1));
  and2  gate997(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate998(.a(s_64), .O(gate440inter3));
  inv1  gate999(.a(s_65), .O(gate440inter4));
  nand2 gate1000(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate1001(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate1002(.a(G1066), .O(gate440inter7));
  inv1  gate1003(.a(G1162), .O(gate440inter8));
  nand2 gate1004(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate1005(.a(s_65), .b(gate440inter3), .O(gate440inter10));
  nor2  gate1006(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate1007(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate1008(.a(gate440inter12), .b(gate440inter1), .O(G1249));
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate827(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate828(.a(gate445inter0), .b(s_40), .O(gate445inter1));
  and2  gate829(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate830(.a(s_40), .O(gate445inter3));
  inv1  gate831(.a(s_41), .O(gate445inter4));
  nand2 gate832(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate833(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate834(.a(G14), .O(gate445inter7));
  inv1  gate835(.a(G1171), .O(gate445inter8));
  nand2 gate836(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate837(.a(s_41), .b(gate445inter3), .O(gate445inter10));
  nor2  gate838(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate839(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate840(.a(gate445inter12), .b(gate445inter1), .O(G1254));

  xor2  gate1037(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate1038(.a(gate446inter0), .b(s_70), .O(gate446inter1));
  and2  gate1039(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate1040(.a(s_70), .O(gate446inter3));
  inv1  gate1041(.a(s_71), .O(gate446inter4));
  nand2 gate1042(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate1043(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate1044(.a(G1075), .O(gate446inter7));
  inv1  gate1045(.a(G1171), .O(gate446inter8));
  nand2 gate1046(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate1047(.a(s_71), .b(gate446inter3), .O(gate446inter10));
  nor2  gate1048(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate1049(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate1050(.a(gate446inter12), .b(gate446inter1), .O(G1255));

  xor2  gate1695(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate1696(.a(gate447inter0), .b(s_164), .O(gate447inter1));
  and2  gate1697(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate1698(.a(s_164), .O(gate447inter3));
  inv1  gate1699(.a(s_165), .O(gate447inter4));
  nand2 gate1700(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate1701(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate1702(.a(G15), .O(gate447inter7));
  inv1  gate1703(.a(G1174), .O(gate447inter8));
  nand2 gate1704(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate1705(.a(s_165), .b(gate447inter3), .O(gate447inter10));
  nor2  gate1706(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate1707(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate1708(.a(gate447inter12), .b(gate447inter1), .O(G1256));
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );

  xor2  gate1121(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate1122(.a(gate449inter0), .b(s_82), .O(gate449inter1));
  and2  gate1123(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate1124(.a(s_82), .O(gate449inter3));
  inv1  gate1125(.a(s_83), .O(gate449inter4));
  nand2 gate1126(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate1127(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate1128(.a(G16), .O(gate449inter7));
  inv1  gate1129(.a(G1177), .O(gate449inter8));
  nand2 gate1130(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate1131(.a(s_83), .b(gate449inter3), .O(gate449inter10));
  nor2  gate1132(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate1133(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate1134(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate1709(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate1710(.a(gate457inter0), .b(s_166), .O(gate457inter1));
  and2  gate1711(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate1712(.a(s_166), .O(gate457inter3));
  inv1  gate1713(.a(s_167), .O(gate457inter4));
  nand2 gate1714(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate1715(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate1716(.a(G20), .O(gate457inter7));
  inv1  gate1717(.a(G1189), .O(gate457inter8));
  nand2 gate1718(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate1719(.a(s_167), .b(gate457inter3), .O(gate457inter10));
  nor2  gate1720(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate1721(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate1722(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );

  xor2  gate1415(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate1416(.a(gate469inter0), .b(s_124), .O(gate469inter1));
  and2  gate1417(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate1418(.a(s_124), .O(gate469inter3));
  inv1  gate1419(.a(s_125), .O(gate469inter4));
  nand2 gate1420(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate1421(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate1422(.a(G26), .O(gate469inter7));
  inv1  gate1423(.a(G1207), .O(gate469inter8));
  nand2 gate1424(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate1425(.a(s_125), .b(gate469inter3), .O(gate469inter10));
  nor2  gate1426(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate1427(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate1428(.a(gate469inter12), .b(gate469inter1), .O(G1278));
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );

  xor2  gate1667(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate1668(.a(gate473inter0), .b(s_160), .O(gate473inter1));
  and2  gate1669(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate1670(.a(s_160), .O(gate473inter3));
  inv1  gate1671(.a(s_161), .O(gate473inter4));
  nand2 gate1672(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate1673(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate1674(.a(G28), .O(gate473inter7));
  inv1  gate1675(.a(G1213), .O(gate473inter8));
  nand2 gate1676(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate1677(.a(s_161), .b(gate473inter3), .O(gate473inter10));
  nor2  gate1678(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate1679(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate1680(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate757(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate758(.a(gate476inter0), .b(s_30), .O(gate476inter1));
  and2  gate759(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate760(.a(s_30), .O(gate476inter3));
  inv1  gate761(.a(s_31), .O(gate476inter4));
  nand2 gate762(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate763(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate764(.a(G1120), .O(gate476inter7));
  inv1  gate765(.a(G1216), .O(gate476inter8));
  nand2 gate766(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate767(.a(s_31), .b(gate476inter3), .O(gate476inter10));
  nor2  gate768(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate769(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate770(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );

  xor2  gate589(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate590(.a(gate479inter0), .b(s_6), .O(gate479inter1));
  and2  gate591(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate592(.a(s_6), .O(gate479inter3));
  inv1  gate593(.a(s_7), .O(gate479inter4));
  nand2 gate594(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate595(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate596(.a(G31), .O(gate479inter7));
  inv1  gate597(.a(G1222), .O(gate479inter8));
  nand2 gate598(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate599(.a(s_7), .b(gate479inter3), .O(gate479inter10));
  nor2  gate600(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate601(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate602(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate743(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate744(.a(gate485inter0), .b(s_28), .O(gate485inter1));
  and2  gate745(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate746(.a(s_28), .O(gate485inter3));
  inv1  gate747(.a(s_29), .O(gate485inter4));
  nand2 gate748(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate749(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate750(.a(G1232), .O(gate485inter7));
  inv1  gate751(.a(G1233), .O(gate485inter8));
  nand2 gate752(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate753(.a(s_29), .b(gate485inter3), .O(gate485inter10));
  nor2  gate754(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate755(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate756(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate897(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate898(.a(gate492inter0), .b(s_50), .O(gate492inter1));
  and2  gate899(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate900(.a(s_50), .O(gate492inter3));
  inv1  gate901(.a(s_51), .O(gate492inter4));
  nand2 gate902(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate903(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate904(.a(G1246), .O(gate492inter7));
  inv1  gate905(.a(G1247), .O(gate492inter8));
  nand2 gate906(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate907(.a(s_51), .b(gate492inter3), .O(gate492inter10));
  nor2  gate908(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate909(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate910(.a(gate492inter12), .b(gate492inter1), .O(G1301));
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate1023(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1024(.a(gate494inter0), .b(s_68), .O(gate494inter1));
  and2  gate1025(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1026(.a(s_68), .O(gate494inter3));
  inv1  gate1027(.a(s_69), .O(gate494inter4));
  nand2 gate1028(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1029(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1030(.a(G1250), .O(gate494inter7));
  inv1  gate1031(.a(G1251), .O(gate494inter8));
  nand2 gate1032(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1033(.a(s_69), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1034(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1035(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1036(.a(gate494inter12), .b(gate494inter1), .O(G1303));

  xor2  gate701(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate702(.a(gate495inter0), .b(s_22), .O(gate495inter1));
  and2  gate703(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate704(.a(s_22), .O(gate495inter3));
  inv1  gate705(.a(s_23), .O(gate495inter4));
  nand2 gate706(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate707(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate708(.a(G1252), .O(gate495inter7));
  inv1  gate709(.a(G1253), .O(gate495inter8));
  nand2 gate710(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate711(.a(s_23), .b(gate495inter3), .O(gate495inter10));
  nor2  gate712(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate713(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate714(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate1723(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate1724(.a(gate500inter0), .b(s_168), .O(gate500inter1));
  and2  gate1725(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate1726(.a(s_168), .O(gate500inter3));
  inv1  gate1727(.a(s_169), .O(gate500inter4));
  nand2 gate1728(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate1729(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate1730(.a(G1262), .O(gate500inter7));
  inv1  gate1731(.a(G1263), .O(gate500inter8));
  nand2 gate1732(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate1733(.a(s_169), .b(gate500inter3), .O(gate500inter10));
  nor2  gate1734(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate1735(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate1736(.a(gate500inter12), .b(gate500inter1), .O(G1309));

  xor2  gate1331(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate1332(.a(gate501inter0), .b(s_112), .O(gate501inter1));
  and2  gate1333(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate1334(.a(s_112), .O(gate501inter3));
  inv1  gate1335(.a(s_113), .O(gate501inter4));
  nand2 gate1336(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1337(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1338(.a(G1264), .O(gate501inter7));
  inv1  gate1339(.a(G1265), .O(gate501inter8));
  nand2 gate1340(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1341(.a(s_113), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1342(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1343(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1344(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate1233(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate1234(.a(gate503inter0), .b(s_98), .O(gate503inter1));
  and2  gate1235(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate1236(.a(s_98), .O(gate503inter3));
  inv1  gate1237(.a(s_99), .O(gate503inter4));
  nand2 gate1238(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate1239(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate1240(.a(G1268), .O(gate503inter7));
  inv1  gate1241(.a(G1269), .O(gate503inter8));
  nand2 gate1242(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate1243(.a(s_99), .b(gate503inter3), .O(gate503inter10));
  nor2  gate1244(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate1245(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate1246(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );

  xor2  gate1303(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate1304(.a(gate507inter0), .b(s_108), .O(gate507inter1));
  and2  gate1305(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate1306(.a(s_108), .O(gate507inter3));
  inv1  gate1307(.a(s_109), .O(gate507inter4));
  nand2 gate1308(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate1309(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate1310(.a(G1276), .O(gate507inter7));
  inv1  gate1311(.a(G1277), .O(gate507inter8));
  nand2 gate1312(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate1313(.a(s_109), .b(gate507inter3), .O(gate507inter10));
  nor2  gate1314(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate1315(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate1316(.a(gate507inter12), .b(gate507inter1), .O(G1316));
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule