module c2670 (N1,N2,N3,N4,N5,N6,N7,N8,N11,N14,
              N15,N16,N19,N20,N21,N22,N23,N24,N25,N26,
              N27,N28,N29,N32,N33,N34,N35,N36,N37,N40,
              N43,N44,N47,N48,N49,N50,N51,N52,N53,N54,
              N55,N56,N57,N60,N61,N62,N63,N64,N65,N66,
              N67,N68,N69,N72,N73,N74,N75,N76,N77,N78,
              N79,N80,N81,N82,N85,N86,N87,N88,N89,N90,
              N91,N92,N93,N94,N95,N96,N99,N100,N101,N102,
              N103,N104,N105,N106,N107,N108,N111,N112,N113,N114,
              N115,N116,N117,N118,N119,N120,N123,N124,N125,N126,
              N127,N128,N129,N130,N131,N132,N135,N136,N137,N138,
              N139,N140,N141,N142,N219,N224,N227,N230,N231,N234,
              N237,N241,N246,N253,N256,N259,N262,N263,N266,N269,
              N272,N275,N278,N281,N284,N287,N290,N294,N297,N301,
              N305,N309,N313,N316,N319,N322,N325,N328,N331,N334,
              N337,N340,N343,N346,N349,N352,N355,N143_I,N144_I,N145_I,
              N146_I,N147_I,N148_I,N149_I,N150_I,N151_I,N152_I,N153_I,N154_I,N155_I,
              N156_I,N157_I,N158_I,N159_I,N160_I,N161_I,N162_I,N163_I,N164_I,N165_I,
              N166_I,N167_I,N168_I,N169_I,N170_I,N171_I,N172_I,N173_I,N174_I,N175_I,
              N176_I,N177_I,N178_I,N179_I,N180_I,N181_I,N182_I,N183_I,N184_I,N185_I,
              N186_I,N187_I,N188_I,N189_I,N190_I,N191_I,N192_I,N193_I,N194_I,N195_I,
              N196_I,N197_I,N198_I,N199_I,N200_I,N201_I,N202_I,N203_I,N204_I,N205_I,
              N206_I,N207_I,N208_I,N209_I,N210_I,N211_I,N212_I,N213_I,N214_I,N215_I,
              N216_I,N217_I,N218_I,N398,N400,N401,N419,N420,N456,N457,
              N458,N487,N488,N489,N490,N491,N492,N493,N494,N792,
              N799,N805,N1026,N1028,N1029,N1269,N1277,N1448,N1726,N1816,
              N1817,N1818,N1819,N1820,N1821,N1969,N1970,N1971,N2010,N2012,
              N2014,N2016,N2018,N2020,N2022,N2387,N2388,N2389,N2390,N2496,
              N2643,N2644,N2891,N2925,N2970,N2971,N3038,N3079,N3546,N3671,
              N3803,N3804,N3809,N3851,N3875,N3881,N3882,N143_O,N144_O,N145_O,
              N146_O,N147_O,N148_O,N149_O,N150_O,N151_O,N152_O,N153_O,N154_O,N155_O,
              N156_O,N157_O,N158_O,N159_O,N160_O,N161_O,N162_O,N163_O,N164_O,N165_O,
              N166_O,N167_O,N168_O,N169_O,N170_O,N171_O,N172_O,N173_O,N174_O,N175_O,
              N176_O,N177_O,N178_O,N179_O,N180_O,N181_O,N182_O,N183_O,N184_O,N185_O,
              N186_O,N187_O,N188_O,N189_O,N190_O,N191_O,N192_O,N193_O,N194_O,N195_O,
              N196_O,N197_O,N198_O,N199_O,N200_O,N201_O,N202_O,N203_O,N204_O,N205_O,
              N206_O,N207_O,N208_O,N209_O,N210_O,N211_O,N212_O,N213_O,N214_O,N215_O,
              N216_O,N217_O,N218_O);
input N1,N2,N3,N4,N5,N6,N7,N8,N11,N14,
      N15,N16,N19,N20,N21,N22,N23,N24,N25,N26,
      N27,N28,N29,N32,N33,N34,N35,N36,N37,N40,
      N43,N44,N47,N48,N49,N50,N51,N52,N53,N54,
      N55,N56,N57,N60,N61,N62,N63,N64,N65,N66,
      N67,N68,N69,N72,N73,N74,N75,N76,N77,N78,
      N79,N80,N81,N82,N85,N86,N87,N88,N89,N90,
      N91,N92,N93,N94,N95,N96,N99,N100,N101,N102,
      N103,N104,N105,N106,N107,N108,N111,N112,N113,N114,
      N115,N116,N117,N118,N119,N120,N123,N124,N125,N126,
      N127,N128,N129,N130,N131,N132,N135,N136,N137,N138,
      N139,N140,N141,N142,N219,N224,N227,N230,N231,N234,
      N237,N241,N246,N253,N256,N259,N262,N263,N266,N269,
      N272,N275,N278,N281,N284,N287,N290,N294,N297,N301,
      N305,N309,N313,N316,N319,N322,N325,N328,N331,N334,
      N337,N340,N343,N346,N349,N352,N355,N143_I,N144_I,N145_I,
      N146_I,N147_I,N148_I,N149_I,N150_I,N151_I,N152_I,N153_I,N154_I,N155_I,
      N156_I,N157_I,N158_I,N159_I,N160_I,N161_I,N162_I,N163_I,N164_I,N165_I,
      N166_I,N167_I,N168_I,N169_I,N170_I,N171_I,N172_I,N173_I,N174_I,N175_I,
      N176_I,N177_I,N178_I,N179_I,N180_I,N181_I,N182_I,N183_I,N184_I,N185_I,
      N186_I,N187_I,N188_I,N189_I,N190_I,N191_I,N192_I,N193_I,N194_I,N195_I,
      N196_I,N197_I,N198_I,N199_I,N200_I,N201_I,N202_I,N203_I,N204_I,N205_I,
      N206_I,N207_I,N208_I,N209_I,N210_I,N211_I,N212_I,N213_I,N214_I,N215_I,
      N216_I,N217_I,N218_I;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251;
output N398,N400,N401,N419,N420,N456,N457,N458,N487,N488,
       N489,N490,N491,N492,N493,N494,N792,N799,N805,N1026,
       N1028,N1029,N1269,N1277,N1448,N1726,N1816,N1817,N1818,N1819,
       N1820,N1821,N1969,N1970,N1971,N2010,N2012,N2014,N2016,N2018,
       N2020,N2022,N2387,N2388,N2389,N2390,N2496,N2643,N2644,N2891,
       N2925,N2970,N2971,N3038,N3079,N3546,N3671,N3803,N3804,N3809,
       N3851,N3875,N3881,N3882,N143_O,N144_O,N145_O,N146_O,N147_O,N148_O,
       N149_O,N150_O,N151_O,N152_O,N153_O,N154_O,N155_O,N156_O,N157_O,N158_O,
       N159_O,N160_O,N161_O,N162_O,N163_O,N164_O,N165_O,N166_O,N167_O,N168_O,
       N169_O,N170_O,N171_O,N172_O,N173_O,N174_O,N175_O,N176_O,N177_O,N178_O,
       N179_O,N180_O,N181_O,N182_O,N183_O,N184_O,N185_O,N186_O,N187_O,N188_O,
       N189_O,N190_O,N191_O,N192_O,N193_O,N194_O,N195_O,N196_O,N197_O,N198_O,
       N199_O,N200_O,N201_O,N202_O,N203_O,N204_O,N205_O,N206_O,N207_O,N208_O,
       N209_O,N210_O,N211_O,N212_O,N213_O,N214_O,N215_O,N216_O,N217_O,N218_O;
wire N405,N408,N425,N485,N486,N495,N496,N499,N500,N503,
     N506,N509,N521,N533,N537,N543,N544,N547,N550,N562,
     N574,N578,N582,N594,N606,N607,N608,N609,N610,N611,
     N612,N613,N625,N637,N643,N650,N651,N655,N659,N663,
     N667,N671,N675,N679,N683,N687,N693,N699,N705,N711,
     N715,N719,N723,N727,N730,N733,N734,N735,N738,N741,
     N744,N747,N750,N753,N756,N759,N762,N765,N768,N771,
     N774,N777,N780,N783,N786,N800,N900,N901,N902,N903,
     N904,N905,N998,N999,N1027,N1032,N1033,N1034,N1037,N1042,
     N1053,N1064,N1065,N1066,N1067,N1068,N1069,N1070,N1075,N1086,
     N1097,N1098,N1099,N1100,N1101,N1102,N1113,N1124,N1125,N1126,
     N1127,N1128,N1129,N1133,N1137,N1140,N1141,N1142,N1143,N1144,
     N1145,N1146,N1157,N1168,N1169,N1170,N1171,N1172,N1173,N1178,
     N1184,N1185,N1186,N1187,N1188,N1189,N1190,N1195,N1200,N1205,
     N1210,N1211,N1212,N1213,N1214,N1215,N1216,N1219,N1222,N1225,
     N1228,N1231,N1234,N1237,N1240,N1243,N1246,N1249,N1250,N1251,
     N1254,N1257,N1260,N1263,N1266,N1275,N1276,N1302,N1351,N1352,
     N1353,N1354,N1355,N1395,N1396,N1397,N1398,N1399,N1422,N1423,
     N1424,N1425,N1426,N1427,N1440,N1441,N1449,N1450,N1451,N1452,
     N1453,N1454,N1455,N1456,N1457,N1458,N1459,N1460,N1461,N1462,
     N1463,N1464,N1465,N1466,N1467,N1468,N1469,N1470,N1471,N1472,
     N1473,N1474,N1475,N1476,N1477,N1478,N1479,N1480,N1481,N1482,
     N1483,N1484,N1485,N1486,N1487,N1488,N1489,N1490,N1491,N1492,
     N1493,N1494,N1495,N1496,N1499,N1502,N1506,N1510,N1513,N1516,
     N1519,N1520,N1521,N1522,N1523,N1524,N1525,N1526,N1527,N1528,
     N1529,N1530,N1531,N1532,N1533,N1534,N1535,N1536,N1537,N1538,
     N1539,N1540,N1541,N1542,N1543,N1544,N1545,N1546,N1547,N1548,
     N1549,N1550,N1551,N1552,N1553,N1557,N1561,N1564,N1565,N1566,
     N1567,N1568,N1569,N1570,N1571,N1572,N1573,N1574,N1575,N1576,
     N1577,N1578,N1581,N1582,N1585,N1588,N1591,N1596,N1600,N1606,
     N1612,N1615,N1619,N1624,N1628,N1631,N1634,N1637,N1642,N1647,
     N1651,N1656,N1676,N1681,N1686,N1690,N1708,N1770,N1773,N1776,
     N1777,N1778,N1781,N1784,N1785,N1795,N1798,N1801,N1804,N1807,
     N1808,N1809,N1810,N1811,N1813,N1814,N1815,N1822,N1823,N1824,
     N1827,N1830,N1831,N1832,N1833,N1836,N1841,N1848,N1852,N1856,
     N1863,N1870,N1875,N1880,N1885,N1888,N1891,N1894,N1897,N1908,
     N1909,N1910,N1911,N1912,N1913,N1914,N1915,N1916,N1917,N1918,
     N1919,N1928,N1929,N1930,N1931,N1932,N1933,N1934,N1935,N1936,
     N1939,N1940,N1941,N1942,N1945,N1948,N1951,N1954,N1957,N1960,
     N1963,N1966,N2028,N2029,N2030,N2031,N2032,N2033,N2034,N2040,
     N2041,N2042,N2043,N2046,N2049,N2052,N2055,N2058,N2061,N2064,
     N2067,N2070,N2073,N2076,N2079,N2095,N2098,N2101,N2104,N2107,
     N2110,N2113,N2119,N2120,N2125,N2126,N2127,N2128,N2135,N2141,
     N2144,N2147,N2150,N2153,N2154,N2155,N2156,N2157,N2158,N2171,
     N2172,N2173,N2174,N2175,N2176,N2177,N2178,N2185,N2188,N2191,
     N2194,N2197,N2200,N2201,N2204,N2207,N2210,N2213,N2216,N2219,
     N2234,N2235,N2236,N2237,N2250,N2266,N2269,N2291,N2294,N2297,
     N2298,N2300,N2301,N2302,N2303,N2304,N2305,N2306,N2307,N2308,
     N2309,N2310,N2311,N2312,N2313,N2314,N2315,N2316,N2317,N2318,
     N2319,N2320,N2321,N2322,N2323,N2324,N2325,N2326,N2327,N2328,
     N2329,N2330,N2331,N2332,N2333,N2334,N2335,N2336,N2337,N2338,
     N2339,N2340,N2354,N2355,N2356,N2357,N2358,N2359,N2364,N2365,
     N2366,N2367,N2368,N2372,N2373,N2374,N2375,N2376,N2377,N2382,
     N2386,N2391,N2395,N2400,N2403,N2406,N2407,N2408,N2409,N2410,
     N2411,N2412,N2413,N2414,N2415,N2416,N2417,N2421,N2425,N2428,
     N2429,N2430,N2431,N2432,N2433,N2434,N2437,N2440,N2443,N2446,
     N2449,N2452,N2453,N2454,N2457,N2460,N2463,N2466,N2469,N2472,
     N2475,N2478,N2481,N2484,N2487,N2490,N2493,N2503,N2504,N2510,
     N2511,N2521,N2528,N2531,N2534,N2537,N2540,N2544,N2545,N2546,
     N2547,N2548,N2549,N2550,N2551,N2552,N2553,N2563,N2564,N2565,
     N2566,N2567,N2568,N2579,N2603,N2607,N2608,N2609,N2610,N2611,
     N2612,N2613,N2617,N2618,N2619,N2620,N2621,N2624,N2628,N2629,
     N2630,N2631,N2632,N2633,N2634,N2635,N2636,N2638,N2645,N2646,
     N2652,N2655,N2656,N2659,N2663,N2664,N2665,N2666,N2667,N2668,
     N2669,N2670,N2671,N2672,N2673,N2674,N2675,N2676,N2677,N2678,
     N2679,N2680,N2681,N2684,N2687,N2690,N2693,N2694,N2695,N2696,
     N2697,N2698,N2699,N2700,N2701,N2702,N2703,N2706,N2707,N2708,
     N2709,N2710,N2719,N2720,N2726,N2729,N2738,N2743,N2747,N2748,
     N2749,N2750,N2751,N2760,N2761,N2766,N2771,N2772,N2773,N2774,
     N2775,N2776,N2777,N2778,N2781,N2782,N2783,N2784,N2789,N2790,
     N2791,N2792,N2793,N2796,N2800,N2803,N2806,N2809,N2810,N2811,
     N2812,N2817,N2820,N2826,N2829,N2830,N2831,N2837,N2838,N2839,
     N2840,N2841,N2844,N2854,N2859,N2869,N2874,N2877,N2880,N2881,
     N2882,N2885,N2888,N2894,N2895,N2896,N2897,N2898,N2899,N2900,
     N2901,N2914,N2915,N2916,N2917,N2918,N2919,N2920,N2921,N2931,
     N2938,N2939,N2963,N2972,N2975,N2978,N2981,N2984,N2985,N2986,
     N2989,N2992,N2995,N2998,N3001,N3004,N3007,N3008,N3009,N3010,
     N3013,N3016,N3019,N3022,N3025,N3028,N3029,N3030,N3035,N3036,
     N3037,N3039,N3044,N3045,N3046,N3047,N3048,N3049,N3050,N3053,
     N3054,N3055,N3056,N3057,N3058,N3059,N3060,N3061,N3064,N3065,
     N3066,N3067,N3068,N3069,N3070,N3071,N3072,N3073,N3074,N3075,
     N3076,N3088,N3091,N3110,N3113,N3137,N3140,N3143,N3146,N3149,
     N3152,N3157,N3160,N3163,N3166,N3169,N3172,N3175,N3176,N3177,
     N3178,N3180,N3187,N3188,N3189,N3190,N3191,N3192,N3193,N3194,
     N3195,N3196,N3197,N3208,N3215,N3216,N3217,N3218,N3219,N3220,
     N3222,N3223,N3230,N3231,N3238,N3241,N3244,N3247,N3250,N3253,
     N3256,N3259,N3262,N3265,N3268,N3271,N3274,N3277,N3281,N3282,
     N3283,N3284,N3286,N3288,N3289,N3291,N3293,N3295,N3296,N3299,
     N3301,N3302,N3304,N3306,N3308,N3309,N3312,N3314,N3315,N3318,
     N3321,N3324,N3327,N3330,N3333,N3334,N3335,N3336,N3337,N3340,
     N3344,N3348,N3352,N3356,N3360,N3364,N3367,N3370,N3374,N3378,
     N3382,N3386,N3390,N3394,N3397,N3400,N3401,N3402,N3403,N3404,
     N3405,N3406,N3409,N3410,N3412,N3414,N3416,N3418,N3420,N3422,
     N3428,N3430,N3432,N3434,N3436,N3438,N3440,N3450,N3453,N3456,
     N3459,N3478,N3479,N3480,N3481,N3482,N3483,N3484,N3485,N3486,
     N3487,N3488,N3489,N3490,N3491,N3492,N3493,N3494,N3496,N3498,
     N3499,N3500,N3501,N3502,N3503,N3504,N3505,N3506,N3507,N3508,
     N3509,N3510,N3511,N3512,N3513,N3515,N3517,N3522,N3525,N3528,
     N3531,N3534,N3537,N3540,N3543,N3551,N3552,N3553,N3554,N3555,
     N3556,N3557,N3558,N3559,N3563,N3564,N3565,N3566,N3567,N3568,
     N3569,N3570,N3576,N3579,N3585,N3588,N3592,N3593,N3594,N3595,
     N3596,N3597,N3598,N3599,N3600,N3603,N3608,N3612,N3615,N3616,
     N3622,N3629,N3630,N3631,N3632,N3633,N3634,N3635,N3640,N3644,
     N3647,N3648,N3654,N3661,N3662,N3667,N3668,N3669,N3670,N3691,
     N3692,N3693,N3694,N3695,N3696,N3697,N3716,N3717,N3718,N3719,
     N3720,N3721,N3722,N3723,N3726,N3727,N3728,N3729,N3730,N3731,
     N3732,N3733,N3734,N3735,N3736,N3737,N3740,N3741,N3742,N3743,
     N3744,N3745,N3746,N3747,N3748,N3749,N3750,N3753,N3754,N3758,
     N3761,N3762,N3767,N3771,N3774,N3775,N3778,N3779,N3780,N3790,
     N3793,N3794,N3802,N3805,N3806,N3807,N3808,N3811,N3812,N3813,
     N3814,N3815,N3816,N3817,N3818,N3819,N3820,N3821,N3822,N3823,
     N3826,N3827,N3834,N3835,N3836,N3837,N3838,N3839,N3840,N3843,
     N3852,N3857,N3858,N3859,N3864,N3869,N3870,N3876,N3877, gate1044inter0, gate1044inter1, gate1044inter2, gate1044inter3, gate1044inter4, gate1044inter5, gate1044inter6, gate1044inter7, gate1044inter8, gate1044inter9, gate1044inter10, gate1044inter11, gate1044inter12, gate526inter0, gate526inter1, gate526inter2, gate526inter3, gate526inter4, gate526inter5, gate526inter6, gate526inter7, gate526inter8, gate526inter9, gate526inter10, gate526inter11, gate526inter12, gate743inter0, gate743inter1, gate743inter2, gate743inter3, gate743inter4, gate743inter5, gate743inter6, gate743inter7, gate743inter8, gate743inter9, gate743inter10, gate743inter11, gate743inter12, gate1025inter0, gate1025inter1, gate1025inter2, gate1025inter3, gate1025inter4, gate1025inter5, gate1025inter6, gate1025inter7, gate1025inter8, gate1025inter9, gate1025inter10, gate1025inter11, gate1025inter12, gate885inter0, gate885inter1, gate885inter2, gate885inter3, gate885inter4, gate885inter5, gate885inter6, gate885inter7, gate885inter8, gate885inter9, gate885inter10, gate885inter11, gate885inter12, gate626inter0, gate626inter1, gate626inter2, gate626inter3, gate626inter4, gate626inter5, gate626inter6, gate626inter7, gate626inter8, gate626inter9, gate626inter10, gate626inter11, gate626inter12, gate1115inter0, gate1115inter1, gate1115inter2, gate1115inter3, gate1115inter4, gate1115inter5, gate1115inter6, gate1115inter7, gate1115inter8, gate1115inter9, gate1115inter10, gate1115inter11, gate1115inter12, gate586inter0, gate586inter1, gate586inter2, gate586inter3, gate586inter4, gate586inter5, gate586inter6, gate586inter7, gate586inter8, gate586inter9, gate586inter10, gate586inter11, gate586inter12, gate1093inter0, gate1093inter1, gate1093inter2, gate1093inter3, gate1093inter4, gate1093inter5, gate1093inter6, gate1093inter7, gate1093inter8, gate1093inter9, gate1093inter10, gate1093inter11, gate1093inter12, gate1034inter0, gate1034inter1, gate1034inter2, gate1034inter3, gate1034inter4, gate1034inter5, gate1034inter6, gate1034inter7, gate1034inter8, gate1034inter9, gate1034inter10, gate1034inter11, gate1034inter12, gate598inter0, gate598inter1, gate598inter2, gate598inter3, gate598inter4, gate598inter5, gate598inter6, gate598inter7, gate598inter8, gate598inter9, gate598inter10, gate598inter11, gate598inter12, gate886inter0, gate886inter1, gate886inter2, gate886inter3, gate886inter4, gate886inter5, gate886inter6, gate886inter7, gate886inter8, gate886inter9, gate886inter10, gate886inter11, gate886inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate1082inter0, gate1082inter1, gate1082inter2, gate1082inter3, gate1082inter4, gate1082inter5, gate1082inter6, gate1082inter7, gate1082inter8, gate1082inter9, gate1082inter10, gate1082inter11, gate1082inter12, gate883inter0, gate883inter1, gate883inter2, gate883inter3, gate883inter4, gate883inter5, gate883inter6, gate883inter7, gate883inter8, gate883inter9, gate883inter10, gate883inter11, gate883inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate1108inter0, gate1108inter1, gate1108inter2, gate1108inter3, gate1108inter4, gate1108inter5, gate1108inter6, gate1108inter7, gate1108inter8, gate1108inter9, gate1108inter10, gate1108inter11, gate1108inter12, gate661inter0, gate661inter1, gate661inter2, gate661inter3, gate661inter4, gate661inter5, gate661inter6, gate661inter7, gate661inter8, gate661inter9, gate661inter10, gate661inter11, gate661inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate594inter0, gate594inter1, gate594inter2, gate594inter3, gate594inter4, gate594inter5, gate594inter6, gate594inter7, gate594inter8, gate594inter9, gate594inter10, gate594inter11, gate594inter12, gate1124inter0, gate1124inter1, gate1124inter2, gate1124inter3, gate1124inter4, gate1124inter5, gate1124inter6, gate1124inter7, gate1124inter8, gate1124inter9, gate1124inter10, gate1124inter11, gate1124inter12, gate763inter0, gate763inter1, gate763inter2, gate763inter3, gate763inter4, gate763inter5, gate763inter6, gate763inter7, gate763inter8, gate763inter9, gate763inter10, gate763inter11, gate763inter12, gate1094inter0, gate1094inter1, gate1094inter2, gate1094inter3, gate1094inter4, gate1094inter5, gate1094inter6, gate1094inter7, gate1094inter8, gate1094inter9, gate1094inter10, gate1094inter11, gate1094inter12, gate520inter0, gate520inter1, gate520inter2, gate520inter3, gate520inter4, gate520inter5, gate520inter6, gate520inter7, gate520inter8, gate520inter9, gate520inter10, gate520inter11, gate520inter12, gate887inter0, gate887inter1, gate887inter2, gate887inter3, gate887inter4, gate887inter5, gate887inter6, gate887inter7, gate887inter8, gate887inter9, gate887inter10, gate887inter11, gate887inter12, gate1125inter0, gate1125inter1, gate1125inter2, gate1125inter3, gate1125inter4, gate1125inter5, gate1125inter6, gate1125inter7, gate1125inter8, gate1125inter9, gate1125inter10, gate1125inter11, gate1125inter12, gate930inter0, gate930inter1, gate930inter2, gate930inter3, gate930inter4, gate930inter5, gate930inter6, gate930inter7, gate930inter8, gate930inter9, gate930inter10, gate930inter11, gate930inter12, gate1123inter0, gate1123inter1, gate1123inter2, gate1123inter3, gate1123inter4, gate1123inter5, gate1123inter6, gate1123inter7, gate1123inter8, gate1123inter9, gate1123inter10, gate1123inter11, gate1123inter12, gate1064inter0, gate1064inter1, gate1064inter2, gate1064inter3, gate1064inter4, gate1064inter5, gate1064inter6, gate1064inter7, gate1064inter8, gate1064inter9, gate1064inter10, gate1064inter11, gate1064inter12, gate1066inter0, gate1066inter1, gate1066inter2, gate1066inter3, gate1066inter4, gate1066inter5, gate1066inter6, gate1066inter7, gate1066inter8, gate1066inter9, gate1066inter10, gate1066inter11, gate1066inter12, gate635inter0, gate635inter1, gate635inter2, gate635inter3, gate635inter4, gate635inter5, gate635inter6, gate635inter7, gate635inter8, gate635inter9, gate635inter10, gate635inter11, gate635inter12, gate590inter0, gate590inter1, gate590inter2, gate590inter3, gate590inter4, gate590inter5, gate590inter6, gate590inter7, gate590inter8, gate590inter9, gate590inter10, gate590inter11, gate590inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate1101inter0, gate1101inter1, gate1101inter2, gate1101inter3, gate1101inter4, gate1101inter5, gate1101inter6, gate1101inter7, gate1101inter8, gate1101inter9, gate1101inter10, gate1101inter11, gate1101inter12, gate587inter0, gate587inter1, gate587inter2, gate587inter3, gate587inter4, gate587inter5, gate587inter6, gate587inter7, gate587inter8, gate587inter9, gate587inter10, gate587inter11, gate587inter12, gate1073inter0, gate1073inter1, gate1073inter2, gate1073inter3, gate1073inter4, gate1073inter5, gate1073inter6, gate1073inter7, gate1073inter8, gate1073inter9, gate1073inter10, gate1073inter11, gate1073inter12, gate545inter0, gate545inter1, gate545inter2, gate545inter3, gate545inter4, gate545inter5, gate545inter6, gate545inter7, gate545inter8, gate545inter9, gate545inter10, gate545inter11, gate545inter12, gate317inter0, gate317inter1, gate317inter2, gate317inter3, gate317inter4, gate317inter5, gate317inter6, gate317inter7, gate317inter8, gate317inter9, gate317inter10, gate317inter11, gate317inter12, gate733inter0, gate733inter1, gate733inter2, gate733inter3, gate733inter4, gate733inter5, gate733inter6, gate733inter7, gate733inter8, gate733inter9, gate733inter10, gate733inter11, gate733inter12, gate625inter0, gate625inter1, gate625inter2, gate625inter3, gate625inter4, gate625inter5, gate625inter6, gate625inter7, gate625inter8, gate625inter9, gate625inter10, gate625inter11, gate625inter12, gate738inter0, gate738inter1, gate738inter2, gate738inter3, gate738inter4, gate738inter5, gate738inter6, gate738inter7, gate738inter8, gate738inter9, gate738inter10, gate738inter11, gate738inter12, gate358inter0, gate358inter1, gate358inter2, gate358inter3, gate358inter4, gate358inter5, gate358inter6, gate358inter7, gate358inter8, gate358inter9, gate358inter10, gate358inter11, gate358inter12, gate1182inter0, gate1182inter1, gate1182inter2, gate1182inter3, gate1182inter4, gate1182inter5, gate1182inter6, gate1182inter7, gate1182inter8, gate1182inter9, gate1182inter10, gate1182inter11, gate1182inter12, gate737inter0, gate737inter1, gate737inter2, gate737inter3, gate737inter4, gate737inter5, gate737inter6, gate737inter7, gate737inter8, gate737inter9, gate737inter10, gate737inter11, gate737inter12, gate551inter0, gate551inter1, gate551inter2, gate551inter3, gate551inter4, gate551inter5, gate551inter6, gate551inter7, gate551inter8, gate551inter9, gate551inter10, gate551inter11, gate551inter12, gate645inter0, gate645inter1, gate645inter2, gate645inter3, gate645inter4, gate645inter5, gate645inter6, gate645inter7, gate645inter8, gate645inter9, gate645inter10, gate645inter11, gate645inter12, gate1046inter0, gate1046inter1, gate1046inter2, gate1046inter3, gate1046inter4, gate1046inter5, gate1046inter6, gate1046inter7, gate1046inter8, gate1046inter9, gate1046inter10, gate1046inter11, gate1046inter12, gate591inter0, gate591inter1, gate591inter2, gate591inter3, gate591inter4, gate591inter5, gate591inter6, gate591inter7, gate591inter8, gate591inter9, gate591inter10, gate591inter11, gate591inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate641inter0, gate641inter1, gate641inter2, gate641inter3, gate641inter4, gate641inter5, gate641inter6, gate641inter7, gate641inter8, gate641inter9, gate641inter10, gate641inter11, gate641inter12, gate739inter0, gate739inter1, gate739inter2, gate739inter3, gate739inter4, gate739inter5, gate739inter6, gate739inter7, gate739inter8, gate739inter9, gate739inter10, gate739inter11, gate739inter12, gate680inter0, gate680inter1, gate680inter2, gate680inter3, gate680inter4, gate680inter5, gate680inter6, gate680inter7, gate680inter8, gate680inter9, gate680inter10, gate680inter11, gate680inter12, gate1077inter0, gate1077inter1, gate1077inter2, gate1077inter3, gate1077inter4, gate1077inter5, gate1077inter6, gate1077inter7, gate1077inter8, gate1077inter9, gate1077inter10, gate1077inter11, gate1077inter12, gate1140inter0, gate1140inter1, gate1140inter2, gate1140inter3, gate1140inter4, gate1140inter5, gate1140inter6, gate1140inter7, gate1140inter8, gate1140inter9, gate1140inter10, gate1140inter11, gate1140inter12, gate1098inter0, gate1098inter1, gate1098inter2, gate1098inter3, gate1098inter4, gate1098inter5, gate1098inter6, gate1098inter7, gate1098inter8, gate1098inter9, gate1098inter10, gate1098inter11, gate1098inter12, gate584inter0, gate584inter1, gate584inter2, gate584inter3, gate584inter4, gate584inter5, gate584inter6, gate584inter7, gate584inter8, gate584inter9, gate584inter10, gate584inter11, gate584inter12, gate754inter0, gate754inter1, gate754inter2, gate754inter3, gate754inter4, gate754inter5, gate754inter6, gate754inter7, gate754inter8, gate754inter9, gate754inter10, gate754inter11, gate754inter12, gate651inter0, gate651inter1, gate651inter2, gate651inter3, gate651inter4, gate651inter5, gate651inter6, gate651inter7, gate651inter8, gate651inter9, gate651inter10, gate651inter11, gate651inter12, gate1055inter0, gate1055inter1, gate1055inter2, gate1055inter3, gate1055inter4, gate1055inter5, gate1055inter6, gate1055inter7, gate1055inter8, gate1055inter9, gate1055inter10, gate1055inter11, gate1055inter12, gate595inter0, gate595inter1, gate595inter2, gate595inter3, gate595inter4, gate595inter5, gate595inter6, gate595inter7, gate595inter8, gate595inter9, gate595inter10, gate595inter11, gate595inter12, gate1004inter0, gate1004inter1, gate1004inter2, gate1004inter3, gate1004inter4, gate1004inter5, gate1004inter6, gate1004inter7, gate1004inter8, gate1004inter9, gate1004inter10, gate1004inter11, gate1004inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate1023inter0, gate1023inter1, gate1023inter2, gate1023inter3, gate1023inter4, gate1023inter5, gate1023inter6, gate1023inter7, gate1023inter8, gate1023inter9, gate1023inter10, gate1023inter11, gate1023inter12, gate1048inter0, gate1048inter1, gate1048inter2, gate1048inter3, gate1048inter4, gate1048inter5, gate1048inter6, gate1048inter7, gate1048inter8, gate1048inter9, gate1048inter10, gate1048inter11, gate1048inter12, gate534inter0, gate534inter1, gate534inter2, gate534inter3, gate534inter4, gate534inter5, gate534inter6, gate534inter7, gate534inter8, gate534inter9, gate534inter10, gate534inter11, gate534inter12, gate518inter0, gate518inter1, gate518inter2, gate518inter3, gate518inter4, gate518inter5, gate518inter6, gate518inter7, gate518inter8, gate518inter9, gate518inter10, gate518inter11, gate518inter12, gate777inter0, gate777inter1, gate777inter2, gate777inter3, gate777inter4, gate777inter5, gate777inter6, gate777inter7, gate777inter8, gate777inter9, gate777inter10, gate777inter11, gate777inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate685inter0, gate685inter1, gate685inter2, gate685inter3, gate685inter4, gate685inter5, gate685inter6, gate685inter7, gate685inter8, gate685inter9, gate685inter10, gate685inter11, gate685inter12, gate1072inter0, gate1072inter1, gate1072inter2, gate1072inter3, gate1072inter4, gate1072inter5, gate1072inter6, gate1072inter7, gate1072inter8, gate1072inter9, gate1072inter10, gate1072inter11, gate1072inter12, gate1136inter0, gate1136inter1, gate1136inter2, gate1136inter3, gate1136inter4, gate1136inter5, gate1136inter6, gate1136inter7, gate1136inter8, gate1136inter9, gate1136inter10, gate1136inter11, gate1136inter12, gate522inter0, gate522inter1, gate522inter2, gate522inter3, gate522inter4, gate522inter5, gate522inter6, gate522inter7, gate522inter8, gate522inter9, gate522inter10, gate522inter11, gate522inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate638inter0, gate638inter1, gate638inter2, gate638inter3, gate638inter4, gate638inter5, gate638inter6, gate638inter7, gate638inter8, gate638inter9, gate638inter10, gate638inter11, gate638inter12, gate537inter0, gate537inter1, gate537inter2, gate537inter3, gate537inter4, gate537inter5, gate537inter6, gate537inter7, gate537inter8, gate537inter9, gate537inter10, gate537inter11, gate537inter12, gate736inter0, gate736inter1, gate736inter2, gate736inter3, gate736inter4, gate736inter5, gate736inter6, gate736inter7, gate736inter8, gate736inter9, gate736inter10, gate736inter11, gate736inter12, gate1105inter0, gate1105inter1, gate1105inter2, gate1105inter3, gate1105inter4, gate1105inter5, gate1105inter6, gate1105inter7, gate1105inter8, gate1105inter9, gate1105inter10, gate1105inter11, gate1105inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate1092inter0, gate1092inter1, gate1092inter2, gate1092inter3, gate1092inter4, gate1092inter5, gate1092inter6, gate1092inter7, gate1092inter8, gate1092inter9, gate1092inter10, gate1092inter11, gate1092inter12, gate910inter0, gate910inter1, gate910inter2, gate910inter3, gate910inter4, gate910inter5, gate910inter6, gate910inter7, gate910inter8, gate910inter9, gate910inter10, gate910inter11, gate910inter12, gate779inter0, gate779inter1, gate779inter2, gate779inter3, gate779inter4, gate779inter5, gate779inter6, gate779inter7, gate779inter8, gate779inter9, gate779inter10, gate779inter11, gate779inter12, gate1085inter0, gate1085inter1, gate1085inter2, gate1085inter3, gate1085inter4, gate1085inter5, gate1085inter6, gate1085inter7, gate1085inter8, gate1085inter9, gate1085inter10, gate1085inter11, gate1085inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate724inter0, gate724inter1, gate724inter2, gate724inter3, gate724inter4, gate724inter5, gate724inter6, gate724inter7, gate724inter8, gate724inter9, gate724inter10, gate724inter11, gate724inter12, gate627inter0, gate627inter1, gate627inter2, gate627inter3, gate627inter4, gate627inter5, gate627inter6, gate627inter7, gate627inter8, gate627inter9, gate627inter10, gate627inter11, gate627inter12, gate753inter0, gate753inter1, gate753inter2, gate753inter3, gate753inter4, gate753inter5, gate753inter6, gate753inter7, gate753inter8, gate753inter9, gate753inter10, gate753inter11, gate753inter12, gate301inter0, gate301inter1, gate301inter2, gate301inter3, gate301inter4, gate301inter5, gate301inter6, gate301inter7, gate301inter8, gate301inter9, gate301inter10, gate301inter11, gate301inter12, gate609inter0, gate609inter1, gate609inter2, gate609inter3, gate609inter4, gate609inter5, gate609inter6, gate609inter7, gate609inter8, gate609inter9, gate609inter10, gate609inter11, gate609inter12, gate971inter0, gate971inter1, gate971inter2, gate971inter3, gate971inter4, gate971inter5, gate971inter6, gate971inter7, gate971inter8, gate971inter9, gate971inter10, gate971inter11, gate971inter12, gate776inter0, gate776inter1, gate776inter2, gate776inter3, gate776inter4, gate776inter5, gate776inter6, gate776inter7, gate776inter8, gate776inter9, gate776inter10, gate776inter11, gate776inter12, gate601inter0, gate601inter1, gate601inter2, gate601inter3, gate601inter4, gate601inter5, gate601inter6, gate601inter7, gate601inter8, gate601inter9, gate601inter10, gate601inter11, gate601inter12, gate975inter0, gate975inter1, gate975inter2, gate975inter3, gate975inter4, gate975inter5, gate975inter6, gate975inter7, gate975inter8, gate975inter9, gate975inter10, gate975inter11, gate975inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate716inter0, gate716inter1, gate716inter2, gate716inter3, gate716inter4, gate716inter5, gate716inter6, gate716inter7, gate716inter8, gate716inter9, gate716inter10, gate716inter11, gate716inter12, gate1116inter0, gate1116inter1, gate1116inter2, gate1116inter3, gate1116inter4, gate1116inter5, gate1116inter6, gate1116inter7, gate1116inter8, gate1116inter9, gate1116inter10, gate1116inter11, gate1116inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate783inter0, gate783inter1, gate783inter2, gate783inter3, gate783inter4, gate783inter5, gate783inter6, gate783inter7, gate783inter8, gate783inter9, gate783inter10, gate783inter11, gate783inter12, gate557inter0, gate557inter1, gate557inter2, gate557inter3, gate557inter4, gate557inter5, gate557inter6, gate557inter7, gate557inter8, gate557inter9, gate557inter10, gate557inter11, gate557inter12, gate1087inter0, gate1087inter1, gate1087inter2, gate1087inter3, gate1087inter4, gate1087inter5, gate1087inter6, gate1087inter7, gate1087inter8, gate1087inter9, gate1087inter10, gate1087inter11, gate1087inter12, gate524inter0, gate524inter1, gate524inter2, gate524inter3, gate524inter4, gate524inter5, gate524inter6, gate524inter7, gate524inter8, gate524inter9, gate524inter10, gate524inter11, gate524inter12, gate620inter0, gate620inter1, gate620inter2, gate620inter3, gate620inter4, gate620inter5, gate620inter6, gate620inter7, gate620inter8, gate620inter9, gate620inter10, gate620inter11, gate620inter12, gate1051inter0, gate1051inter1, gate1051inter2, gate1051inter3, gate1051inter4, gate1051inter5, gate1051inter6, gate1051inter7, gate1051inter8, gate1051inter9, gate1051inter10, gate1051inter11, gate1051inter12, gate321inter0, gate321inter1, gate321inter2, gate321inter3, gate321inter4, gate321inter5, gate321inter6, gate321inter7, gate321inter8, gate321inter9, gate321inter10, gate321inter11, gate321inter12, gate630inter0, gate630inter1, gate630inter2, gate630inter3, gate630inter4, gate630inter5, gate630inter6, gate630inter7, gate630inter8, gate630inter9, gate630inter10, gate630inter11, gate630inter12, gate1100inter0, gate1100inter1, gate1100inter2, gate1100inter3, gate1100inter4, gate1100inter5, gate1100inter6, gate1100inter7, gate1100inter8, gate1100inter9, gate1100inter10, gate1100inter11, gate1100inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate756inter0, gate756inter1, gate756inter2, gate756inter3, gate756inter4, gate756inter5, gate756inter6, gate756inter7, gate756inter8, gate756inter9, gate756inter10, gate756inter11, gate756inter12, gate556inter0, gate556inter1, gate556inter2, gate556inter3, gate556inter4, gate556inter5, gate556inter6, gate556inter7, gate556inter8, gate556inter9, gate556inter10, gate556inter11, gate556inter12, gate928inter0, gate928inter1, gate928inter2, gate928inter3, gate928inter4, gate928inter5, gate928inter6, gate928inter7, gate928inter8, gate928inter9, gate928inter10, gate928inter11, gate928inter12, gate530inter0, gate530inter1, gate530inter2, gate530inter3, gate530inter4, gate530inter5, gate530inter6, gate530inter7, gate530inter8, gate530inter9, gate530inter10, gate530inter11, gate530inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate1012inter0, gate1012inter1, gate1012inter2, gate1012inter3, gate1012inter4, gate1012inter5, gate1012inter6, gate1012inter7, gate1012inter8, gate1012inter9, gate1012inter10, gate1012inter11, gate1012inter12, gate722inter0, gate722inter1, gate722inter2, gate722inter3, gate722inter4, gate722inter5, gate722inter6, gate722inter7, gate722inter8, gate722inter9, gate722inter10, gate722inter11, gate722inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate662inter0, gate662inter1, gate662inter2, gate662inter3, gate662inter4, gate662inter5, gate662inter6, gate662inter7, gate662inter8, gate662inter9, gate662inter10, gate662inter11, gate662inter12, gate1107inter0, gate1107inter1, gate1107inter2, gate1107inter3, gate1107inter4, gate1107inter5, gate1107inter6, gate1107inter7, gate1107inter8, gate1107inter9, gate1107inter10, gate1107inter11, gate1107inter12, gate979inter0, gate979inter1, gate979inter2, gate979inter3, gate979inter4, gate979inter5, gate979inter6, gate979inter7, gate979inter8, gate979inter9, gate979inter10, gate979inter11, gate979inter12, gate896inter0, gate896inter1, gate896inter2, gate896inter3, gate896inter4, gate896inter5, gate896inter6, gate896inter7, gate896inter8, gate896inter9, gate896inter10, gate896inter11, gate896inter12, gate320inter0, gate320inter1, gate320inter2, gate320inter3, gate320inter4, gate320inter5, gate320inter6, gate320inter7, gate320inter8, gate320inter9, gate320inter10, gate320inter11, gate320inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate1002inter0, gate1002inter1, gate1002inter2, gate1002inter3, gate1002inter4, gate1002inter5, gate1002inter6, gate1002inter7, gate1002inter8, gate1002inter9, gate1002inter10, gate1002inter11, gate1002inter12;


buf1 gate1( .a(N219), .O(N398) );
buf1 gate2( .a(N219), .O(N400) );
buf1 gate3( .a(N219), .O(N401) );
and2 gate4( .a(N1), .b(N3), .O(N405) );
inv1 gate5( .a(N230), .O(N408) );
buf1 gate6( .a(N253), .O(N419) );
buf1 gate7( .a(N253), .O(N420) );
inv1 gate8( .a(N262), .O(N425) );
buf1 gate9( .a(N290), .O(N456) );
buf1 gate10( .a(N290), .O(N457) );
buf1 gate11( .a(N290), .O(N458) );
and4 gate12( .a(N309), .b(N305), .c(N301), .d(N297), .O(N485) );
inv1 gate13( .a(N405), .O(N486) );
inv1 gate14( .a(N44), .O(N487) );
inv1 gate15( .a(N132), .O(N488) );
inv1 gate16( .a(N82), .O(N489) );
inv1 gate17( .a(N96), .O(N490) );
inv1 gate18( .a(N69), .O(N491) );
inv1 gate19( .a(N120), .O(N492) );
inv1 gate20( .a(N57), .O(N493) );
inv1 gate21( .a(N108), .O(N494) );
and3 gate22( .a(N2), .b(N15), .c(N237), .O(N495) );
buf1 gate23( .a(N237), .O(N496) );
and2 gate24( .a(N37), .b(N37), .O(N499) );
buf1 gate25( .a(N219), .O(N500) );
buf1 gate26( .a(N8), .O(N503) );
buf1 gate27( .a(N8), .O(N506) );
buf1 gate28( .a(N227), .O(N509) );
buf1 gate29( .a(N234), .O(N521) );
inv1 gate30( .a(N241), .O(N533) );
inv1 gate31( .a(N246), .O(N537) );
and2 gate32( .a(N11), .b(N246), .O(N543) );
and4 gate33( .a(N132), .b(N82), .c(N96), .d(N44), .O(N544) );
and4 gate34( .a(N120), .b(N57), .c(N108), .d(N69), .O(N547) );
buf1 gate35( .a(N227), .O(N550) );
buf1 gate36( .a(N234), .O(N562) );
inv1 gate37( .a(N256), .O(N574) );
inv1 gate38( .a(N259), .O(N578) );
buf1 gate39( .a(N319), .O(N582) );
buf1 gate40( .a(N322), .O(N594) );
inv1 gate41( .a(N328), .O(N606) );
inv1 gate42( .a(N331), .O(N607) );
inv1 gate43( .a(N334), .O(N608) );
inv1 gate44( .a(N337), .O(N609) );
inv1 gate45( .a(N340), .O(N610) );
inv1 gate46( .a(N343), .O(N611) );
inv1 gate47( .a(N352), .O(N612) );
buf1 gate48( .a(N319), .O(N613) );
buf1 gate49( .a(N322), .O(N625) );
buf1 gate50( .a(N16), .O(N637) );
buf1 gate51( .a(N16), .O(N643) );
inv1 gate52( .a(N355), .O(N650) );
and2 gate53( .a(N7), .b(N237), .O(N651) );
inv1 gate54( .a(N263), .O(N655) );
inv1 gate55( .a(N266), .O(N659) );
inv1 gate56( .a(N269), .O(N663) );
inv1 gate57( .a(N272), .O(N667) );
inv1 gate58( .a(N275), .O(N671) );
inv1 gate59( .a(N278), .O(N675) );
inv1 gate60( .a(N281), .O(N679) );
inv1 gate61( .a(N284), .O(N683) );
inv1 gate62( .a(N287), .O(N687) );
buf1 gate63( .a(N29), .O(N693) );
buf1 gate64( .a(N29), .O(N699) );
inv1 gate65( .a(N294), .O(N705) );
inv1 gate66( .a(N297), .O(N711) );
inv1 gate67( .a(N301), .O(N715) );
inv1 gate68( .a(N305), .O(N719) );
inv1 gate69( .a(N309), .O(N723) );
inv1 gate70( .a(N313), .O(N727) );
inv1 gate71( .a(N316), .O(N730) );
inv1 gate72( .a(N346), .O(N733) );
inv1 gate73( .a(N349), .O(N734) );
buf1 gate74( .a(N259), .O(N735) );
buf1 gate75( .a(N256), .O(N738) );
buf1 gate76( .a(N263), .O(N741) );
buf1 gate77( .a(N269), .O(N744) );
buf1 gate78( .a(N266), .O(N747) );
buf1 gate79( .a(N275), .O(N750) );
buf1 gate80( .a(N272), .O(N753) );
buf1 gate81( .a(N281), .O(N756) );
buf1 gate82( .a(N278), .O(N759) );
buf1 gate83( .a(N287), .O(N762) );
buf1 gate84( .a(N284), .O(N765) );
buf1 gate85( .a(N294), .O(N768) );
buf1 gate86( .a(N301), .O(N771) );
buf1 gate87( .a(N297), .O(N774) );
buf1 gate88( .a(N309), .O(N777) );
buf1 gate89( .a(N305), .O(N780) );
buf1 gate90( .a(N316), .O(N783) );
buf1 gate91( .a(N313), .O(N786) );
inv1 gate92( .a(N485), .O(N792) );
inv1 gate93( .a(N495), .O(N799) );
inv1 gate94( .a(N499), .O(N800) );
buf1 gate95( .a(N500), .O(N805) );
nand2 gate96( .a(N331), .b(N606), .O(N900) );
nand2 gate97( .a(N328), .b(N607), .O(N901) );

  xor2  gate2320(.a(N608), .b(N337), .O(gate98inter0));
  nand2 gate2321(.a(gate98inter0), .b(s_150), .O(gate98inter1));
  and2  gate2322(.a(N608), .b(N337), .O(gate98inter2));
  inv1  gate2323(.a(s_150), .O(gate98inter3));
  inv1  gate2324(.a(s_151), .O(gate98inter4));
  nand2 gate2325(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate2326(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate2327(.a(N337), .O(gate98inter7));
  inv1  gate2328(.a(N608), .O(gate98inter8));
  nand2 gate2329(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate2330(.a(s_151), .b(gate98inter3), .O(gate98inter10));
  nor2  gate2331(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate2332(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate2333(.a(gate98inter12), .b(gate98inter1), .O(N902));

  xor2  gate2908(.a(N609), .b(N334), .O(gate99inter0));
  nand2 gate2909(.a(gate99inter0), .b(s_234), .O(gate99inter1));
  and2  gate2910(.a(N609), .b(N334), .O(gate99inter2));
  inv1  gate2911(.a(s_234), .O(gate99inter3));
  inv1  gate2912(.a(s_235), .O(gate99inter4));
  nand2 gate2913(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate2914(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate2915(.a(N334), .O(gate99inter7));
  inv1  gate2916(.a(N609), .O(gate99inter8));
  nand2 gate2917(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate2918(.a(s_235), .b(gate99inter3), .O(gate99inter10));
  nor2  gate2919(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate2920(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate2921(.a(gate99inter12), .b(gate99inter1), .O(N903));
nand2 gate100( .a(N343), .b(N610), .O(N904) );
nand2 gate101( .a(N340), .b(N611), .O(N905) );
nand2 gate102( .a(N349), .b(N733), .O(N998) );
nand2 gate103( .a(N346), .b(N734), .O(N999) );
and2 gate104( .a(N94), .b(N500), .O(N1026) );
and2 gate105( .a(N325), .b(N651), .O(N1027) );
inv1 gate106( .a(N651), .O(N1028) );

  xor2  gate1536(.a(N651), .b(N231), .O(gate107inter0));
  nand2 gate1537(.a(gate107inter0), .b(s_38), .O(gate107inter1));
  and2  gate1538(.a(N651), .b(N231), .O(gate107inter2));
  inv1  gate1539(.a(s_38), .O(gate107inter3));
  inv1  gate1540(.a(s_39), .O(gate107inter4));
  nand2 gate1541(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate1542(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate1543(.a(N231), .O(gate107inter7));
  inv1  gate1544(.a(N651), .O(gate107inter8));
  nand2 gate1545(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate1546(.a(s_39), .b(gate107inter3), .O(gate107inter10));
  nor2  gate1547(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate1548(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate1549(.a(gate107inter12), .b(gate107inter1), .O(N1029));
inv1 gate108( .a(N544), .O(N1032) );
inv1 gate109( .a(N547), .O(N1033) );
and2 gate110( .a(N547), .b(N544), .O(N1034) );
buf1 gate111( .a(N503), .O(N1037) );
inv1 gate112( .a(N509), .O(N1042) );
inv1 gate113( .a(N521), .O(N1053) );
and3 gate114( .a(N80), .b(N509), .c(N521), .O(N1064) );
and3 gate115( .a(N68), .b(N509), .c(N521), .O(N1065) );
and3 gate116( .a(N79), .b(N509), .c(N521), .O(N1066) );
and3 gate117( .a(N78), .b(N509), .c(N521), .O(N1067) );
and3 gate118( .a(N77), .b(N509), .c(N521), .O(N1068) );
and2 gate119( .a(N11), .b(N537), .O(N1069) );
buf1 gate120( .a(N503), .O(N1070) );
inv1 gate121( .a(N550), .O(N1075) );
inv1 gate122( .a(N562), .O(N1086) );
and3 gate123( .a(N76), .b(N550), .c(N562), .O(N1097) );
and3 gate124( .a(N75), .b(N550), .c(N562), .O(N1098) );
and3 gate125( .a(N74), .b(N550), .c(N562), .O(N1099) );
and3 gate126( .a(N73), .b(N550), .c(N562), .O(N1100) );
and3 gate127( .a(N72), .b(N550), .c(N562), .O(N1101) );
inv1 gate128( .a(N582), .O(N1102) );
inv1 gate129( .a(N594), .O(N1113) );
and3 gate130( .a(N114), .b(N582), .c(N594), .O(N1124) );
and3 gate131( .a(N113), .b(N582), .c(N594), .O(N1125) );
and3 gate132( .a(N112), .b(N582), .c(N594), .O(N1126) );
and3 gate133( .a(N111), .b(N582), .c(N594), .O(N1127) );
and2 gate134( .a(N582), .b(N594), .O(N1128) );
nand2 gate135( .a(N900), .b(N901), .O(N1129) );
nand2 gate136( .a(N902), .b(N903), .O(N1133) );

  xor2  gate2782(.a(N905), .b(N904), .O(gate137inter0));
  nand2 gate2783(.a(gate137inter0), .b(s_216), .O(gate137inter1));
  and2  gate2784(.a(N905), .b(N904), .O(gate137inter2));
  inv1  gate2785(.a(s_216), .O(gate137inter3));
  inv1  gate2786(.a(s_217), .O(gate137inter4));
  nand2 gate2787(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate2788(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate2789(.a(N904), .O(gate137inter7));
  inv1  gate2790(.a(N905), .O(gate137inter8));
  nand2 gate2791(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate2792(.a(s_217), .b(gate137inter3), .O(gate137inter10));
  nor2  gate2793(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate2794(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate2795(.a(gate137inter12), .b(gate137inter1), .O(N1137));
inv1 gate138( .a(N741), .O(N1140) );
nand2 gate139( .a(N741), .b(N612), .O(N1141) );
inv1 gate140( .a(N744), .O(N1142) );
inv1 gate141( .a(N747), .O(N1143) );
inv1 gate142( .a(N750), .O(N1144) );
inv1 gate143( .a(N753), .O(N1145) );
inv1 gate144( .a(N613), .O(N1146) );
inv1 gate145( .a(N625), .O(N1157) );
and3 gate146( .a(N118), .b(N613), .c(N625), .O(N1168) );
and3 gate147( .a(N107), .b(N613), .c(N625), .O(N1169) );
and3 gate148( .a(N117), .b(N613), .c(N625), .O(N1170) );
and3 gate149( .a(N116), .b(N613), .c(N625), .O(N1171) );
and3 gate150( .a(N115), .b(N613), .c(N625), .O(N1172) );
inv1 gate151( .a(N637), .O(N1173) );
inv1 gate152( .a(N643), .O(N1178) );
inv1 gate153( .a(N768), .O(N1184) );
nand2 gate154( .a(N768), .b(N650), .O(N1185) );
inv1 gate155( .a(N771), .O(N1186) );
inv1 gate156( .a(N774), .O(N1187) );
inv1 gate157( .a(N777), .O(N1188) );
inv1 gate158( .a(N780), .O(N1189) );
buf1 gate159( .a(N506), .O(N1190) );
buf1 gate160( .a(N506), .O(N1195) );
inv1 gate161( .a(N693), .O(N1200) );
inv1 gate162( .a(N699), .O(N1205) );
inv1 gate163( .a(N735), .O(N1210) );
inv1 gate164( .a(N738), .O(N1211) );
inv1 gate165( .a(N756), .O(N1212) );
inv1 gate166( .a(N759), .O(N1213) );
inv1 gate167( .a(N762), .O(N1214) );
inv1 gate168( .a(N765), .O(N1215) );
nand2 gate169( .a(N998), .b(N999), .O(N1216) );
buf1 gate170( .a(N574), .O(N1219) );
buf1 gate171( .a(N578), .O(N1222) );
buf1 gate172( .a(N655), .O(N1225) );
buf1 gate173( .a(N659), .O(N1228) );
buf1 gate174( .a(N663), .O(N1231) );
buf1 gate175( .a(N667), .O(N1234) );
buf1 gate176( .a(N671), .O(N1237) );
buf1 gate177( .a(N675), .O(N1240) );
buf1 gate178( .a(N679), .O(N1243) );
buf1 gate179( .a(N683), .O(N1246) );
inv1 gate180( .a(N783), .O(N1249) );
inv1 gate181( .a(N786), .O(N1250) );
buf1 gate182( .a(N687), .O(N1251) );
buf1 gate183( .a(N705), .O(N1254) );
buf1 gate184( .a(N711), .O(N1257) );
buf1 gate185( .a(N715), .O(N1260) );
buf1 gate186( .a(N719), .O(N1263) );
buf1 gate187( .a(N723), .O(N1266) );
inv1 gate188( .a(N1027), .O(N1269) );
and2 gate189( .a(N325), .b(N1032), .O(N1275) );
and2 gate190( .a(N231), .b(N1033), .O(N1276) );
buf1 gate191( .a(N1034), .O(N1277) );
or2 gate192( .a(N1069), .b(N543), .O(N1302) );

  xor2  gate1746(.a(N1140), .b(N352), .O(gate193inter0));
  nand2 gate1747(.a(gate193inter0), .b(s_68), .O(gate193inter1));
  and2  gate1748(.a(N1140), .b(N352), .O(gate193inter2));
  inv1  gate1749(.a(s_68), .O(gate193inter3));
  inv1  gate1750(.a(s_69), .O(gate193inter4));
  nand2 gate1751(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate1752(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate1753(.a(N352), .O(gate193inter7));
  inv1  gate1754(.a(N1140), .O(gate193inter8));
  nand2 gate1755(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate1756(.a(s_69), .b(gate193inter3), .O(gate193inter10));
  nor2  gate1757(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate1758(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate1759(.a(gate193inter12), .b(gate193inter1), .O(N1351));
nand2 gate194( .a(N747), .b(N1142), .O(N1352) );

  xor2  gate1480(.a(N1143), .b(N744), .O(gate195inter0));
  nand2 gate1481(.a(gate195inter0), .b(s_30), .O(gate195inter1));
  and2  gate1482(.a(N1143), .b(N744), .O(gate195inter2));
  inv1  gate1483(.a(s_30), .O(gate195inter3));
  inv1  gate1484(.a(s_31), .O(gate195inter4));
  nand2 gate1485(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate1486(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate1487(.a(N744), .O(gate195inter7));
  inv1  gate1488(.a(N1143), .O(gate195inter8));
  nand2 gate1489(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate1490(.a(s_31), .b(gate195inter3), .O(gate195inter10));
  nor2  gate1491(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate1492(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate1493(.a(gate195inter12), .b(gate195inter1), .O(N1353));

  xor2  gate1550(.a(N1144), .b(N753), .O(gate196inter0));
  nand2 gate1551(.a(gate196inter0), .b(s_40), .O(gate196inter1));
  and2  gate1552(.a(N1144), .b(N753), .O(gate196inter2));
  inv1  gate1553(.a(s_40), .O(gate196inter3));
  inv1  gate1554(.a(s_41), .O(gate196inter4));
  nand2 gate1555(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate1556(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate1557(.a(N753), .O(gate196inter7));
  inv1  gate1558(.a(N1144), .O(gate196inter8));
  nand2 gate1559(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate1560(.a(s_41), .b(gate196inter3), .O(gate196inter10));
  nor2  gate1561(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate1562(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate1563(.a(gate196inter12), .b(gate196inter1), .O(N1354));
nand2 gate197( .a(N750), .b(N1145), .O(N1355) );
nand2 gate198( .a(N355), .b(N1184), .O(N1395) );
nand2 gate199( .a(N774), .b(N1186), .O(N1396) );

  xor2  gate2460(.a(N1187), .b(N771), .O(gate200inter0));
  nand2 gate2461(.a(gate200inter0), .b(s_170), .O(gate200inter1));
  and2  gate2462(.a(N1187), .b(N771), .O(gate200inter2));
  inv1  gate2463(.a(s_170), .O(gate200inter3));
  inv1  gate2464(.a(s_171), .O(gate200inter4));
  nand2 gate2465(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate2466(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate2467(.a(N771), .O(gate200inter7));
  inv1  gate2468(.a(N1187), .O(gate200inter8));
  nand2 gate2469(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate2470(.a(s_171), .b(gate200inter3), .O(gate200inter10));
  nor2  gate2471(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate2472(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate2473(.a(gate200inter12), .b(gate200inter1), .O(N1397));

  xor2  gate2866(.a(N1188), .b(N780), .O(gate201inter0));
  nand2 gate2867(.a(gate201inter0), .b(s_228), .O(gate201inter1));
  and2  gate2868(.a(N1188), .b(N780), .O(gate201inter2));
  inv1  gate2869(.a(s_228), .O(gate201inter3));
  inv1  gate2870(.a(s_229), .O(gate201inter4));
  nand2 gate2871(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate2872(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate2873(.a(N780), .O(gate201inter7));
  inv1  gate2874(.a(N1188), .O(gate201inter8));
  nand2 gate2875(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate2876(.a(s_229), .b(gate201inter3), .O(gate201inter10));
  nor2  gate2877(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate2878(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate2879(.a(gate201inter12), .b(gate201inter1), .O(N1398));
nand2 gate202( .a(N777), .b(N1189), .O(N1399) );
nand2 gate203( .a(N738), .b(N1210), .O(N1422) );
nand2 gate204( .a(N735), .b(N1211), .O(N1423) );
nand2 gate205( .a(N759), .b(N1212), .O(N1424) );

  xor2  gate1438(.a(N1213), .b(N756), .O(gate206inter0));
  nand2 gate1439(.a(gate206inter0), .b(s_24), .O(gate206inter1));
  and2  gate1440(.a(N1213), .b(N756), .O(gate206inter2));
  inv1  gate1441(.a(s_24), .O(gate206inter3));
  inv1  gate1442(.a(s_25), .O(gate206inter4));
  nand2 gate1443(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate1444(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate1445(.a(N756), .O(gate206inter7));
  inv1  gate1446(.a(N1213), .O(gate206inter8));
  nand2 gate1447(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate1448(.a(s_25), .b(gate206inter3), .O(gate206inter10));
  nor2  gate1449(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate1450(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate1451(.a(gate206inter12), .b(gate206inter1), .O(N1425));
nand2 gate207( .a(N765), .b(N1214), .O(N1426) );

  xor2  gate2600(.a(N1215), .b(N762), .O(gate208inter0));
  nand2 gate2601(.a(gate208inter0), .b(s_190), .O(gate208inter1));
  and2  gate2602(.a(N1215), .b(N762), .O(gate208inter2));
  inv1  gate2603(.a(s_190), .O(gate208inter3));
  inv1  gate2604(.a(s_191), .O(gate208inter4));
  nand2 gate2605(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate2606(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate2607(.a(N762), .O(gate208inter7));
  inv1  gate2608(.a(N1215), .O(gate208inter8));
  nand2 gate2609(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate2610(.a(s_191), .b(gate208inter3), .O(gate208inter10));
  nor2  gate2611(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate2612(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate2613(.a(gate208inter12), .b(gate208inter1), .O(N1427));
nand2 gate209( .a(N786), .b(N1249), .O(N1440) );
nand2 gate210( .a(N783), .b(N1250), .O(N1441) );
inv1 gate211( .a(N1034), .O(N1448) );
inv1 gate212( .a(N1275), .O(N1449) );
inv1 gate213( .a(N1276), .O(N1450) );
and3 gate214( .a(N93), .b(N1042), .c(N1053), .O(N1451) );
and3 gate215( .a(N55), .b(N509), .c(N1053), .O(N1452) );
and3 gate216( .a(N67), .b(N1042), .c(N521), .O(N1453) );
and3 gate217( .a(N81), .b(N1042), .c(N1053), .O(N1454) );
and3 gate218( .a(N43), .b(N509), .c(N1053), .O(N1455) );
and3 gate219( .a(N56), .b(N1042), .c(N521), .O(N1456) );
and3 gate220( .a(N92), .b(N1042), .c(N1053), .O(N1457) );
and3 gate221( .a(N54), .b(N509), .c(N1053), .O(N1458) );
and3 gate222( .a(N66), .b(N1042), .c(N521), .O(N1459) );
and3 gate223( .a(N91), .b(N1042), .c(N1053), .O(N1460) );
and3 gate224( .a(N53), .b(N509), .c(N1053), .O(N1461) );
and3 gate225( .a(N65), .b(N1042), .c(N521), .O(N1462) );
and3 gate226( .a(N90), .b(N1042), .c(N1053), .O(N1463) );
and3 gate227( .a(N52), .b(N509), .c(N1053), .O(N1464) );
and3 gate228( .a(N64), .b(N1042), .c(N521), .O(N1465) );
and3 gate229( .a(N89), .b(N1075), .c(N1086), .O(N1466) );
and3 gate230( .a(N51), .b(N550), .c(N1086), .O(N1467) );
and3 gate231( .a(N63), .b(N1075), .c(N562), .O(N1468) );
and3 gate232( .a(N88), .b(N1075), .c(N1086), .O(N1469) );
and3 gate233( .a(N50), .b(N550), .c(N1086), .O(N1470) );
and3 gate234( .a(N62), .b(N1075), .c(N562), .O(N1471) );
and3 gate235( .a(N87), .b(N1075), .c(N1086), .O(N1472) );
and3 gate236( .a(N49), .b(N550), .c(N1086), .O(N1473) );
and2 gate237( .a(N1075), .b(N562), .O(N1474) );
and3 gate238( .a(N86), .b(N1075), .c(N1086), .O(N1475) );
and3 gate239( .a(N48), .b(N550), .c(N1086), .O(N1476) );
and3 gate240( .a(N61), .b(N1075), .c(N562), .O(N1477) );
and3 gate241( .a(N85), .b(N1075), .c(N1086), .O(N1478) );
and3 gate242( .a(N47), .b(N550), .c(N1086), .O(N1479) );
and3 gate243( .a(N60), .b(N1075), .c(N562), .O(N1480) );
and3 gate244( .a(N138), .b(N1102), .c(N1113), .O(N1481) );
and3 gate245( .a(N102), .b(N582), .c(N1113), .O(N1482) );
and3 gate246( .a(N126), .b(N1102), .c(N594), .O(N1483) );
and3 gate247( .a(N137), .b(N1102), .c(N1113), .O(N1484) );
and3 gate248( .a(N101), .b(N582), .c(N1113), .O(N1485) );
and3 gate249( .a(N125), .b(N1102), .c(N594), .O(N1486) );
and3 gate250( .a(N136), .b(N1102), .c(N1113), .O(N1487) );
and3 gate251( .a(N100), .b(N582), .c(N1113), .O(N1488) );
and3 gate252( .a(N124), .b(N1102), .c(N594), .O(N1489) );
and3 gate253( .a(N135), .b(N1102), .c(N1113), .O(N1490) );
and3 gate254( .a(N99), .b(N582), .c(N1113), .O(N1491) );
and3 gate255( .a(N123), .b(N1102), .c(N594), .O(N1492) );
and2 gate256( .a(N1102), .b(N1113), .O(N1493) );
and2 gate257( .a(N582), .b(N1113), .O(N1494) );
and2 gate258( .a(N1102), .b(N594), .O(N1495) );
inv1 gate259( .a(N1129), .O(N1496) );
inv1 gate260( .a(N1133), .O(N1499) );

  xor2  gate2390(.a(N1141), .b(N1351), .O(gate261inter0));
  nand2 gate2391(.a(gate261inter0), .b(s_160), .O(gate261inter1));
  and2  gate2392(.a(N1141), .b(N1351), .O(gate261inter2));
  inv1  gate2393(.a(s_160), .O(gate261inter3));
  inv1  gate2394(.a(s_161), .O(gate261inter4));
  nand2 gate2395(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate2396(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate2397(.a(N1351), .O(gate261inter7));
  inv1  gate2398(.a(N1141), .O(gate261inter8));
  nand2 gate2399(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate2400(.a(s_161), .b(gate261inter3), .O(gate261inter10));
  nor2  gate2401(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate2402(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate2403(.a(gate261inter12), .b(gate261inter1), .O(N1502));

  xor2  gate1970(.a(N1353), .b(N1352), .O(gate262inter0));
  nand2 gate1971(.a(gate262inter0), .b(s_100), .O(gate262inter1));
  and2  gate1972(.a(N1353), .b(N1352), .O(gate262inter2));
  inv1  gate1973(.a(s_100), .O(gate262inter3));
  inv1  gate1974(.a(s_101), .O(gate262inter4));
  nand2 gate1975(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate1976(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate1977(.a(N1352), .O(gate262inter7));
  inv1  gate1978(.a(N1353), .O(gate262inter8));
  nand2 gate1979(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate1980(.a(s_101), .b(gate262inter3), .O(gate262inter10));
  nor2  gate1981(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate1982(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate1983(.a(gate262inter12), .b(gate262inter1), .O(N1506));
nand2 gate263( .a(N1354), .b(N1355), .O(N1510) );
buf1 gate264( .a(N1137), .O(N1513) );
buf1 gate265( .a(N1137), .O(N1516) );
inv1 gate266( .a(N1219), .O(N1519) );
inv1 gate267( .a(N1222), .O(N1520) );
inv1 gate268( .a(N1225), .O(N1521) );
inv1 gate269( .a(N1228), .O(N1522) );
inv1 gate270( .a(N1231), .O(N1523) );
inv1 gate271( .a(N1234), .O(N1524) );
inv1 gate272( .a(N1237), .O(N1525) );
inv1 gate273( .a(N1240), .O(N1526) );
inv1 gate274( .a(N1243), .O(N1527) );
inv1 gate275( .a(N1246), .O(N1528) );
and3 gate276( .a(N142), .b(N1146), .c(N1157), .O(N1529) );
and3 gate277( .a(N106), .b(N613), .c(N1157), .O(N1530) );
and3 gate278( .a(N130), .b(N1146), .c(N625), .O(N1531) );
and3 gate279( .a(N131), .b(N1146), .c(N1157), .O(N1532) );
and3 gate280( .a(N95), .b(N613), .c(N1157), .O(N1533) );
and3 gate281( .a(N119), .b(N1146), .c(N625), .O(N1534) );
and3 gate282( .a(N141), .b(N1146), .c(N1157), .O(N1535) );
and3 gate283( .a(N105), .b(N613), .c(N1157), .O(N1536) );
and3 gate284( .a(N129), .b(N1146), .c(N625), .O(N1537) );
and3 gate285( .a(N140), .b(N1146), .c(N1157), .O(N1538) );
and3 gate286( .a(N104), .b(N613), .c(N1157), .O(N1539) );
and3 gate287( .a(N128), .b(N1146), .c(N625), .O(N1540) );
and3 gate288( .a(N139), .b(N1146), .c(N1157), .O(N1541) );
and3 gate289( .a(N103), .b(N613), .c(N1157), .O(N1542) );
and3 gate290( .a(N127), .b(N1146), .c(N625), .O(N1543) );
and2 gate291( .a(N19), .b(N1173), .O(N1544) );
and2 gate292( .a(N4), .b(N1173), .O(N1545) );
and2 gate293( .a(N20), .b(N1173), .O(N1546) );
and2 gate294( .a(N5), .b(N1173), .O(N1547) );
and2 gate295( .a(N21), .b(N1178), .O(N1548) );
and2 gate296( .a(N22), .b(N1178), .O(N1549) );
and2 gate297( .a(N23), .b(N1178), .O(N1550) );
and2 gate298( .a(N6), .b(N1178), .O(N1551) );
and2 gate299( .a(N24), .b(N1178), .O(N1552) );
nand2 gate300( .a(N1395), .b(N1185), .O(N1553) );

  xor2  gate2516(.a(N1397), .b(N1396), .O(gate301inter0));
  nand2 gate2517(.a(gate301inter0), .b(s_178), .O(gate301inter1));
  and2  gate2518(.a(N1397), .b(N1396), .O(gate301inter2));
  inv1  gate2519(.a(s_178), .O(gate301inter3));
  inv1  gate2520(.a(s_179), .O(gate301inter4));
  nand2 gate2521(.a(gate301inter4), .b(gate301inter3), .O(gate301inter5));
  nor2  gate2522(.a(gate301inter5), .b(gate301inter2), .O(gate301inter6));
  inv1  gate2523(.a(N1396), .O(gate301inter7));
  inv1  gate2524(.a(N1397), .O(gate301inter8));
  nand2 gate2525(.a(gate301inter8), .b(gate301inter7), .O(gate301inter9));
  nand2 gate2526(.a(s_179), .b(gate301inter3), .O(gate301inter10));
  nor2  gate2527(.a(gate301inter10), .b(gate301inter9), .O(gate301inter11));
  nor2  gate2528(.a(gate301inter11), .b(gate301inter6), .O(gate301inter12));
  nand2 gate2529(.a(gate301inter12), .b(gate301inter1), .O(N1557));
nand2 gate302( .a(N1398), .b(N1399), .O(N1561) );
and2 gate303( .a(N25), .b(N1200), .O(N1564) );
and2 gate304( .a(N32), .b(N1200), .O(N1565) );
and2 gate305( .a(N26), .b(N1200), .O(N1566) );
and2 gate306( .a(N33), .b(N1200), .O(N1567) );
and2 gate307( .a(N27), .b(N1205), .O(N1568) );
and2 gate308( .a(N34), .b(N1205), .O(N1569) );
and2 gate309( .a(N35), .b(N1205), .O(N1570) );
and2 gate310( .a(N28), .b(N1205), .O(N1571) );
inv1 gate311( .a(N1251), .O(N1572) );
inv1 gate312( .a(N1254), .O(N1573) );
inv1 gate313( .a(N1257), .O(N1574) );
inv1 gate314( .a(N1260), .O(N1575) );
inv1 gate315( .a(N1263), .O(N1576) );
inv1 gate316( .a(N1266), .O(N1577) );

  xor2  gate1816(.a(N1423), .b(N1422), .O(gate317inter0));
  nand2 gate1817(.a(gate317inter0), .b(s_78), .O(gate317inter1));
  and2  gate1818(.a(N1423), .b(N1422), .O(gate317inter2));
  inv1  gate1819(.a(s_78), .O(gate317inter3));
  inv1  gate1820(.a(s_79), .O(gate317inter4));
  nand2 gate1821(.a(gate317inter4), .b(gate317inter3), .O(gate317inter5));
  nor2  gate1822(.a(gate317inter5), .b(gate317inter2), .O(gate317inter6));
  inv1  gate1823(.a(N1422), .O(gate317inter7));
  inv1  gate1824(.a(N1423), .O(gate317inter8));
  nand2 gate1825(.a(gate317inter8), .b(gate317inter7), .O(gate317inter9));
  nand2 gate1826(.a(s_79), .b(gate317inter3), .O(gate317inter10));
  nor2  gate1827(.a(gate317inter10), .b(gate317inter9), .O(gate317inter11));
  nor2  gate1828(.a(gate317inter11), .b(gate317inter6), .O(gate317inter12));
  nand2 gate1829(.a(gate317inter12), .b(gate317inter1), .O(N1578));
inv1 gate318( .a(N1216), .O(N1581) );
nand2 gate319( .a(N1426), .b(N1427), .O(N1582) );

  xor2  gate2978(.a(N1425), .b(N1424), .O(gate320inter0));
  nand2 gate2979(.a(gate320inter0), .b(s_244), .O(gate320inter1));
  and2  gate2980(.a(N1425), .b(N1424), .O(gate320inter2));
  inv1  gate2981(.a(s_244), .O(gate320inter3));
  inv1  gate2982(.a(s_245), .O(gate320inter4));
  nand2 gate2983(.a(gate320inter4), .b(gate320inter3), .O(gate320inter5));
  nor2  gate2984(.a(gate320inter5), .b(gate320inter2), .O(gate320inter6));
  inv1  gate2985(.a(N1424), .O(gate320inter7));
  inv1  gate2986(.a(N1425), .O(gate320inter8));
  nand2 gate2987(.a(gate320inter8), .b(gate320inter7), .O(gate320inter9));
  nand2 gate2988(.a(s_245), .b(gate320inter3), .O(gate320inter10));
  nor2  gate2989(.a(gate320inter10), .b(gate320inter9), .O(gate320inter11));
  nor2  gate2990(.a(gate320inter11), .b(gate320inter6), .O(gate320inter12));
  nand2 gate2991(.a(gate320inter12), .b(gate320inter1), .O(N1585));

  xor2  gate2740(.a(N1441), .b(N1440), .O(gate321inter0));
  nand2 gate2741(.a(gate321inter0), .b(s_210), .O(gate321inter1));
  and2  gate2742(.a(N1441), .b(N1440), .O(gate321inter2));
  inv1  gate2743(.a(s_210), .O(gate321inter3));
  inv1  gate2744(.a(s_211), .O(gate321inter4));
  nand2 gate2745(.a(gate321inter4), .b(gate321inter3), .O(gate321inter5));
  nor2  gate2746(.a(gate321inter5), .b(gate321inter2), .O(gate321inter6));
  inv1  gate2747(.a(N1440), .O(gate321inter7));
  inv1  gate2748(.a(N1441), .O(gate321inter8));
  nand2 gate2749(.a(gate321inter8), .b(gate321inter7), .O(gate321inter9));
  nand2 gate2750(.a(s_211), .b(gate321inter3), .O(gate321inter10));
  nor2  gate2751(.a(gate321inter10), .b(gate321inter9), .O(gate321inter11));
  nor2  gate2752(.a(gate321inter11), .b(gate321inter6), .O(gate321inter12));
  nand2 gate2753(.a(gate321inter12), .b(gate321inter1), .O(N1588));
and2 gate322( .a(N1449), .b(N1450), .O(N1591) );
or4 gate323( .a(N1451), .b(N1452), .c(N1453), .d(N1064), .O(N1596) );
or4 gate324( .a(N1454), .b(N1455), .c(N1456), .d(N1065), .O(N1600) );
or4 gate325( .a(N1457), .b(N1458), .c(N1459), .d(N1066), .O(N1606) );
or4 gate326( .a(N1460), .b(N1461), .c(N1462), .d(N1067), .O(N1612) );
or4 gate327( .a(N1463), .b(N1464), .c(N1465), .d(N1068), .O(N1615) );
or4 gate328( .a(N1466), .b(N1467), .c(N1468), .d(N1097), .O(N1619) );
or4 gate329( .a(N1469), .b(N1470), .c(N1471), .d(N1098), .O(N1624) );
or4 gate330( .a(N1472), .b(N1473), .c(N1474), .d(N1099), .O(N1628) );
or4 gate331( .a(N1475), .b(N1476), .c(N1477), .d(N1100), .O(N1631) );
or4 gate332( .a(N1478), .b(N1479), .c(N1480), .d(N1101), .O(N1634) );
or4 gate333( .a(N1481), .b(N1482), .c(N1483), .d(N1124), .O(N1637) );
or4 gate334( .a(N1484), .b(N1485), .c(N1486), .d(N1125), .O(N1642) );
or4 gate335( .a(N1487), .b(N1488), .c(N1489), .d(N1126), .O(N1647) );
or4 gate336( .a(N1490), .b(N1491), .c(N1492), .d(N1127), .O(N1651) );
or4 gate337( .a(N1493), .b(N1494), .c(N1495), .d(N1128), .O(N1656) );
or4 gate338( .a(N1532), .b(N1533), .c(N1534), .d(N1169), .O(N1676) );
or4 gate339( .a(N1535), .b(N1536), .c(N1537), .d(N1170), .O(N1681) );
or4 gate340( .a(N1538), .b(N1539), .c(N1540), .d(N1171), .O(N1686) );
or4 gate341( .a(N1541), .b(N1542), .c(N1543), .d(N1172), .O(N1690) );
or4 gate342( .a(N1529), .b(N1530), .c(N1531), .d(N1168), .O(N1708) );
buf1 gate343( .a(N1591), .O(N1726) );
inv1 gate344( .a(N1502), .O(N1770) );
inv1 gate345( .a(N1506), .O(N1773) );
inv1 gate346( .a(N1513), .O(N1776) );
inv1 gate347( .a(N1516), .O(N1777) );
buf1 gate348( .a(N1510), .O(N1778) );
buf1 gate349( .a(N1510), .O(N1781) );
and3 gate350( .a(N1133), .b(N1129), .c(N1513), .O(N1784) );
and3 gate351( .a(N1499), .b(N1496), .c(N1516), .O(N1785) );
inv1 gate352( .a(N1553), .O(N1795) );
inv1 gate353( .a(N1557), .O(N1798) );
buf1 gate354( .a(N1561), .O(N1801) );
buf1 gate355( .a(N1561), .O(N1804) );
inv1 gate356( .a(N1588), .O(N1807) );
inv1 gate357( .a(N1578), .O(N1808) );

  xor2  gate1872(.a(N1581), .b(N1578), .O(gate358inter0));
  nand2 gate1873(.a(gate358inter0), .b(s_86), .O(gate358inter1));
  and2  gate1874(.a(N1581), .b(N1578), .O(gate358inter2));
  inv1  gate1875(.a(s_86), .O(gate358inter3));
  inv1  gate1876(.a(s_87), .O(gate358inter4));
  nand2 gate1877(.a(gate358inter4), .b(gate358inter3), .O(gate358inter5));
  nor2  gate1878(.a(gate358inter5), .b(gate358inter2), .O(gate358inter6));
  inv1  gate1879(.a(N1578), .O(gate358inter7));
  inv1  gate1880(.a(N1581), .O(gate358inter8));
  nand2 gate1881(.a(gate358inter8), .b(gate358inter7), .O(gate358inter9));
  nand2 gate1882(.a(s_87), .b(gate358inter3), .O(gate358inter10));
  nor2  gate1883(.a(gate358inter10), .b(gate358inter9), .O(gate358inter11));
  nor2  gate1884(.a(gate358inter11), .b(gate358inter6), .O(gate358inter12));
  nand2 gate1885(.a(gate358inter12), .b(gate358inter1), .O(N1809));
inv1 gate359( .a(N1582), .O(N1810) );
inv1 gate360( .a(N1585), .O(N1811) );
and2 gate361( .a(N1596), .b(N241), .O(N1813) );
and2 gate362( .a(N1606), .b(N241), .O(N1814) );
and2 gate363( .a(N1600), .b(N241), .O(N1815) );
inv1 gate364( .a(N1642), .O(N1816) );
inv1 gate365( .a(N1647), .O(N1817) );
inv1 gate366( .a(N1637), .O(N1818) );
inv1 gate367( .a(N1624), .O(N1819) );
inv1 gate368( .a(N1619), .O(N1820) );
inv1 gate369( .a(N1615), .O(N1821) );
and4 gate370( .a(N496), .b(N224), .c(N36), .d(N1591), .O(N1822) );
and4 gate371( .a(N496), .b(N224), .c(N1591), .d(N486), .O(N1823) );
buf1 gate372( .a(N1596), .O(N1824) );
inv1 gate373( .a(N1606), .O(N1827) );
and2 gate374( .a(N1600), .b(N537), .O(N1830) );
and2 gate375( .a(N1606), .b(N537), .O(N1831) );
and2 gate376( .a(N1619), .b(N246), .O(N1832) );
inv1 gate377( .a(N1596), .O(N1833) );
inv1 gate378( .a(N1600), .O(N1836) );
inv1 gate379( .a(N1606), .O(N1841) );
buf1 gate380( .a(N1612), .O(N1848) );
buf1 gate381( .a(N1615), .O(N1852) );
buf1 gate382( .a(N1619), .O(N1856) );
buf1 gate383( .a(N1624), .O(N1863) );
buf1 gate384( .a(N1628), .O(N1870) );
buf1 gate385( .a(N1631), .O(N1875) );
buf1 gate386( .a(N1634), .O(N1880) );

  xor2  gate3006(.a(N1651), .b(N727), .O(gate387inter0));
  nand2 gate3007(.a(gate387inter0), .b(s_248), .O(gate387inter1));
  and2  gate3008(.a(N1651), .b(N727), .O(gate387inter2));
  inv1  gate3009(.a(s_248), .O(gate387inter3));
  inv1  gate3010(.a(s_249), .O(gate387inter4));
  nand2 gate3011(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate3012(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate3013(.a(N727), .O(gate387inter7));
  inv1  gate3014(.a(N1651), .O(gate387inter8));
  nand2 gate3015(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate3016(.a(s_249), .b(gate387inter3), .O(gate387inter10));
  nor2  gate3017(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate3018(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate3019(.a(gate387inter12), .b(gate387inter1), .O(N1885));
nand2 gate388( .a(N730), .b(N1656), .O(N1888) );
buf1 gate389( .a(N1686), .O(N1891) );
and2 gate390( .a(N1637), .b(N425), .O(N1894) );
inv1 gate391( .a(N1642), .O(N1897) );
and3 gate392( .a(N1496), .b(N1133), .c(N1776), .O(N1908) );
and3 gate393( .a(N1129), .b(N1499), .c(N1777), .O(N1909) );
and2 gate394( .a(N1600), .b(N637), .O(N1910) );
and2 gate395( .a(N1606), .b(N637), .O(N1911) );
and2 gate396( .a(N1612), .b(N637), .O(N1912) );
and2 gate397( .a(N1615), .b(N637), .O(N1913) );
and2 gate398( .a(N1619), .b(N643), .O(N1914) );
and2 gate399( .a(N1624), .b(N643), .O(N1915) );
and2 gate400( .a(N1628), .b(N643), .O(N1916) );
and2 gate401( .a(N1631), .b(N643), .O(N1917) );
and2 gate402( .a(N1634), .b(N643), .O(N1918) );
inv1 gate403( .a(N1708), .O(N1919) );
and2 gate404( .a(N1676), .b(N693), .O(N1928) );
and2 gate405( .a(N1681), .b(N693), .O(N1929) );
and2 gate406( .a(N1686), .b(N693), .O(N1930) );
and2 gate407( .a(N1690), .b(N693), .O(N1931) );
and2 gate408( .a(N1637), .b(N699), .O(N1932) );
and2 gate409( .a(N1642), .b(N699), .O(N1933) );
and2 gate410( .a(N1647), .b(N699), .O(N1934) );
and2 gate411( .a(N1651), .b(N699), .O(N1935) );
buf1 gate412( .a(N1600), .O(N1936) );
nand2 gate413( .a(N1216), .b(N1808), .O(N1939) );
nand2 gate414( .a(N1585), .b(N1810), .O(N1940) );

  xor2  gate2642(.a(N1811), .b(N1582), .O(gate415inter0));
  nand2 gate2643(.a(gate415inter0), .b(s_196), .O(gate415inter1));
  and2  gate2644(.a(N1811), .b(N1582), .O(gate415inter2));
  inv1  gate2645(.a(s_196), .O(gate415inter3));
  inv1  gate2646(.a(s_197), .O(gate415inter4));
  nand2 gate2647(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate2648(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate2649(.a(N1582), .O(gate415inter7));
  inv1  gate2650(.a(N1811), .O(gate415inter8));
  nand2 gate2651(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate2652(.a(s_197), .b(gate415inter3), .O(gate415inter10));
  nor2  gate2653(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate2654(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate2655(.a(gate415inter12), .b(gate415inter1), .O(N1941));
buf1 gate416( .a(N1676), .O(N1942) );
buf1 gate417( .a(N1686), .O(N1945) );
buf1 gate418( .a(N1681), .O(N1948) );
buf1 gate419( .a(N1637), .O(N1951) );
buf1 gate420( .a(N1690), .O(N1954) );
buf1 gate421( .a(N1647), .O(N1957) );
buf1 gate422( .a(N1642), .O(N1960) );
buf1 gate423( .a(N1656), .O(N1963) );
buf1 gate424( .a(N1651), .O(N1966) );
or2 gate425( .a(N533), .b(N1815), .O(N1969) );
inv1 gate426( .a(N1822), .O(N1970) );
inv1 gate427( .a(N1823), .O(N1971) );
buf1 gate428( .a(N1848), .O(N2010) );
buf1 gate429( .a(N1852), .O(N2012) );
buf1 gate430( .a(N1856), .O(N2014) );
buf1 gate431( .a(N1863), .O(N2016) );
buf1 gate432( .a(N1870), .O(N2018) );
buf1 gate433( .a(N1875), .O(N2020) );
buf1 gate434( .a(N1880), .O(N2022) );
inv1 gate435( .a(N1778), .O(N2028) );
inv1 gate436( .a(N1781), .O(N2029) );

  xor2  gate1522(.a(N1784), .b(N1908), .O(gate437inter0));
  nand2 gate1523(.a(gate437inter0), .b(s_36), .O(gate437inter1));
  and2  gate1524(.a(N1784), .b(N1908), .O(gate437inter2));
  inv1  gate1525(.a(s_36), .O(gate437inter3));
  inv1  gate1526(.a(s_37), .O(gate437inter4));
  nand2 gate1527(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate1528(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate1529(.a(N1908), .O(gate437inter7));
  inv1  gate1530(.a(N1784), .O(gate437inter8));
  nand2 gate1531(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate1532(.a(s_37), .b(gate437inter3), .O(gate437inter10));
  nor2  gate1533(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate1534(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate1535(.a(gate437inter12), .b(gate437inter1), .O(N2030));

  xor2  gate2236(.a(N1785), .b(N1909), .O(gate438inter0));
  nand2 gate2237(.a(gate438inter0), .b(s_138), .O(gate438inter1));
  and2  gate2238(.a(N1785), .b(N1909), .O(gate438inter2));
  inv1  gate2239(.a(s_138), .O(gate438inter3));
  inv1  gate2240(.a(s_139), .O(gate438inter4));
  nand2 gate2241(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate2242(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate2243(.a(N1909), .O(gate438inter7));
  inv1  gate2244(.a(N1785), .O(gate438inter8));
  nand2 gate2245(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate2246(.a(s_139), .b(gate438inter3), .O(gate438inter10));
  nor2  gate2247(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate2248(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate2249(.a(gate438inter12), .b(gate438inter1), .O(N2031));
and3 gate439( .a(N1506), .b(N1502), .c(N1778), .O(N2032) );
and3 gate440( .a(N1773), .b(N1770), .c(N1781), .O(N2033) );
or2 gate441( .a(N1571), .b(N1935), .O(N2034) );
inv1 gate442( .a(N1801), .O(N2040) );
inv1 gate443( .a(N1804), .O(N2041) );
and3 gate444( .a(N1557), .b(N1553), .c(N1801), .O(N2042) );
and3 gate445( .a(N1798), .b(N1795), .c(N1804), .O(N2043) );

  xor2  gate2306(.a(N1809), .b(N1939), .O(gate446inter0));
  nand2 gate2307(.a(gate446inter0), .b(s_148), .O(gate446inter1));
  and2  gate2308(.a(N1809), .b(N1939), .O(gate446inter2));
  inv1  gate2309(.a(s_148), .O(gate446inter3));
  inv1  gate2310(.a(s_149), .O(gate446inter4));
  nand2 gate2311(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate2312(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate2313(.a(N1939), .O(gate446inter7));
  inv1  gate2314(.a(N1809), .O(gate446inter8));
  nand2 gate2315(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate2316(.a(s_149), .b(gate446inter3), .O(gate446inter10));
  nor2  gate2317(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate2318(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate2319(.a(gate446inter12), .b(gate446inter1), .O(N2046));
nand2 gate447( .a(N1940), .b(N1941), .O(N2049) );
or2 gate448( .a(N1544), .b(N1910), .O(N2052) );
or2 gate449( .a(N1545), .b(N1911), .O(N2055) );
or2 gate450( .a(N1546), .b(N1912), .O(N2058) );
or2 gate451( .a(N1547), .b(N1913), .O(N2061) );
or2 gate452( .a(N1548), .b(N1914), .O(N2064) );
or2 gate453( .a(N1549), .b(N1915), .O(N2067) );
or2 gate454( .a(N1550), .b(N1916), .O(N2070) );
or2 gate455( .a(N1551), .b(N1917), .O(N2073) );
or2 gate456( .a(N1552), .b(N1918), .O(N2076) );
or2 gate457( .a(N1564), .b(N1928), .O(N2079) );
or2 gate458( .a(N1565), .b(N1929), .O(N2095) );
or2 gate459( .a(N1566), .b(N1930), .O(N2098) );
or2 gate460( .a(N1567), .b(N1931), .O(N2101) );
or2 gate461( .a(N1568), .b(N1932), .O(N2104) );
or2 gate462( .a(N1569), .b(N1933), .O(N2107) );
or2 gate463( .a(N1570), .b(N1934), .O(N2110) );
and3 gate464( .a(N1897), .b(N1894), .c(N40), .O(N2113) );
inv1 gate465( .a(N1894), .O(N2119) );

  xor2  gate2152(.a(N1827), .b(N408), .O(gate466inter0));
  nand2 gate2153(.a(gate466inter0), .b(s_126), .O(gate466inter1));
  and2  gate2154(.a(N1827), .b(N408), .O(gate466inter2));
  inv1  gate2155(.a(s_126), .O(gate466inter3));
  inv1  gate2156(.a(s_127), .O(gate466inter4));
  nand2 gate2157(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate2158(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate2159(.a(N408), .O(gate466inter7));
  inv1  gate2160(.a(N1827), .O(gate466inter8));
  nand2 gate2161(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate2162(.a(s_127), .b(gate466inter3), .O(gate466inter10));
  nor2  gate2163(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate2164(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate2165(.a(gate466inter12), .b(gate466inter1), .O(N2120));
and2 gate467( .a(N1824), .b(N537), .O(N2125) );
and2 gate468( .a(N1852), .b(N246), .O(N2126) );
and2 gate469( .a(N1848), .b(N537), .O(N2127) );
inv1 gate470( .a(N1848), .O(N2128) );
inv1 gate471( .a(N1852), .O(N2135) );
inv1 gate472( .a(N1863), .O(N2141) );
inv1 gate473( .a(N1870), .O(N2144) );
inv1 gate474( .a(N1875), .O(N2147) );
inv1 gate475( .a(N1880), .O(N2150) );
and2 gate476( .a(N727), .b(N1885), .O(N2153) );
and2 gate477( .a(N1885), .b(N1651), .O(N2154) );
and2 gate478( .a(N730), .b(N1888), .O(N2155) );
and2 gate479( .a(N1888), .b(N1656), .O(N2156) );
and3 gate480( .a(N1770), .b(N1506), .c(N2028), .O(N2157) );
and3 gate481( .a(N1502), .b(N1773), .c(N2029), .O(N2158) );
inv1 gate482( .a(N1942), .O(N2171) );
nand2 gate483( .a(N1942), .b(N1919), .O(N2172) );
inv1 gate484( .a(N1945), .O(N2173) );
inv1 gate485( .a(N1948), .O(N2174) );
inv1 gate486( .a(N1951), .O(N2175) );
inv1 gate487( .a(N1954), .O(N2176) );
and3 gate488( .a(N1795), .b(N1557), .c(N2040), .O(N2177) );
and3 gate489( .a(N1553), .b(N1798), .c(N2041), .O(N2178) );
buf1 gate490( .a(N1836), .O(N2185) );
buf1 gate491( .a(N1833), .O(N2188) );
buf1 gate492( .a(N1841), .O(N2191) );
inv1 gate493( .a(N1856), .O(N2194) );
inv1 gate494( .a(N1827), .O(N2197) );
inv1 gate495( .a(N1936), .O(N2200) );
buf1 gate496( .a(N1836), .O(N2201) );
buf1 gate497( .a(N1833), .O(N2204) );
buf1 gate498( .a(N1841), .O(N2207) );
buf1 gate499( .a(N1824), .O(N2210) );
buf1 gate500( .a(N1841), .O(N2213) );
buf1 gate501( .a(N1841), .O(N2216) );
nand2 gate502( .a(N2031), .b(N2030), .O(N2219) );
inv1 gate503( .a(N1957), .O(N2234) );
inv1 gate504( .a(N1960), .O(N2235) );
inv1 gate505( .a(N1963), .O(N2236) );
inv1 gate506( .a(N1966), .O(N2237) );
and3 gate507( .a(N40), .b(N1897), .c(N2119), .O(N2250) );
or2 gate508( .a(N1831), .b(N2126), .O(N2266) );
or2 gate509( .a(N2127), .b(N1832), .O(N2269) );
or2 gate510( .a(N2153), .b(N2154), .O(N2291) );
or2 gate511( .a(N2155), .b(N2156), .O(N2294) );

  xor2  gate2796(.a(N2032), .b(N2157), .O(gate512inter0));
  nand2 gate2797(.a(gate512inter0), .b(s_218), .O(gate512inter1));
  and2  gate2798(.a(N2032), .b(N2157), .O(gate512inter2));
  inv1  gate2799(.a(s_218), .O(gate512inter3));
  inv1  gate2800(.a(s_219), .O(gate512inter4));
  nand2 gate2801(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate2802(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate2803(.a(N2157), .O(gate512inter7));
  inv1  gate2804(.a(N2032), .O(gate512inter8));
  nand2 gate2805(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate2806(.a(s_219), .b(gate512inter3), .O(gate512inter10));
  nor2  gate2807(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate2808(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate2809(.a(gate512inter12), .b(gate512inter1), .O(N2297));

  xor2  gate2992(.a(N2033), .b(N2158), .O(gate513inter0));
  nand2 gate2993(.a(gate513inter0), .b(s_246), .O(gate513inter1));
  and2  gate2994(.a(N2033), .b(N2158), .O(gate513inter2));
  inv1  gate2995(.a(s_246), .O(gate513inter3));
  inv1  gate2996(.a(s_247), .O(gate513inter4));
  nand2 gate2997(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate2998(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate2999(.a(N2158), .O(gate513inter7));
  inv1  gate3000(.a(N2033), .O(gate513inter8));
  nand2 gate3001(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate3002(.a(s_247), .b(gate513inter3), .O(gate513inter10));
  nor2  gate3003(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate3004(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate3005(.a(gate513inter12), .b(gate513inter1), .O(N2298));
inv1 gate514( .a(N2046), .O(N2300) );
inv1 gate515( .a(N2049), .O(N2301) );
nand2 gate516( .a(N2052), .b(N1519), .O(N2302) );
inv1 gate517( .a(N2052), .O(N2303) );

  xor2  gate2208(.a(N1520), .b(N2055), .O(gate518inter0));
  nand2 gate2209(.a(gate518inter0), .b(s_134), .O(gate518inter1));
  and2  gate2210(.a(N1520), .b(N2055), .O(gate518inter2));
  inv1  gate2211(.a(s_134), .O(gate518inter3));
  inv1  gate2212(.a(s_135), .O(gate518inter4));
  nand2 gate2213(.a(gate518inter4), .b(gate518inter3), .O(gate518inter5));
  nor2  gate2214(.a(gate518inter5), .b(gate518inter2), .O(gate518inter6));
  inv1  gate2215(.a(N2055), .O(gate518inter7));
  inv1  gate2216(.a(N1520), .O(gate518inter8));
  nand2 gate2217(.a(gate518inter8), .b(gate518inter7), .O(gate518inter9));
  nand2 gate2218(.a(s_135), .b(gate518inter3), .O(gate518inter10));
  nor2  gate2219(.a(gate518inter10), .b(gate518inter9), .O(gate518inter11));
  nor2  gate2220(.a(gate518inter11), .b(gate518inter6), .O(gate518inter12));
  nand2 gate2221(.a(gate518inter12), .b(gate518inter1), .O(N2304));
inv1 gate519( .a(N2055), .O(N2305) );

  xor2  gate1620(.a(N1521), .b(N2058), .O(gate520inter0));
  nand2 gate1621(.a(gate520inter0), .b(s_50), .O(gate520inter1));
  and2  gate1622(.a(N1521), .b(N2058), .O(gate520inter2));
  inv1  gate1623(.a(s_50), .O(gate520inter3));
  inv1  gate1624(.a(s_51), .O(gate520inter4));
  nand2 gate1625(.a(gate520inter4), .b(gate520inter3), .O(gate520inter5));
  nor2  gate1626(.a(gate520inter5), .b(gate520inter2), .O(gate520inter6));
  inv1  gate1627(.a(N2058), .O(gate520inter7));
  inv1  gate1628(.a(N1521), .O(gate520inter8));
  nand2 gate1629(.a(gate520inter8), .b(gate520inter7), .O(gate520inter9));
  nand2 gate1630(.a(s_51), .b(gate520inter3), .O(gate520inter10));
  nor2  gate1631(.a(gate520inter10), .b(gate520inter9), .O(gate520inter11));
  nor2  gate1632(.a(gate520inter11), .b(gate520inter6), .O(gate520inter12));
  nand2 gate1633(.a(gate520inter12), .b(gate520inter1), .O(N2306));
inv1 gate521( .a(N2058), .O(N2307) );

  xor2  gate2292(.a(N1522), .b(N2061), .O(gate522inter0));
  nand2 gate2293(.a(gate522inter0), .b(s_146), .O(gate522inter1));
  and2  gate2294(.a(N1522), .b(N2061), .O(gate522inter2));
  inv1  gate2295(.a(s_146), .O(gate522inter3));
  inv1  gate2296(.a(s_147), .O(gate522inter4));
  nand2 gate2297(.a(gate522inter4), .b(gate522inter3), .O(gate522inter5));
  nor2  gate2298(.a(gate522inter5), .b(gate522inter2), .O(gate522inter6));
  inv1  gate2299(.a(N2061), .O(gate522inter7));
  inv1  gate2300(.a(N1522), .O(gate522inter8));
  nand2 gate2301(.a(gate522inter8), .b(gate522inter7), .O(gate522inter9));
  nand2 gate2302(.a(s_147), .b(gate522inter3), .O(gate522inter10));
  nor2  gate2303(.a(gate522inter10), .b(gate522inter9), .O(gate522inter11));
  nor2  gate2304(.a(gate522inter11), .b(gate522inter6), .O(gate522inter12));
  nand2 gate2305(.a(gate522inter12), .b(gate522inter1), .O(N2308));
inv1 gate523( .a(N2061), .O(N2309) );

  xor2  gate2698(.a(N1523), .b(N2064), .O(gate524inter0));
  nand2 gate2699(.a(gate524inter0), .b(s_204), .O(gate524inter1));
  and2  gate2700(.a(N1523), .b(N2064), .O(gate524inter2));
  inv1  gate2701(.a(s_204), .O(gate524inter3));
  inv1  gate2702(.a(s_205), .O(gate524inter4));
  nand2 gate2703(.a(gate524inter4), .b(gate524inter3), .O(gate524inter5));
  nor2  gate2704(.a(gate524inter5), .b(gate524inter2), .O(gate524inter6));
  inv1  gate2705(.a(N2064), .O(gate524inter7));
  inv1  gate2706(.a(N1523), .O(gate524inter8));
  nand2 gate2707(.a(gate524inter8), .b(gate524inter7), .O(gate524inter9));
  nand2 gate2708(.a(s_205), .b(gate524inter3), .O(gate524inter10));
  nor2  gate2709(.a(gate524inter10), .b(gate524inter9), .O(gate524inter11));
  nor2  gate2710(.a(gate524inter11), .b(gate524inter6), .O(gate524inter12));
  nand2 gate2711(.a(gate524inter12), .b(gate524inter1), .O(N2310));
inv1 gate525( .a(N2064), .O(N2311) );

  xor2  gate1284(.a(N1524), .b(N2067), .O(gate526inter0));
  nand2 gate1285(.a(gate526inter0), .b(s_2), .O(gate526inter1));
  and2  gate1286(.a(N1524), .b(N2067), .O(gate526inter2));
  inv1  gate1287(.a(s_2), .O(gate526inter3));
  inv1  gate1288(.a(s_3), .O(gate526inter4));
  nand2 gate1289(.a(gate526inter4), .b(gate526inter3), .O(gate526inter5));
  nor2  gate1290(.a(gate526inter5), .b(gate526inter2), .O(gate526inter6));
  inv1  gate1291(.a(N2067), .O(gate526inter7));
  inv1  gate1292(.a(N1524), .O(gate526inter8));
  nand2 gate1293(.a(gate526inter8), .b(gate526inter7), .O(gate526inter9));
  nand2 gate1294(.a(s_3), .b(gate526inter3), .O(gate526inter10));
  nor2  gate1295(.a(gate526inter10), .b(gate526inter9), .O(gate526inter11));
  nor2  gate1296(.a(gate526inter11), .b(gate526inter6), .O(gate526inter12));
  nand2 gate1297(.a(gate526inter12), .b(gate526inter1), .O(N2312));
inv1 gate527( .a(N2067), .O(N2313) );
nand2 gate528( .a(N2070), .b(N1525), .O(N2314) );
inv1 gate529( .a(N2070), .O(N2315) );

  xor2  gate2852(.a(N1526), .b(N2073), .O(gate530inter0));
  nand2 gate2853(.a(gate530inter0), .b(s_226), .O(gate530inter1));
  and2  gate2854(.a(N1526), .b(N2073), .O(gate530inter2));
  inv1  gate2855(.a(s_226), .O(gate530inter3));
  inv1  gate2856(.a(s_227), .O(gate530inter4));
  nand2 gate2857(.a(gate530inter4), .b(gate530inter3), .O(gate530inter5));
  nor2  gate2858(.a(gate530inter5), .b(gate530inter2), .O(gate530inter6));
  inv1  gate2859(.a(N2073), .O(gate530inter7));
  inv1  gate2860(.a(N1526), .O(gate530inter8));
  nand2 gate2861(.a(gate530inter8), .b(gate530inter7), .O(gate530inter9));
  nand2 gate2862(.a(s_227), .b(gate530inter3), .O(gate530inter10));
  nor2  gate2863(.a(gate530inter10), .b(gate530inter9), .O(gate530inter11));
  nor2  gate2864(.a(gate530inter11), .b(gate530inter6), .O(gate530inter12));
  nand2 gate2865(.a(gate530inter12), .b(gate530inter1), .O(N2316));
inv1 gate531( .a(N2073), .O(N2317) );
nand2 gate532( .a(N2076), .b(N1527), .O(N2318) );
inv1 gate533( .a(N2076), .O(N2319) );

  xor2  gate2194(.a(N1528), .b(N2079), .O(gate534inter0));
  nand2 gate2195(.a(gate534inter0), .b(s_132), .O(gate534inter1));
  and2  gate2196(.a(N1528), .b(N2079), .O(gate534inter2));
  inv1  gate2197(.a(s_132), .O(gate534inter3));
  inv1  gate2198(.a(s_133), .O(gate534inter4));
  nand2 gate2199(.a(gate534inter4), .b(gate534inter3), .O(gate534inter5));
  nor2  gate2200(.a(gate534inter5), .b(gate534inter2), .O(gate534inter6));
  inv1  gate2201(.a(N2079), .O(gate534inter7));
  inv1  gate2202(.a(N1528), .O(gate534inter8));
  nand2 gate2203(.a(gate534inter8), .b(gate534inter7), .O(gate534inter9));
  nand2 gate2204(.a(s_133), .b(gate534inter3), .O(gate534inter10));
  nor2  gate2205(.a(gate534inter10), .b(gate534inter9), .O(gate534inter11));
  nor2  gate2206(.a(gate534inter11), .b(gate534inter6), .O(gate534inter12));
  nand2 gate2207(.a(gate534inter12), .b(gate534inter1), .O(N2320));
inv1 gate535( .a(N2079), .O(N2321) );
nand2 gate536( .a(N1708), .b(N2171), .O(N2322) );

  xor2  gate2348(.a(N2173), .b(N1948), .O(gate537inter0));
  nand2 gate2349(.a(gate537inter0), .b(s_154), .O(gate537inter1));
  and2  gate2350(.a(N2173), .b(N1948), .O(gate537inter2));
  inv1  gate2351(.a(s_154), .O(gate537inter3));
  inv1  gate2352(.a(s_155), .O(gate537inter4));
  nand2 gate2353(.a(gate537inter4), .b(gate537inter3), .O(gate537inter5));
  nor2  gate2354(.a(gate537inter5), .b(gate537inter2), .O(gate537inter6));
  inv1  gate2355(.a(N1948), .O(gate537inter7));
  inv1  gate2356(.a(N2173), .O(gate537inter8));
  nand2 gate2357(.a(gate537inter8), .b(gate537inter7), .O(gate537inter9));
  nand2 gate2358(.a(s_155), .b(gate537inter3), .O(gate537inter10));
  nor2  gate2359(.a(gate537inter10), .b(gate537inter9), .O(gate537inter11));
  nor2  gate2360(.a(gate537inter11), .b(gate537inter6), .O(gate537inter12));
  nand2 gate2361(.a(gate537inter12), .b(gate537inter1), .O(N2323));
nand2 gate538( .a(N1945), .b(N2174), .O(N2324) );
nand2 gate539( .a(N1954), .b(N2175), .O(N2325) );
nand2 gate540( .a(N1951), .b(N2176), .O(N2326) );
nor2 gate541( .a(N2177), .b(N2042), .O(N2327) );
nor2 gate542( .a(N2178), .b(N2043), .O(N2328) );
nand2 gate543( .a(N2095), .b(N1572), .O(N2329) );
inv1 gate544( .a(N2095), .O(N2330) );

  xor2  gate1802(.a(N1573), .b(N2098), .O(gate545inter0));
  nand2 gate1803(.a(gate545inter0), .b(s_76), .O(gate545inter1));
  and2  gate1804(.a(N1573), .b(N2098), .O(gate545inter2));
  inv1  gate1805(.a(s_76), .O(gate545inter3));
  inv1  gate1806(.a(s_77), .O(gate545inter4));
  nand2 gate1807(.a(gate545inter4), .b(gate545inter3), .O(gate545inter5));
  nor2  gate1808(.a(gate545inter5), .b(gate545inter2), .O(gate545inter6));
  inv1  gate1809(.a(N2098), .O(gate545inter7));
  inv1  gate1810(.a(N1573), .O(gate545inter8));
  nand2 gate1811(.a(gate545inter8), .b(gate545inter7), .O(gate545inter9));
  nand2 gate1812(.a(s_77), .b(gate545inter3), .O(gate545inter10));
  nor2  gate1813(.a(gate545inter10), .b(gate545inter9), .O(gate545inter11));
  nor2  gate1814(.a(gate545inter11), .b(gate545inter6), .O(gate545inter12));
  nand2 gate1815(.a(gate545inter12), .b(gate545inter1), .O(N2331));
inv1 gate546( .a(N2098), .O(N2332) );
nand2 gate547( .a(N2101), .b(N1574), .O(N2333) );
inv1 gate548( .a(N2101), .O(N2334) );
nand2 gate549( .a(N2104), .b(N1575), .O(N2335) );
inv1 gate550( .a(N2104), .O(N2336) );

  xor2  gate1914(.a(N1576), .b(N2107), .O(gate551inter0));
  nand2 gate1915(.a(gate551inter0), .b(s_92), .O(gate551inter1));
  and2  gate1916(.a(N1576), .b(N2107), .O(gate551inter2));
  inv1  gate1917(.a(s_92), .O(gate551inter3));
  inv1  gate1918(.a(s_93), .O(gate551inter4));
  nand2 gate1919(.a(gate551inter4), .b(gate551inter3), .O(gate551inter5));
  nor2  gate1920(.a(gate551inter5), .b(gate551inter2), .O(gate551inter6));
  inv1  gate1921(.a(N2107), .O(gate551inter7));
  inv1  gate1922(.a(N1576), .O(gate551inter8));
  nand2 gate1923(.a(gate551inter8), .b(gate551inter7), .O(gate551inter9));
  nand2 gate1924(.a(s_93), .b(gate551inter3), .O(gate551inter10));
  nor2  gate1925(.a(gate551inter10), .b(gate551inter9), .O(gate551inter11));
  nor2  gate1926(.a(gate551inter11), .b(gate551inter6), .O(gate551inter12));
  nand2 gate1927(.a(gate551inter12), .b(gate551inter1), .O(N2337));
inv1 gate552( .a(N2107), .O(N2338) );
nand2 gate553( .a(N2110), .b(N1577), .O(N2339) );
inv1 gate554( .a(N2110), .O(N2340) );
nand2 gate555( .a(N1960), .b(N2234), .O(N2354) );

  xor2  gate2824(.a(N2235), .b(N1957), .O(gate556inter0));
  nand2 gate2825(.a(gate556inter0), .b(s_222), .O(gate556inter1));
  and2  gate2826(.a(N2235), .b(N1957), .O(gate556inter2));
  inv1  gate2827(.a(s_222), .O(gate556inter3));
  inv1  gate2828(.a(s_223), .O(gate556inter4));
  nand2 gate2829(.a(gate556inter4), .b(gate556inter3), .O(gate556inter5));
  nor2  gate2830(.a(gate556inter5), .b(gate556inter2), .O(gate556inter6));
  inv1  gate2831(.a(N1957), .O(gate556inter7));
  inv1  gate2832(.a(N2235), .O(gate556inter8));
  nand2 gate2833(.a(gate556inter8), .b(gate556inter7), .O(gate556inter9));
  nand2 gate2834(.a(s_223), .b(gate556inter3), .O(gate556inter10));
  nor2  gate2835(.a(gate556inter10), .b(gate556inter9), .O(gate556inter11));
  nor2  gate2836(.a(gate556inter11), .b(gate556inter6), .O(gate556inter12));
  nand2 gate2837(.a(gate556inter12), .b(gate556inter1), .O(N2355));

  xor2  gate2670(.a(N2236), .b(N1966), .O(gate557inter0));
  nand2 gate2671(.a(gate557inter0), .b(s_200), .O(gate557inter1));
  and2  gate2672(.a(N2236), .b(N1966), .O(gate557inter2));
  inv1  gate2673(.a(s_200), .O(gate557inter3));
  inv1  gate2674(.a(s_201), .O(gate557inter4));
  nand2 gate2675(.a(gate557inter4), .b(gate557inter3), .O(gate557inter5));
  nor2  gate2676(.a(gate557inter5), .b(gate557inter2), .O(gate557inter6));
  inv1  gate2677(.a(N1966), .O(gate557inter7));
  inv1  gate2678(.a(N2236), .O(gate557inter8));
  nand2 gate2679(.a(gate557inter8), .b(gate557inter7), .O(gate557inter9));
  nand2 gate2680(.a(s_201), .b(gate557inter3), .O(gate557inter10));
  nor2  gate2681(.a(gate557inter10), .b(gate557inter9), .O(gate557inter11));
  nor2  gate2682(.a(gate557inter11), .b(gate557inter6), .O(gate557inter12));
  nand2 gate2683(.a(gate557inter12), .b(gate557inter1), .O(N2356));
nand2 gate558( .a(N1963), .b(N2237), .O(N2357) );
and2 gate559( .a(N2120), .b(N533), .O(N2358) );
inv1 gate560( .a(N2113), .O(N2359) );
inv1 gate561( .a(N2185), .O(N2364) );
inv1 gate562( .a(N2188), .O(N2365) );
inv1 gate563( .a(N2191), .O(N2366) );
inv1 gate564( .a(N2194), .O(N2367) );
buf1 gate565( .a(N2120), .O(N2368) );
inv1 gate566( .a(N2201), .O(N2372) );
inv1 gate567( .a(N2204), .O(N2373) );
inv1 gate568( .a(N2207), .O(N2374) );
inv1 gate569( .a(N2210), .O(N2375) );
inv1 gate570( .a(N2213), .O(N2376) );
inv1 gate571( .a(N2113), .O(N2377) );
buf1 gate572( .a(N2113), .O(N2382) );
and2 gate573( .a(N2120), .b(N246), .O(N2386) );
buf1 gate574( .a(N2266), .O(N2387) );
buf1 gate575( .a(N2266), .O(N2388) );
buf1 gate576( .a(N2269), .O(N2389) );
buf1 gate577( .a(N2269), .O(N2390) );
buf1 gate578( .a(N2113), .O(N2391) );
inv1 gate579( .a(N2113), .O(N2395) );
nand2 gate580( .a(N2219), .b(N2300), .O(N2400) );
inv1 gate581( .a(N2216), .O(N2403) );
inv1 gate582( .a(N2219), .O(N2406) );
nand2 gate583( .a(N1219), .b(N2303), .O(N2407) );

  xor2  gate2068(.a(N2305), .b(N1222), .O(gate584inter0));
  nand2 gate2069(.a(gate584inter0), .b(s_114), .O(gate584inter1));
  and2  gate2070(.a(N2305), .b(N1222), .O(gate584inter2));
  inv1  gate2071(.a(s_114), .O(gate584inter3));
  inv1  gate2072(.a(s_115), .O(gate584inter4));
  nand2 gate2073(.a(gate584inter4), .b(gate584inter3), .O(gate584inter5));
  nor2  gate2074(.a(gate584inter5), .b(gate584inter2), .O(gate584inter6));
  inv1  gate2075(.a(N1222), .O(gate584inter7));
  inv1  gate2076(.a(N2305), .O(gate584inter8));
  nand2 gate2077(.a(gate584inter8), .b(gate584inter7), .O(gate584inter9));
  nand2 gate2078(.a(s_115), .b(gate584inter3), .O(gate584inter10));
  nor2  gate2079(.a(gate584inter10), .b(gate584inter9), .O(gate584inter11));
  nor2  gate2080(.a(gate584inter11), .b(gate584inter6), .O(gate584inter12));
  nand2 gate2081(.a(gate584inter12), .b(gate584inter1), .O(N2408));
nand2 gate585( .a(N1225), .b(N2307), .O(N2409) );

  xor2  gate1368(.a(N2309), .b(N1228), .O(gate586inter0));
  nand2 gate1369(.a(gate586inter0), .b(s_14), .O(gate586inter1));
  and2  gate1370(.a(N2309), .b(N1228), .O(gate586inter2));
  inv1  gate1371(.a(s_14), .O(gate586inter3));
  inv1  gate1372(.a(s_15), .O(gate586inter4));
  nand2 gate1373(.a(gate586inter4), .b(gate586inter3), .O(gate586inter5));
  nor2  gate1374(.a(gate586inter5), .b(gate586inter2), .O(gate586inter6));
  inv1  gate1375(.a(N1228), .O(gate586inter7));
  inv1  gate1376(.a(N2309), .O(gate586inter8));
  nand2 gate1377(.a(gate586inter8), .b(gate586inter7), .O(gate586inter9));
  nand2 gate1378(.a(s_15), .b(gate586inter3), .O(gate586inter10));
  nor2  gate1379(.a(gate586inter10), .b(gate586inter9), .O(gate586inter11));
  nor2  gate1380(.a(gate586inter11), .b(gate586inter6), .O(gate586inter12));
  nand2 gate1381(.a(gate586inter12), .b(gate586inter1), .O(N2410));

  xor2  gate1774(.a(N2311), .b(N1231), .O(gate587inter0));
  nand2 gate1775(.a(gate587inter0), .b(s_72), .O(gate587inter1));
  and2  gate1776(.a(N2311), .b(N1231), .O(gate587inter2));
  inv1  gate1777(.a(s_72), .O(gate587inter3));
  inv1  gate1778(.a(s_73), .O(gate587inter4));
  nand2 gate1779(.a(gate587inter4), .b(gate587inter3), .O(gate587inter5));
  nor2  gate1780(.a(gate587inter5), .b(gate587inter2), .O(gate587inter6));
  inv1  gate1781(.a(N1231), .O(gate587inter7));
  inv1  gate1782(.a(N2311), .O(gate587inter8));
  nand2 gate1783(.a(gate587inter8), .b(gate587inter7), .O(gate587inter9));
  nand2 gate1784(.a(s_73), .b(gate587inter3), .O(gate587inter10));
  nor2  gate1785(.a(gate587inter10), .b(gate587inter9), .O(gate587inter11));
  nor2  gate1786(.a(gate587inter11), .b(gate587inter6), .O(gate587inter12));
  nand2 gate1787(.a(gate587inter12), .b(gate587inter1), .O(N2411));
nand2 gate588( .a(N1234), .b(N2313), .O(N2412) );
nand2 gate589( .a(N1237), .b(N2315), .O(N2413) );

  xor2  gate1732(.a(N2317), .b(N1240), .O(gate590inter0));
  nand2 gate1733(.a(gate590inter0), .b(s_66), .O(gate590inter1));
  and2  gate1734(.a(N2317), .b(N1240), .O(gate590inter2));
  inv1  gate1735(.a(s_66), .O(gate590inter3));
  inv1  gate1736(.a(s_67), .O(gate590inter4));
  nand2 gate1737(.a(gate590inter4), .b(gate590inter3), .O(gate590inter5));
  nor2  gate1738(.a(gate590inter5), .b(gate590inter2), .O(gate590inter6));
  inv1  gate1739(.a(N1240), .O(gate590inter7));
  inv1  gate1740(.a(N2317), .O(gate590inter8));
  nand2 gate1741(.a(gate590inter8), .b(gate590inter7), .O(gate590inter9));
  nand2 gate1742(.a(s_67), .b(gate590inter3), .O(gate590inter10));
  nor2  gate1743(.a(gate590inter10), .b(gate590inter9), .O(gate590inter11));
  nor2  gate1744(.a(gate590inter11), .b(gate590inter6), .O(gate590inter12));
  nand2 gate1745(.a(gate590inter12), .b(gate590inter1), .O(N2414));

  xor2  gate1956(.a(N2319), .b(N1243), .O(gate591inter0));
  nand2 gate1957(.a(gate591inter0), .b(s_98), .O(gate591inter1));
  and2  gate1958(.a(N2319), .b(N1243), .O(gate591inter2));
  inv1  gate1959(.a(s_98), .O(gate591inter3));
  inv1  gate1960(.a(s_99), .O(gate591inter4));
  nand2 gate1961(.a(gate591inter4), .b(gate591inter3), .O(gate591inter5));
  nor2  gate1962(.a(gate591inter5), .b(gate591inter2), .O(gate591inter6));
  inv1  gate1963(.a(N1243), .O(gate591inter7));
  inv1  gate1964(.a(N2319), .O(gate591inter8));
  nand2 gate1965(.a(gate591inter8), .b(gate591inter7), .O(gate591inter9));
  nand2 gate1966(.a(s_99), .b(gate591inter3), .O(gate591inter10));
  nor2  gate1967(.a(gate591inter10), .b(gate591inter9), .O(gate591inter11));
  nor2  gate1968(.a(gate591inter11), .b(gate591inter6), .O(gate591inter12));
  nand2 gate1969(.a(gate591inter12), .b(gate591inter1), .O(N2415));
nand2 gate592( .a(N1246), .b(N2321), .O(N2416) );
nand2 gate593( .a(N2322), .b(N2172), .O(N2417) );

  xor2  gate1564(.a(N2324), .b(N2323), .O(gate594inter0));
  nand2 gate1565(.a(gate594inter0), .b(s_42), .O(gate594inter1));
  and2  gate1566(.a(N2324), .b(N2323), .O(gate594inter2));
  inv1  gate1567(.a(s_42), .O(gate594inter3));
  inv1  gate1568(.a(s_43), .O(gate594inter4));
  nand2 gate1569(.a(gate594inter4), .b(gate594inter3), .O(gate594inter5));
  nor2  gate1570(.a(gate594inter5), .b(gate594inter2), .O(gate594inter6));
  inv1  gate1571(.a(N2323), .O(gate594inter7));
  inv1  gate1572(.a(N2324), .O(gate594inter8));
  nand2 gate1573(.a(gate594inter8), .b(gate594inter7), .O(gate594inter9));
  nand2 gate1574(.a(s_43), .b(gate594inter3), .O(gate594inter10));
  nor2  gate1575(.a(gate594inter10), .b(gate594inter9), .O(gate594inter11));
  nor2  gate1576(.a(gate594inter11), .b(gate594inter6), .O(gate594inter12));
  nand2 gate1577(.a(gate594inter12), .b(gate594inter1), .O(N2421));

  xor2  gate2124(.a(N2326), .b(N2325), .O(gate595inter0));
  nand2 gate2125(.a(gate595inter0), .b(s_122), .O(gate595inter1));
  and2  gate2126(.a(N2326), .b(N2325), .O(gate595inter2));
  inv1  gate2127(.a(s_122), .O(gate595inter3));
  inv1  gate2128(.a(s_123), .O(gate595inter4));
  nand2 gate2129(.a(gate595inter4), .b(gate595inter3), .O(gate595inter5));
  nor2  gate2130(.a(gate595inter5), .b(gate595inter2), .O(gate595inter6));
  inv1  gate2131(.a(N2325), .O(gate595inter7));
  inv1  gate2132(.a(N2326), .O(gate595inter8));
  nand2 gate2133(.a(gate595inter8), .b(gate595inter7), .O(gate595inter9));
  nand2 gate2134(.a(s_123), .b(gate595inter3), .O(gate595inter10));
  nor2  gate2135(.a(gate595inter10), .b(gate595inter9), .O(gate595inter11));
  nor2  gate2136(.a(gate595inter11), .b(gate595inter6), .O(gate595inter12));
  nand2 gate2137(.a(gate595inter12), .b(gate595inter1), .O(N2425));
nand2 gate596( .a(N1251), .b(N2330), .O(N2428) );
nand2 gate597( .a(N1254), .b(N2332), .O(N2429) );

  xor2  gate1410(.a(N2334), .b(N1257), .O(gate598inter0));
  nand2 gate1411(.a(gate598inter0), .b(s_20), .O(gate598inter1));
  and2  gate1412(.a(N2334), .b(N1257), .O(gate598inter2));
  inv1  gate1413(.a(s_20), .O(gate598inter3));
  inv1  gate1414(.a(s_21), .O(gate598inter4));
  nand2 gate1415(.a(gate598inter4), .b(gate598inter3), .O(gate598inter5));
  nor2  gate1416(.a(gate598inter5), .b(gate598inter2), .O(gate598inter6));
  inv1  gate1417(.a(N1257), .O(gate598inter7));
  inv1  gate1418(.a(N2334), .O(gate598inter8));
  nand2 gate1419(.a(gate598inter8), .b(gate598inter7), .O(gate598inter9));
  nand2 gate1420(.a(s_21), .b(gate598inter3), .O(gate598inter10));
  nor2  gate1421(.a(gate598inter10), .b(gate598inter9), .O(gate598inter11));
  nor2  gate1422(.a(gate598inter11), .b(gate598inter6), .O(gate598inter12));
  nand2 gate1423(.a(gate598inter12), .b(gate598inter1), .O(N2430));
nand2 gate599( .a(N1260), .b(N2336), .O(N2431) );
nand2 gate600( .a(N1263), .b(N2338), .O(N2432) );

  xor2  gate2572(.a(N2340), .b(N1266), .O(gate601inter0));
  nand2 gate2573(.a(gate601inter0), .b(s_186), .O(gate601inter1));
  and2  gate2574(.a(N2340), .b(N1266), .O(gate601inter2));
  inv1  gate2575(.a(s_186), .O(gate601inter3));
  inv1  gate2576(.a(s_187), .O(gate601inter4));
  nand2 gate2577(.a(gate601inter4), .b(gate601inter3), .O(gate601inter5));
  nor2  gate2578(.a(gate601inter5), .b(gate601inter2), .O(gate601inter6));
  inv1  gate2579(.a(N1266), .O(gate601inter7));
  inv1  gate2580(.a(N2340), .O(gate601inter8));
  nand2 gate2581(.a(gate601inter8), .b(gate601inter7), .O(gate601inter9));
  nand2 gate2582(.a(s_187), .b(gate601inter3), .O(gate601inter10));
  nor2  gate2583(.a(gate601inter10), .b(gate601inter9), .O(gate601inter11));
  nor2  gate2584(.a(gate601inter11), .b(gate601inter6), .O(gate601inter12));
  nand2 gate2585(.a(gate601inter12), .b(gate601inter1), .O(N2433));
buf1 gate602( .a(N2128), .O(N2434) );
buf1 gate603( .a(N2135), .O(N2437) );
buf1 gate604( .a(N2144), .O(N2440) );
buf1 gate605( .a(N2141), .O(N2443) );
buf1 gate606( .a(N2150), .O(N2446) );
buf1 gate607( .a(N2147), .O(N2449) );
inv1 gate608( .a(N2197), .O(N2452) );

  xor2  gate2530(.a(N2200), .b(N2197), .O(gate609inter0));
  nand2 gate2531(.a(gate609inter0), .b(s_180), .O(gate609inter1));
  and2  gate2532(.a(N2200), .b(N2197), .O(gate609inter2));
  inv1  gate2533(.a(s_180), .O(gate609inter3));
  inv1  gate2534(.a(s_181), .O(gate609inter4));
  nand2 gate2535(.a(gate609inter4), .b(gate609inter3), .O(gate609inter5));
  nor2  gate2536(.a(gate609inter5), .b(gate609inter2), .O(gate609inter6));
  inv1  gate2537(.a(N2197), .O(gate609inter7));
  inv1  gate2538(.a(N2200), .O(gate609inter8));
  nand2 gate2539(.a(gate609inter8), .b(gate609inter7), .O(gate609inter9));
  nand2 gate2540(.a(s_181), .b(gate609inter3), .O(gate609inter10));
  nor2  gate2541(.a(gate609inter10), .b(gate609inter9), .O(gate609inter11));
  nor2  gate2542(.a(gate609inter11), .b(gate609inter6), .O(gate609inter12));
  nand2 gate2543(.a(gate609inter12), .b(gate609inter1), .O(N2453));
buf1 gate610( .a(N2128), .O(N2454) );
buf1 gate611( .a(N2144), .O(N2457) );
buf1 gate612( .a(N2141), .O(N2460) );
buf1 gate613( .a(N2150), .O(N2463) );
buf1 gate614( .a(N2147), .O(N2466) );
inv1 gate615( .a(N2120), .O(N2469) );
buf1 gate616( .a(N2128), .O(N2472) );
buf1 gate617( .a(N2135), .O(N2475) );
buf1 gate618( .a(N2128), .O(N2478) );
buf1 gate619( .a(N2135), .O(N2481) );

  xor2  gate2712(.a(N2297), .b(N2298), .O(gate620inter0));
  nand2 gate2713(.a(gate620inter0), .b(s_206), .O(gate620inter1));
  and2  gate2714(.a(N2297), .b(N2298), .O(gate620inter2));
  inv1  gate2715(.a(s_206), .O(gate620inter3));
  inv1  gate2716(.a(s_207), .O(gate620inter4));
  nand2 gate2717(.a(gate620inter4), .b(gate620inter3), .O(gate620inter5));
  nor2  gate2718(.a(gate620inter5), .b(gate620inter2), .O(gate620inter6));
  inv1  gate2719(.a(N2298), .O(gate620inter7));
  inv1  gate2720(.a(N2297), .O(gate620inter8));
  nand2 gate2721(.a(gate620inter8), .b(gate620inter7), .O(gate620inter9));
  nand2 gate2722(.a(s_207), .b(gate620inter3), .O(gate620inter10));
  nor2  gate2723(.a(gate620inter10), .b(gate620inter9), .O(gate620inter11));
  nor2  gate2724(.a(gate620inter11), .b(gate620inter6), .O(gate620inter12));
  nand2 gate2725(.a(gate620inter12), .b(gate620inter1), .O(N2484));
nand2 gate621( .a(N2356), .b(N2357), .O(N2487) );
nand2 gate622( .a(N2354), .b(N2355), .O(N2490) );
nand2 gate623( .a(N2328), .b(N2327), .O(N2493) );
or2 gate624( .a(N2358), .b(N1814), .O(N2496) );

  xor2  gate1844(.a(N2364), .b(N2188), .O(gate625inter0));
  nand2 gate1845(.a(gate625inter0), .b(s_82), .O(gate625inter1));
  and2  gate1846(.a(N2364), .b(N2188), .O(gate625inter2));
  inv1  gate1847(.a(s_82), .O(gate625inter3));
  inv1  gate1848(.a(s_83), .O(gate625inter4));
  nand2 gate1849(.a(gate625inter4), .b(gate625inter3), .O(gate625inter5));
  nor2  gate1850(.a(gate625inter5), .b(gate625inter2), .O(gate625inter6));
  inv1  gate1851(.a(N2188), .O(gate625inter7));
  inv1  gate1852(.a(N2364), .O(gate625inter8));
  nand2 gate1853(.a(gate625inter8), .b(gate625inter7), .O(gate625inter9));
  nand2 gate1854(.a(s_83), .b(gate625inter3), .O(gate625inter10));
  nor2  gate1855(.a(gate625inter10), .b(gate625inter9), .O(gate625inter11));
  nor2  gate1856(.a(gate625inter11), .b(gate625inter6), .O(gate625inter12));
  nand2 gate1857(.a(gate625inter12), .b(gate625inter1), .O(N2503));

  xor2  gate1340(.a(N2365), .b(N2185), .O(gate626inter0));
  nand2 gate1341(.a(gate626inter0), .b(s_10), .O(gate626inter1));
  and2  gate1342(.a(N2365), .b(N2185), .O(gate626inter2));
  inv1  gate1343(.a(s_10), .O(gate626inter3));
  inv1  gate1344(.a(s_11), .O(gate626inter4));
  nand2 gate1345(.a(gate626inter4), .b(gate626inter3), .O(gate626inter5));
  nor2  gate1346(.a(gate626inter5), .b(gate626inter2), .O(gate626inter6));
  inv1  gate1347(.a(N2185), .O(gate626inter7));
  inv1  gate1348(.a(N2365), .O(gate626inter8));
  nand2 gate1349(.a(gate626inter8), .b(gate626inter7), .O(gate626inter9));
  nand2 gate1350(.a(s_11), .b(gate626inter3), .O(gate626inter10));
  nor2  gate1351(.a(gate626inter10), .b(gate626inter9), .O(gate626inter11));
  nor2  gate1352(.a(gate626inter11), .b(gate626inter6), .O(gate626inter12));
  nand2 gate1353(.a(gate626inter12), .b(gate626inter1), .O(N2504));

  xor2  gate2488(.a(N2372), .b(N2204), .O(gate627inter0));
  nand2 gate2489(.a(gate627inter0), .b(s_174), .O(gate627inter1));
  and2  gate2490(.a(N2372), .b(N2204), .O(gate627inter2));
  inv1  gate2491(.a(s_174), .O(gate627inter3));
  inv1  gate2492(.a(s_175), .O(gate627inter4));
  nand2 gate2493(.a(gate627inter4), .b(gate627inter3), .O(gate627inter5));
  nor2  gate2494(.a(gate627inter5), .b(gate627inter2), .O(gate627inter6));
  inv1  gate2495(.a(N2204), .O(gate627inter7));
  inv1  gate2496(.a(N2372), .O(gate627inter8));
  nand2 gate2497(.a(gate627inter8), .b(gate627inter7), .O(gate627inter9));
  nand2 gate2498(.a(s_175), .b(gate627inter3), .O(gate627inter10));
  nor2  gate2499(.a(gate627inter10), .b(gate627inter9), .O(gate627inter11));
  nor2  gate2500(.a(gate627inter11), .b(gate627inter6), .O(gate627inter12));
  nand2 gate2501(.a(gate627inter12), .b(gate627inter1), .O(N2510));
nand2 gate628( .a(N2201), .b(N2373), .O(N2511) );
or2 gate629( .a(N1830), .b(N2386), .O(N2521) );

  xor2  gate2754(.a(N2406), .b(N2046), .O(gate630inter0));
  nand2 gate2755(.a(gate630inter0), .b(s_212), .O(gate630inter1));
  and2  gate2756(.a(N2406), .b(N2046), .O(gate630inter2));
  inv1  gate2757(.a(s_212), .O(gate630inter3));
  inv1  gate2758(.a(s_213), .O(gate630inter4));
  nand2 gate2759(.a(gate630inter4), .b(gate630inter3), .O(gate630inter5));
  nor2  gate2760(.a(gate630inter5), .b(gate630inter2), .O(gate630inter6));
  inv1  gate2761(.a(N2046), .O(gate630inter7));
  inv1  gate2762(.a(N2406), .O(gate630inter8));
  nand2 gate2763(.a(gate630inter8), .b(gate630inter7), .O(gate630inter9));
  nand2 gate2764(.a(s_213), .b(gate630inter3), .O(gate630inter10));
  nor2  gate2765(.a(gate630inter10), .b(gate630inter9), .O(gate630inter11));
  nor2  gate2766(.a(gate630inter11), .b(gate630inter6), .O(gate630inter12));
  nand2 gate2767(.a(gate630inter12), .b(gate630inter1), .O(N2528));
inv1 gate631( .a(N2291), .O(N2531) );
inv1 gate632( .a(N2294), .O(N2534) );
buf1 gate633( .a(N2250), .O(N2537) );
buf1 gate634( .a(N2250), .O(N2540) );

  xor2  gate1718(.a(N2407), .b(N2302), .O(gate635inter0));
  nand2 gate1719(.a(gate635inter0), .b(s_64), .O(gate635inter1));
  and2  gate1720(.a(N2407), .b(N2302), .O(gate635inter2));
  inv1  gate1721(.a(s_64), .O(gate635inter3));
  inv1  gate1722(.a(s_65), .O(gate635inter4));
  nand2 gate1723(.a(gate635inter4), .b(gate635inter3), .O(gate635inter5));
  nor2  gate1724(.a(gate635inter5), .b(gate635inter2), .O(gate635inter6));
  inv1  gate1725(.a(N2302), .O(gate635inter7));
  inv1  gate1726(.a(N2407), .O(gate635inter8));
  nand2 gate1727(.a(gate635inter8), .b(gate635inter7), .O(gate635inter9));
  nand2 gate1728(.a(s_65), .b(gate635inter3), .O(gate635inter10));
  nor2  gate1729(.a(gate635inter10), .b(gate635inter9), .O(gate635inter11));
  nor2  gate1730(.a(gate635inter11), .b(gate635inter6), .O(gate635inter12));
  nand2 gate1731(.a(gate635inter12), .b(gate635inter1), .O(N2544));
nand2 gate636( .a(N2304), .b(N2408), .O(N2545) );
nand2 gate637( .a(N2306), .b(N2409), .O(N2546) );

  xor2  gate2334(.a(N2410), .b(N2308), .O(gate638inter0));
  nand2 gate2335(.a(gate638inter0), .b(s_152), .O(gate638inter1));
  and2  gate2336(.a(N2410), .b(N2308), .O(gate638inter2));
  inv1  gate2337(.a(s_152), .O(gate638inter3));
  inv1  gate2338(.a(s_153), .O(gate638inter4));
  nand2 gate2339(.a(gate638inter4), .b(gate638inter3), .O(gate638inter5));
  nor2  gate2340(.a(gate638inter5), .b(gate638inter2), .O(gate638inter6));
  inv1  gate2341(.a(N2308), .O(gate638inter7));
  inv1  gate2342(.a(N2410), .O(gate638inter8));
  nand2 gate2343(.a(gate638inter8), .b(gate638inter7), .O(gate638inter9));
  nand2 gate2344(.a(s_153), .b(gate638inter3), .O(gate638inter10));
  nor2  gate2345(.a(gate638inter10), .b(gate638inter9), .O(gate638inter11));
  nor2  gate2346(.a(gate638inter11), .b(gate638inter6), .O(gate638inter12));
  nand2 gate2347(.a(gate638inter12), .b(gate638inter1), .O(N2547));
nand2 gate639( .a(N2310), .b(N2411), .O(N2548) );
nand2 gate640( .a(N2312), .b(N2412), .O(N2549) );

  xor2  gate1984(.a(N2413), .b(N2314), .O(gate641inter0));
  nand2 gate1985(.a(gate641inter0), .b(s_102), .O(gate641inter1));
  and2  gate1986(.a(N2413), .b(N2314), .O(gate641inter2));
  inv1  gate1987(.a(s_102), .O(gate641inter3));
  inv1  gate1988(.a(s_103), .O(gate641inter4));
  nand2 gate1989(.a(gate641inter4), .b(gate641inter3), .O(gate641inter5));
  nor2  gate1990(.a(gate641inter5), .b(gate641inter2), .O(gate641inter6));
  inv1  gate1991(.a(N2314), .O(gate641inter7));
  inv1  gate1992(.a(N2413), .O(gate641inter8));
  nand2 gate1993(.a(gate641inter8), .b(gate641inter7), .O(gate641inter9));
  nand2 gate1994(.a(s_103), .b(gate641inter3), .O(gate641inter10));
  nor2  gate1995(.a(gate641inter10), .b(gate641inter9), .O(gate641inter11));
  nor2  gate1996(.a(gate641inter11), .b(gate641inter6), .O(gate641inter12));
  nand2 gate1997(.a(gate641inter12), .b(gate641inter1), .O(N2550));
nand2 gate642( .a(N2316), .b(N2414), .O(N2551) );
nand2 gate643( .a(N2318), .b(N2415), .O(N2552) );
nand2 gate644( .a(N2320), .b(N2416), .O(N2553) );

  xor2  gate1928(.a(N2428), .b(N2329), .O(gate645inter0));
  nand2 gate1929(.a(gate645inter0), .b(s_94), .O(gate645inter1));
  and2  gate1930(.a(N2428), .b(N2329), .O(gate645inter2));
  inv1  gate1931(.a(s_94), .O(gate645inter3));
  inv1  gate1932(.a(s_95), .O(gate645inter4));
  nand2 gate1933(.a(gate645inter4), .b(gate645inter3), .O(gate645inter5));
  nor2  gate1934(.a(gate645inter5), .b(gate645inter2), .O(gate645inter6));
  inv1  gate1935(.a(N2329), .O(gate645inter7));
  inv1  gate1936(.a(N2428), .O(gate645inter8));
  nand2 gate1937(.a(gate645inter8), .b(gate645inter7), .O(gate645inter9));
  nand2 gate1938(.a(s_95), .b(gate645inter3), .O(gate645inter10));
  nor2  gate1939(.a(gate645inter10), .b(gate645inter9), .O(gate645inter11));
  nor2  gate1940(.a(gate645inter11), .b(gate645inter6), .O(gate645inter12));
  nand2 gate1941(.a(gate645inter12), .b(gate645inter1), .O(N2563));
nand2 gate646( .a(N2331), .b(N2429), .O(N2564) );
nand2 gate647( .a(N2333), .b(N2430), .O(N2565) );
nand2 gate648( .a(N2335), .b(N2431), .O(N2566) );
nand2 gate649( .a(N2337), .b(N2432), .O(N2567) );
nand2 gate650( .a(N2339), .b(N2433), .O(N2568) );

  xor2  gate2096(.a(N2452), .b(N1936), .O(gate651inter0));
  nand2 gate2097(.a(gate651inter0), .b(s_118), .O(gate651inter1));
  and2  gate2098(.a(N2452), .b(N1936), .O(gate651inter2));
  inv1  gate2099(.a(s_118), .O(gate651inter3));
  inv1  gate2100(.a(s_119), .O(gate651inter4));
  nand2 gate2101(.a(gate651inter4), .b(gate651inter3), .O(gate651inter5));
  nor2  gate2102(.a(gate651inter5), .b(gate651inter2), .O(gate651inter6));
  inv1  gate2103(.a(N1936), .O(gate651inter7));
  inv1  gate2104(.a(N2452), .O(gate651inter8));
  nand2 gate2105(.a(gate651inter8), .b(gate651inter7), .O(gate651inter9));
  nand2 gate2106(.a(s_119), .b(gate651inter3), .O(gate651inter10));
  nor2  gate2107(.a(gate651inter10), .b(gate651inter9), .O(gate651inter11));
  nor2  gate2108(.a(gate651inter11), .b(gate651inter6), .O(gate651inter12));
  nand2 gate2109(.a(gate651inter12), .b(gate651inter1), .O(N2579));
buf1 gate652( .a(N2359), .O(N2603) );
and2 gate653( .a(N1880), .b(N2377), .O(N2607) );
and2 gate654( .a(N1676), .b(N2377), .O(N2608) );
and2 gate655( .a(N1681), .b(N2377), .O(N2609) );
and2 gate656( .a(N1891), .b(N2377), .O(N2610) );
and2 gate657( .a(N1856), .b(N2382), .O(N2611) );
and2 gate658( .a(N1863), .b(N2382), .O(N2612) );
nand2 gate659( .a(N2503), .b(N2504), .O(N2613) );
inv1 gate660( .a(N2434), .O(N2617) );

  xor2  gate1508(.a(N2366), .b(N2434), .O(gate661inter0));
  nand2 gate1509(.a(gate661inter0), .b(s_34), .O(gate661inter1));
  and2  gate1510(.a(N2366), .b(N2434), .O(gate661inter2));
  inv1  gate1511(.a(s_34), .O(gate661inter3));
  inv1  gate1512(.a(s_35), .O(gate661inter4));
  nand2 gate1513(.a(gate661inter4), .b(gate661inter3), .O(gate661inter5));
  nor2  gate1514(.a(gate661inter5), .b(gate661inter2), .O(gate661inter6));
  inv1  gate1515(.a(N2434), .O(gate661inter7));
  inv1  gate1516(.a(N2366), .O(gate661inter8));
  nand2 gate1517(.a(gate661inter8), .b(gate661inter7), .O(gate661inter9));
  nand2 gate1518(.a(s_35), .b(gate661inter3), .O(gate661inter10));
  nor2  gate1519(.a(gate661inter10), .b(gate661inter9), .O(gate661inter11));
  nor2  gate1520(.a(gate661inter11), .b(gate661inter6), .O(gate661inter12));
  nand2 gate1521(.a(gate661inter12), .b(gate661inter1), .O(N2618));

  xor2  gate2922(.a(N2367), .b(N2437), .O(gate662inter0));
  nand2 gate2923(.a(gate662inter0), .b(s_236), .O(gate662inter1));
  and2  gate2924(.a(N2367), .b(N2437), .O(gate662inter2));
  inv1  gate2925(.a(s_236), .O(gate662inter3));
  inv1  gate2926(.a(s_237), .O(gate662inter4));
  nand2 gate2927(.a(gate662inter4), .b(gate662inter3), .O(gate662inter5));
  nor2  gate2928(.a(gate662inter5), .b(gate662inter2), .O(gate662inter6));
  inv1  gate2929(.a(N2437), .O(gate662inter7));
  inv1  gate2930(.a(N2367), .O(gate662inter8));
  nand2 gate2931(.a(gate662inter8), .b(gate662inter7), .O(gate662inter9));
  nand2 gate2932(.a(s_237), .b(gate662inter3), .O(gate662inter10));
  nor2  gate2933(.a(gate662inter10), .b(gate662inter9), .O(gate662inter11));
  nor2  gate2934(.a(gate662inter11), .b(gate662inter6), .O(gate662inter12));
  nand2 gate2935(.a(gate662inter12), .b(gate662inter1), .O(N2619));
inv1 gate663( .a(N2437), .O(N2620) );
inv1 gate664( .a(N2368), .O(N2621) );
nand2 gate665( .a(N2510), .b(N2511), .O(N2624) );
inv1 gate666( .a(N2454), .O(N2628) );
nand2 gate667( .a(N2454), .b(N2374), .O(N2629) );
inv1 gate668( .a(N2472), .O(N2630) );
and2 gate669( .a(N1856), .b(N2391), .O(N2631) );
and2 gate670( .a(N1863), .b(N2391), .O(N2632) );
and2 gate671( .a(N1880), .b(N2395), .O(N2633) );
and2 gate672( .a(N1676), .b(N2395), .O(N2634) );
and2 gate673( .a(N1681), .b(N2395), .O(N2635) );
and2 gate674( .a(N1891), .b(N2395), .O(N2636) );
inv1 gate675( .a(N2382), .O(N2638) );
buf1 gate676( .a(N2521), .O(N2643) );
buf1 gate677( .a(N2521), .O(N2644) );
inv1 gate678( .a(N2475), .O(N2645) );
inv1 gate679( .a(N2391), .O(N2646) );

  xor2  gate2012(.a(N2400), .b(N2528), .O(gate680inter0));
  nand2 gate2013(.a(gate680inter0), .b(s_106), .O(gate680inter1));
  and2  gate2014(.a(N2400), .b(N2528), .O(gate680inter2));
  inv1  gate2015(.a(s_106), .O(gate680inter3));
  inv1  gate2016(.a(s_107), .O(gate680inter4));
  nand2 gate2017(.a(gate680inter4), .b(gate680inter3), .O(gate680inter5));
  nor2  gate2018(.a(gate680inter5), .b(gate680inter2), .O(gate680inter6));
  inv1  gate2019(.a(N2528), .O(gate680inter7));
  inv1  gate2020(.a(N2400), .O(gate680inter8));
  nand2 gate2021(.a(gate680inter8), .b(gate680inter7), .O(gate680inter9));
  nand2 gate2022(.a(s_107), .b(gate680inter3), .O(gate680inter10));
  nor2  gate2023(.a(gate680inter10), .b(gate680inter9), .O(gate680inter11));
  nor2  gate2024(.a(gate680inter11), .b(gate680inter6), .O(gate680inter12));
  nand2 gate2025(.a(gate680inter12), .b(gate680inter1), .O(N2652));
inv1 gate681( .a(N2478), .O(N2655) );
inv1 gate682( .a(N2481), .O(N2656) );
buf1 gate683( .a(N2359), .O(N2659) );
inv1 gate684( .a(N2484), .O(N2663) );

  xor2  gate2250(.a(N2301), .b(N2484), .O(gate685inter0));
  nand2 gate2251(.a(gate685inter0), .b(s_140), .O(gate685inter1));
  and2  gate2252(.a(N2301), .b(N2484), .O(gate685inter2));
  inv1  gate2253(.a(s_140), .O(gate685inter3));
  inv1  gate2254(.a(s_141), .O(gate685inter4));
  nand2 gate2255(.a(gate685inter4), .b(gate685inter3), .O(gate685inter5));
  nor2  gate2256(.a(gate685inter5), .b(gate685inter2), .O(gate685inter6));
  inv1  gate2257(.a(N2484), .O(gate685inter7));
  inv1  gate2258(.a(N2301), .O(gate685inter8));
  nand2 gate2259(.a(gate685inter8), .b(gate685inter7), .O(gate685inter9));
  nand2 gate2260(.a(s_141), .b(gate685inter3), .O(gate685inter10));
  nor2  gate2261(.a(gate685inter10), .b(gate685inter9), .O(gate685inter11));
  nor2  gate2262(.a(gate685inter11), .b(gate685inter6), .O(gate685inter12));
  nand2 gate2263(.a(gate685inter12), .b(gate685inter1), .O(N2664));
inv1 gate686( .a(N2553), .O(N2665) );
inv1 gate687( .a(N2552), .O(N2666) );
inv1 gate688( .a(N2551), .O(N2667) );
inv1 gate689( .a(N2550), .O(N2668) );
inv1 gate690( .a(N2549), .O(N2669) );
inv1 gate691( .a(N2548), .O(N2670) );
inv1 gate692( .a(N2547), .O(N2671) );
inv1 gate693( .a(N2546), .O(N2672) );
inv1 gate694( .a(N2545), .O(N2673) );
inv1 gate695( .a(N2544), .O(N2674) );
inv1 gate696( .a(N2568), .O(N2675) );
inv1 gate697( .a(N2567), .O(N2676) );
inv1 gate698( .a(N2566), .O(N2677) );
inv1 gate699( .a(N2565), .O(N2678) );
inv1 gate700( .a(N2564), .O(N2679) );
inv1 gate701( .a(N2563), .O(N2680) );
inv1 gate702( .a(N2417), .O(N2681) );
inv1 gate703( .a(N2421), .O(N2684) );
buf1 gate704( .a(N2425), .O(N2687) );
buf1 gate705( .a(N2425), .O(N2690) );
inv1 gate706( .a(N2493), .O(N2693) );
nand2 gate707( .a(N2493), .b(N1807), .O(N2694) );
inv1 gate708( .a(N2440), .O(N2695) );
inv1 gate709( .a(N2443), .O(N2696) );
inv1 gate710( .a(N2446), .O(N2697) );
inv1 gate711( .a(N2449), .O(N2698) );
inv1 gate712( .a(N2457), .O(N2699) );
inv1 gate713( .a(N2460), .O(N2700) );
inv1 gate714( .a(N2463), .O(N2701) );
inv1 gate715( .a(N2466), .O(N2702) );

  xor2  gate2614(.a(N2453), .b(N2579), .O(gate716inter0));
  nand2 gate2615(.a(gate716inter0), .b(s_192), .O(gate716inter1));
  and2  gate2616(.a(N2453), .b(N2579), .O(gate716inter2));
  inv1  gate2617(.a(s_192), .O(gate716inter3));
  inv1  gate2618(.a(s_193), .O(gate716inter4));
  nand2 gate2619(.a(gate716inter4), .b(gate716inter3), .O(gate716inter5));
  nor2  gate2620(.a(gate716inter5), .b(gate716inter2), .O(gate716inter6));
  inv1  gate2621(.a(N2579), .O(gate716inter7));
  inv1  gate2622(.a(N2453), .O(gate716inter8));
  nand2 gate2623(.a(gate716inter8), .b(gate716inter7), .O(gate716inter9));
  nand2 gate2624(.a(s_193), .b(gate716inter3), .O(gate716inter10));
  nor2  gate2625(.a(gate716inter10), .b(gate716inter9), .O(gate716inter11));
  nor2  gate2626(.a(gate716inter11), .b(gate716inter6), .O(gate716inter12));
  nand2 gate2627(.a(gate716inter12), .b(gate716inter1), .O(N2703));
inv1 gate717( .a(N2469), .O(N2706) );
inv1 gate718( .a(N2487), .O(N2707) );
inv1 gate719( .a(N2490), .O(N2708) );
and2 gate720( .a(N2294), .b(N2534), .O(N2709) );
and2 gate721( .a(N2291), .b(N2531), .O(N2710) );

  xor2  gate2894(.a(N2617), .b(N2191), .O(gate722inter0));
  nand2 gate2895(.a(gate722inter0), .b(s_232), .O(gate722inter1));
  and2  gate2896(.a(N2617), .b(N2191), .O(gate722inter2));
  inv1  gate2897(.a(s_232), .O(gate722inter3));
  inv1  gate2898(.a(s_233), .O(gate722inter4));
  nand2 gate2899(.a(gate722inter4), .b(gate722inter3), .O(gate722inter5));
  nor2  gate2900(.a(gate722inter5), .b(gate722inter2), .O(gate722inter6));
  inv1  gate2901(.a(N2191), .O(gate722inter7));
  inv1  gate2902(.a(N2617), .O(gate722inter8));
  nand2 gate2903(.a(gate722inter8), .b(gate722inter7), .O(gate722inter9));
  nand2 gate2904(.a(s_233), .b(gate722inter3), .O(gate722inter10));
  nor2  gate2905(.a(gate722inter10), .b(gate722inter9), .O(gate722inter11));
  nor2  gate2906(.a(gate722inter11), .b(gate722inter6), .O(gate722inter12));
  nand2 gate2907(.a(gate722inter12), .b(gate722inter1), .O(N2719));
nand2 gate723( .a(N2194), .b(N2620), .O(N2720) );

  xor2  gate2474(.a(N2628), .b(N2207), .O(gate724inter0));
  nand2 gate2475(.a(gate724inter0), .b(s_172), .O(gate724inter1));
  and2  gate2476(.a(N2628), .b(N2207), .O(gate724inter2));
  inv1  gate2477(.a(s_172), .O(gate724inter3));
  inv1  gate2478(.a(s_173), .O(gate724inter4));
  nand2 gate2479(.a(gate724inter4), .b(gate724inter3), .O(gate724inter5));
  nor2  gate2480(.a(gate724inter5), .b(gate724inter2), .O(gate724inter6));
  inv1  gate2481(.a(N2207), .O(gate724inter7));
  inv1  gate2482(.a(N2628), .O(gate724inter8));
  nand2 gate2483(.a(gate724inter8), .b(gate724inter7), .O(gate724inter9));
  nand2 gate2484(.a(s_173), .b(gate724inter3), .O(gate724inter10));
  nor2  gate2485(.a(gate724inter10), .b(gate724inter9), .O(gate724inter11));
  nor2  gate2486(.a(gate724inter11), .b(gate724inter6), .O(gate724inter12));
  nand2 gate2487(.a(gate724inter12), .b(gate724inter1), .O(N2726));
buf1 gate725( .a(N2537), .O(N2729) );
buf1 gate726( .a(N2537), .O(N2738) );
inv1 gate727( .a(N2652), .O(N2743) );
nand2 gate728( .a(N2049), .b(N2663), .O(N2747) );
and5 gate729( .a(N2665), .b(N2666), .c(N2667), .d(N2668), .e(N2669), .O(N2748) );
and5 gate730( .a(N2670), .b(N2671), .c(N2672), .d(N2673), .e(N2674), .O(N2749) );
and2 gate731( .a(N2034), .b(N2675), .O(N2750) );
and5 gate732( .a(N2676), .b(N2677), .c(N2678), .d(N2679), .e(N2680), .O(N2751) );

  xor2  gate1830(.a(N2693), .b(N1588), .O(gate733inter0));
  nand2 gate1831(.a(gate733inter0), .b(s_80), .O(gate733inter1));
  and2  gate1832(.a(N2693), .b(N1588), .O(gate733inter2));
  inv1  gate1833(.a(s_80), .O(gate733inter3));
  inv1  gate1834(.a(s_81), .O(gate733inter4));
  nand2 gate1835(.a(gate733inter4), .b(gate733inter3), .O(gate733inter5));
  nor2  gate1836(.a(gate733inter5), .b(gate733inter2), .O(gate733inter6));
  inv1  gate1837(.a(N1588), .O(gate733inter7));
  inv1  gate1838(.a(N2693), .O(gate733inter8));
  nand2 gate1839(.a(gate733inter8), .b(gate733inter7), .O(gate733inter9));
  nand2 gate1840(.a(s_81), .b(gate733inter3), .O(gate733inter10));
  nor2  gate1841(.a(gate733inter10), .b(gate733inter9), .O(gate733inter11));
  nor2  gate1842(.a(gate733inter11), .b(gate733inter6), .O(gate733inter12));
  nand2 gate1843(.a(gate733inter12), .b(gate733inter1), .O(N2760));
buf1 gate734( .a(N2540), .O(N2761) );
buf1 gate735( .a(N2540), .O(N2766) );

  xor2  gate2362(.a(N2695), .b(N2443), .O(gate736inter0));
  nand2 gate2363(.a(gate736inter0), .b(s_156), .O(gate736inter1));
  and2  gate2364(.a(N2695), .b(N2443), .O(gate736inter2));
  inv1  gate2365(.a(s_156), .O(gate736inter3));
  inv1  gate2366(.a(s_157), .O(gate736inter4));
  nand2 gate2367(.a(gate736inter4), .b(gate736inter3), .O(gate736inter5));
  nor2  gate2368(.a(gate736inter5), .b(gate736inter2), .O(gate736inter6));
  inv1  gate2369(.a(N2443), .O(gate736inter7));
  inv1  gate2370(.a(N2695), .O(gate736inter8));
  nand2 gate2371(.a(gate736inter8), .b(gate736inter7), .O(gate736inter9));
  nand2 gate2372(.a(s_157), .b(gate736inter3), .O(gate736inter10));
  nor2  gate2373(.a(gate736inter10), .b(gate736inter9), .O(gate736inter11));
  nor2  gate2374(.a(gate736inter11), .b(gate736inter6), .O(gate736inter12));
  nand2 gate2375(.a(gate736inter12), .b(gate736inter1), .O(N2771));

  xor2  gate1900(.a(N2696), .b(N2440), .O(gate737inter0));
  nand2 gate1901(.a(gate737inter0), .b(s_90), .O(gate737inter1));
  and2  gate1902(.a(N2696), .b(N2440), .O(gate737inter2));
  inv1  gate1903(.a(s_90), .O(gate737inter3));
  inv1  gate1904(.a(s_91), .O(gate737inter4));
  nand2 gate1905(.a(gate737inter4), .b(gate737inter3), .O(gate737inter5));
  nor2  gate1906(.a(gate737inter5), .b(gate737inter2), .O(gate737inter6));
  inv1  gate1907(.a(N2440), .O(gate737inter7));
  inv1  gate1908(.a(N2696), .O(gate737inter8));
  nand2 gate1909(.a(gate737inter8), .b(gate737inter7), .O(gate737inter9));
  nand2 gate1910(.a(s_91), .b(gate737inter3), .O(gate737inter10));
  nor2  gate1911(.a(gate737inter10), .b(gate737inter9), .O(gate737inter11));
  nor2  gate1912(.a(gate737inter11), .b(gate737inter6), .O(gate737inter12));
  nand2 gate1913(.a(gate737inter12), .b(gate737inter1), .O(N2772));

  xor2  gate1858(.a(N2697), .b(N2449), .O(gate738inter0));
  nand2 gate1859(.a(gate738inter0), .b(s_84), .O(gate738inter1));
  and2  gate1860(.a(N2697), .b(N2449), .O(gate738inter2));
  inv1  gate1861(.a(s_84), .O(gate738inter3));
  inv1  gate1862(.a(s_85), .O(gate738inter4));
  nand2 gate1863(.a(gate738inter4), .b(gate738inter3), .O(gate738inter5));
  nor2  gate1864(.a(gate738inter5), .b(gate738inter2), .O(gate738inter6));
  inv1  gate1865(.a(N2449), .O(gate738inter7));
  inv1  gate1866(.a(N2697), .O(gate738inter8));
  nand2 gate1867(.a(gate738inter8), .b(gate738inter7), .O(gate738inter9));
  nand2 gate1868(.a(s_85), .b(gate738inter3), .O(gate738inter10));
  nor2  gate1869(.a(gate738inter10), .b(gate738inter9), .O(gate738inter11));
  nor2  gate1870(.a(gate738inter11), .b(gate738inter6), .O(gate738inter12));
  nand2 gate1871(.a(gate738inter12), .b(gate738inter1), .O(N2773));

  xor2  gate1998(.a(N2698), .b(N2446), .O(gate739inter0));
  nand2 gate1999(.a(gate739inter0), .b(s_104), .O(gate739inter1));
  and2  gate2000(.a(N2698), .b(N2446), .O(gate739inter2));
  inv1  gate2001(.a(s_104), .O(gate739inter3));
  inv1  gate2002(.a(s_105), .O(gate739inter4));
  nand2 gate2003(.a(gate739inter4), .b(gate739inter3), .O(gate739inter5));
  nor2  gate2004(.a(gate739inter5), .b(gate739inter2), .O(gate739inter6));
  inv1  gate2005(.a(N2446), .O(gate739inter7));
  inv1  gate2006(.a(N2698), .O(gate739inter8));
  nand2 gate2007(.a(gate739inter8), .b(gate739inter7), .O(gate739inter9));
  nand2 gate2008(.a(s_105), .b(gate739inter3), .O(gate739inter10));
  nor2  gate2009(.a(gate739inter10), .b(gate739inter9), .O(gate739inter11));
  nor2  gate2010(.a(gate739inter11), .b(gate739inter6), .O(gate739inter12));
  nand2 gate2011(.a(gate739inter12), .b(gate739inter1), .O(N2774));
nand2 gate740( .a(N2460), .b(N2699), .O(N2775) );
nand2 gate741( .a(N2457), .b(N2700), .O(N2776) );
nand2 gate742( .a(N2466), .b(N2701), .O(N2777) );

  xor2  gate1298(.a(N2702), .b(N2463), .O(gate743inter0));
  nand2 gate1299(.a(gate743inter0), .b(s_4), .O(gate743inter1));
  and2  gate1300(.a(N2702), .b(N2463), .O(gate743inter2));
  inv1  gate1301(.a(s_4), .O(gate743inter3));
  inv1  gate1302(.a(s_5), .O(gate743inter4));
  nand2 gate1303(.a(gate743inter4), .b(gate743inter3), .O(gate743inter5));
  nor2  gate1304(.a(gate743inter5), .b(gate743inter2), .O(gate743inter6));
  inv1  gate1305(.a(N2463), .O(gate743inter7));
  inv1  gate1306(.a(N2702), .O(gate743inter8));
  nand2 gate1307(.a(gate743inter8), .b(gate743inter7), .O(gate743inter9));
  nand2 gate1308(.a(s_5), .b(gate743inter3), .O(gate743inter10));
  nor2  gate1309(.a(gate743inter10), .b(gate743inter9), .O(gate743inter11));
  nor2  gate1310(.a(gate743inter11), .b(gate743inter6), .O(gate743inter12));
  nand2 gate1311(.a(gate743inter12), .b(gate743inter1), .O(N2778));
nand2 gate744( .a(N2490), .b(N2707), .O(N2781) );
nand2 gate745( .a(N2487), .b(N2708), .O(N2782) );
or2 gate746( .a(N2709), .b(N2534), .O(N2783) );
or2 gate747( .a(N2710), .b(N2531), .O(N2784) );
and2 gate748( .a(N1856), .b(N2638), .O(N2789) );
and2 gate749( .a(N1863), .b(N2638), .O(N2790) );
and2 gate750( .a(N1870), .b(N2638), .O(N2791) );
and2 gate751( .a(N1875), .b(N2638), .O(N2792) );
inv1 gate752( .a(N2613), .O(N2793) );

  xor2  gate2502(.a(N2618), .b(N2719), .O(gate753inter0));
  nand2 gate2503(.a(gate753inter0), .b(s_176), .O(gate753inter1));
  and2  gate2504(.a(N2618), .b(N2719), .O(gate753inter2));
  inv1  gate2505(.a(s_176), .O(gate753inter3));
  inv1  gate2506(.a(s_177), .O(gate753inter4));
  nand2 gate2507(.a(gate753inter4), .b(gate753inter3), .O(gate753inter5));
  nor2  gate2508(.a(gate753inter5), .b(gate753inter2), .O(gate753inter6));
  inv1  gate2509(.a(N2719), .O(gate753inter7));
  inv1  gate2510(.a(N2618), .O(gate753inter8));
  nand2 gate2511(.a(gate753inter8), .b(gate753inter7), .O(gate753inter9));
  nand2 gate2512(.a(s_177), .b(gate753inter3), .O(gate753inter10));
  nor2  gate2513(.a(gate753inter10), .b(gate753inter9), .O(gate753inter11));
  nor2  gate2514(.a(gate753inter11), .b(gate753inter6), .O(gate753inter12));
  nand2 gate2515(.a(gate753inter12), .b(gate753inter1), .O(N2796));

  xor2  gate2082(.a(N2720), .b(N2619), .O(gate754inter0));
  nand2 gate2083(.a(gate754inter0), .b(s_116), .O(gate754inter1));
  and2  gate2084(.a(N2720), .b(N2619), .O(gate754inter2));
  inv1  gate2085(.a(s_116), .O(gate754inter3));
  inv1  gate2086(.a(s_117), .O(gate754inter4));
  nand2 gate2087(.a(gate754inter4), .b(gate754inter3), .O(gate754inter5));
  nor2  gate2088(.a(gate754inter5), .b(gate754inter2), .O(gate754inter6));
  inv1  gate2089(.a(N2619), .O(gate754inter7));
  inv1  gate2090(.a(N2720), .O(gate754inter8));
  nand2 gate2091(.a(gate754inter8), .b(gate754inter7), .O(gate754inter9));
  nand2 gate2092(.a(s_117), .b(gate754inter3), .O(gate754inter10));
  nor2  gate2093(.a(gate754inter10), .b(gate754inter9), .O(gate754inter11));
  nor2  gate2094(.a(gate754inter11), .b(gate754inter6), .O(gate754inter12));
  nand2 gate2095(.a(gate754inter12), .b(gate754inter1), .O(N2800));
inv1 gate755( .a(N2624), .O(N2803) );

  xor2  gate2810(.a(N2629), .b(N2726), .O(gate756inter0));
  nand2 gate2811(.a(gate756inter0), .b(s_220), .O(gate756inter1));
  and2  gate2812(.a(N2629), .b(N2726), .O(gate756inter2));
  inv1  gate2813(.a(s_220), .O(gate756inter3));
  inv1  gate2814(.a(s_221), .O(gate756inter4));
  nand2 gate2815(.a(gate756inter4), .b(gate756inter3), .O(gate756inter5));
  nor2  gate2816(.a(gate756inter5), .b(gate756inter2), .O(gate756inter6));
  inv1  gate2817(.a(N2726), .O(gate756inter7));
  inv1  gate2818(.a(N2629), .O(gate756inter8));
  nand2 gate2819(.a(gate756inter8), .b(gate756inter7), .O(gate756inter9));
  nand2 gate2820(.a(s_221), .b(gate756inter3), .O(gate756inter10));
  nor2  gate2821(.a(gate756inter10), .b(gate756inter9), .O(gate756inter11));
  nor2  gate2822(.a(gate756inter11), .b(gate756inter6), .O(gate756inter12));
  nand2 gate2823(.a(gate756inter12), .b(gate756inter1), .O(N2806));
and2 gate757( .a(N1856), .b(N2646), .O(N2809) );
and2 gate758( .a(N1863), .b(N2646), .O(N2810) );
and2 gate759( .a(N1870), .b(N2646), .O(N2811) );
and2 gate760( .a(N1875), .b(N2646), .O(N2812) );
and2 gate761( .a(N2743), .b(N14), .O(N2817) );
buf1 gate762( .a(N2603), .O(N2820) );

  xor2  gate1592(.a(N2664), .b(N2747), .O(gate763inter0));
  nand2 gate1593(.a(gate763inter0), .b(s_46), .O(gate763inter1));
  and2  gate1594(.a(N2664), .b(N2747), .O(gate763inter2));
  inv1  gate1595(.a(s_46), .O(gate763inter3));
  inv1  gate1596(.a(s_47), .O(gate763inter4));
  nand2 gate1597(.a(gate763inter4), .b(gate763inter3), .O(gate763inter5));
  nor2  gate1598(.a(gate763inter5), .b(gate763inter2), .O(gate763inter6));
  inv1  gate1599(.a(N2747), .O(gate763inter7));
  inv1  gate1600(.a(N2664), .O(gate763inter8));
  nand2 gate1601(.a(gate763inter8), .b(gate763inter7), .O(gate763inter9));
  nand2 gate1602(.a(s_47), .b(gate763inter3), .O(gate763inter10));
  nor2  gate1603(.a(gate763inter10), .b(gate763inter9), .O(gate763inter11));
  nor2  gate1604(.a(gate763inter11), .b(gate763inter6), .O(gate763inter12));
  nand2 gate1605(.a(gate763inter12), .b(gate763inter1), .O(N2826));
and2 gate764( .a(N2748), .b(N2749), .O(N2829) );
and2 gate765( .a(N2750), .b(N2751), .O(N2830) );
buf1 gate766( .a(N2659), .O(N2831) );
inv1 gate767( .a(N2687), .O(N2837) );
inv1 gate768( .a(N2690), .O(N2838) );
and3 gate769( .a(N2421), .b(N2417), .c(N2687), .O(N2839) );
and3 gate770( .a(N2684), .b(N2681), .c(N2690), .O(N2840) );
nand2 gate771( .a(N2760), .b(N2694), .O(N2841) );
buf1 gate772( .a(N2603), .O(N2844) );
buf1 gate773( .a(N2603), .O(N2854) );
buf1 gate774( .a(N2659), .O(N2859) );
buf1 gate775( .a(N2659), .O(N2869) );

  xor2  gate2558(.a(N2774), .b(N2773), .O(gate776inter0));
  nand2 gate2559(.a(gate776inter0), .b(s_184), .O(gate776inter1));
  and2  gate2560(.a(N2774), .b(N2773), .O(gate776inter2));
  inv1  gate2561(.a(s_184), .O(gate776inter3));
  inv1  gate2562(.a(s_185), .O(gate776inter4));
  nand2 gate2563(.a(gate776inter4), .b(gate776inter3), .O(gate776inter5));
  nor2  gate2564(.a(gate776inter5), .b(gate776inter2), .O(gate776inter6));
  inv1  gate2565(.a(N2773), .O(gate776inter7));
  inv1  gate2566(.a(N2774), .O(gate776inter8));
  nand2 gate2567(.a(gate776inter8), .b(gate776inter7), .O(gate776inter9));
  nand2 gate2568(.a(s_185), .b(gate776inter3), .O(gate776inter10));
  nor2  gate2569(.a(gate776inter10), .b(gate776inter9), .O(gate776inter11));
  nor2  gate2570(.a(gate776inter11), .b(gate776inter6), .O(gate776inter12));
  nand2 gate2571(.a(gate776inter12), .b(gate776inter1), .O(N2874));

  xor2  gate2222(.a(N2772), .b(N2771), .O(gate777inter0));
  nand2 gate2223(.a(gate777inter0), .b(s_136), .O(gate777inter1));
  and2  gate2224(.a(N2772), .b(N2771), .O(gate777inter2));
  inv1  gate2225(.a(s_136), .O(gate777inter3));
  inv1  gate2226(.a(s_137), .O(gate777inter4));
  nand2 gate2227(.a(gate777inter4), .b(gate777inter3), .O(gate777inter5));
  nor2  gate2228(.a(gate777inter5), .b(gate777inter2), .O(gate777inter6));
  inv1  gate2229(.a(N2771), .O(gate777inter7));
  inv1  gate2230(.a(N2772), .O(gate777inter8));
  nand2 gate2231(.a(gate777inter8), .b(gate777inter7), .O(gate777inter9));
  nand2 gate2232(.a(s_137), .b(gate777inter3), .O(gate777inter10));
  nor2  gate2233(.a(gate777inter10), .b(gate777inter9), .O(gate777inter11));
  nor2  gate2234(.a(gate777inter11), .b(gate777inter6), .O(gate777inter12));
  nand2 gate2235(.a(gate777inter12), .b(gate777inter1), .O(N2877));
inv1 gate778( .a(N2703), .O(N2880) );

  xor2  gate2432(.a(N2706), .b(N2703), .O(gate779inter0));
  nand2 gate2433(.a(gate779inter0), .b(s_166), .O(gate779inter1));
  and2  gate2434(.a(N2706), .b(N2703), .O(gate779inter2));
  inv1  gate2435(.a(s_166), .O(gate779inter3));
  inv1  gate2436(.a(s_167), .O(gate779inter4));
  nand2 gate2437(.a(gate779inter4), .b(gate779inter3), .O(gate779inter5));
  nor2  gate2438(.a(gate779inter5), .b(gate779inter2), .O(gate779inter6));
  inv1  gate2439(.a(N2703), .O(gate779inter7));
  inv1  gate2440(.a(N2706), .O(gate779inter8));
  nand2 gate2441(.a(gate779inter8), .b(gate779inter7), .O(gate779inter9));
  nand2 gate2442(.a(s_167), .b(gate779inter3), .O(gate779inter10));
  nor2  gate2443(.a(gate779inter10), .b(gate779inter9), .O(gate779inter11));
  nor2  gate2444(.a(gate779inter11), .b(gate779inter6), .O(gate779inter12));
  nand2 gate2445(.a(gate779inter12), .b(gate779inter1), .O(N2881));
nand2 gate780( .a(N2777), .b(N2778), .O(N2882) );
nand2 gate781( .a(N2775), .b(N2776), .O(N2885) );
nand2 gate782( .a(N2781), .b(N2782), .O(N2888) );

  xor2  gate2656(.a(N2784), .b(N2783), .O(gate783inter0));
  nand2 gate2657(.a(gate783inter0), .b(s_198), .O(gate783inter1));
  and2  gate2658(.a(N2784), .b(N2783), .O(gate783inter2));
  inv1  gate2659(.a(s_198), .O(gate783inter3));
  inv1  gate2660(.a(s_199), .O(gate783inter4));
  nand2 gate2661(.a(gate783inter4), .b(gate783inter3), .O(gate783inter5));
  nor2  gate2662(.a(gate783inter5), .b(gate783inter2), .O(gate783inter6));
  inv1  gate2663(.a(N2783), .O(gate783inter7));
  inv1  gate2664(.a(N2784), .O(gate783inter8));
  nand2 gate2665(.a(gate783inter8), .b(gate783inter7), .O(gate783inter9));
  nand2 gate2666(.a(s_199), .b(gate783inter3), .O(gate783inter10));
  nor2  gate2667(.a(gate783inter10), .b(gate783inter9), .O(gate783inter11));
  nor2  gate2668(.a(gate783inter11), .b(gate783inter6), .O(gate783inter12));
  nand2 gate2669(.a(gate783inter12), .b(gate783inter1), .O(N2891));
and2 gate784( .a(N2607), .b(N2729), .O(N2894) );
and2 gate785( .a(N2608), .b(N2729), .O(N2895) );
and2 gate786( .a(N2609), .b(N2729), .O(N2896) );
and2 gate787( .a(N2610), .b(N2729), .O(N2897) );
or2 gate788( .a(N2789), .b(N2611), .O(N2898) );
or2 gate789( .a(N2790), .b(N2612), .O(N2899) );
and2 gate790( .a(N2791), .b(N1037), .O(N2900) );
and2 gate791( .a(N2792), .b(N1037), .O(N2901) );
or2 gate792( .a(N2809), .b(N2631), .O(N2914) );
or2 gate793( .a(N2810), .b(N2632), .O(N2915) );
and2 gate794( .a(N2811), .b(N1070), .O(N2916) );
and2 gate795( .a(N2812), .b(N1070), .O(N2917) );
and2 gate796( .a(N2633), .b(N2738), .O(N2918) );
and2 gate797( .a(N2634), .b(N2738), .O(N2919) );
and2 gate798( .a(N2635), .b(N2738), .O(N2920) );
and2 gate799( .a(N2636), .b(N2738), .O(N2921) );
buf1 gate800( .a(N2817), .O(N2925) );
and3 gate801( .a(N2829), .b(N2830), .c(N1302), .O(N2931) );
and3 gate802( .a(N2681), .b(N2421), .c(N2837), .O(N2938) );
and3 gate803( .a(N2417), .b(N2684), .c(N2838), .O(N2939) );
nand2 gate804( .a(N2469), .b(N2880), .O(N2963) );
inv1 gate805( .a(N2841), .O(N2970) );
inv1 gate806( .a(N2826), .O(N2971) );
inv1 gate807( .a(N2894), .O(N2972) );
inv1 gate808( .a(N2895), .O(N2975) );
inv1 gate809( .a(N2896), .O(N2978) );
inv1 gate810( .a(N2897), .O(N2981) );
and2 gate811( .a(N2898), .b(N1037), .O(N2984) );
and2 gate812( .a(N2899), .b(N1037), .O(N2985) );
inv1 gate813( .a(N2900), .O(N2986) );
inv1 gate814( .a(N2901), .O(N2989) );
inv1 gate815( .a(N2796), .O(N2992) );
buf1 gate816( .a(N2800), .O(N2995) );
buf1 gate817( .a(N2800), .O(N2998) );
buf1 gate818( .a(N2806), .O(N3001) );
buf1 gate819( .a(N2806), .O(N3004) );
and2 gate820( .a(N574), .b(N2820), .O(N3007) );
and2 gate821( .a(N2914), .b(N1070), .O(N3008) );
and2 gate822( .a(N2915), .b(N1070), .O(N3009) );
inv1 gate823( .a(N2916), .O(N3010) );
inv1 gate824( .a(N2917), .O(N3013) );
inv1 gate825( .a(N2918), .O(N3016) );
inv1 gate826( .a(N2919), .O(N3019) );
inv1 gate827( .a(N2920), .O(N3022) );
inv1 gate828( .a(N2921), .O(N3025) );
inv1 gate829( .a(N2817), .O(N3028) );
and2 gate830( .a(N574), .b(N2831), .O(N3029) );
inv1 gate831( .a(N2820), .O(N3030) );
and2 gate832( .a(N578), .b(N2820), .O(N3035) );
and2 gate833( .a(N655), .b(N2820), .O(N3036) );
and2 gate834( .a(N659), .b(N2820), .O(N3037) );
buf1 gate835( .a(N2931), .O(N3038) );
inv1 gate836( .a(N2831), .O(N3039) );
and2 gate837( .a(N578), .b(N2831), .O(N3044) );
and2 gate838( .a(N655), .b(N2831), .O(N3045) );
and2 gate839( .a(N659), .b(N2831), .O(N3046) );
nor2 gate840( .a(N2938), .b(N2839), .O(N3047) );
nor2 gate841( .a(N2939), .b(N2840), .O(N3048) );
inv1 gate842( .a(N2888), .O(N3049) );
inv1 gate843( .a(N2844), .O(N3050) );
and2 gate844( .a(N663), .b(N2844), .O(N3053) );
and2 gate845( .a(N667), .b(N2844), .O(N3054) );
and2 gate846( .a(N671), .b(N2844), .O(N3055) );
and2 gate847( .a(N675), .b(N2844), .O(N3056) );
and2 gate848( .a(N679), .b(N2854), .O(N3057) );
and2 gate849( .a(N683), .b(N2854), .O(N3058) );
and2 gate850( .a(N687), .b(N2854), .O(N3059) );
and2 gate851( .a(N705), .b(N2854), .O(N3060) );
inv1 gate852( .a(N2859), .O(N3061) );
and2 gate853( .a(N663), .b(N2859), .O(N3064) );
and2 gate854( .a(N667), .b(N2859), .O(N3065) );
and2 gate855( .a(N671), .b(N2859), .O(N3066) );
and2 gate856( .a(N675), .b(N2859), .O(N3067) );
and2 gate857( .a(N679), .b(N2869), .O(N3068) );
and2 gate858( .a(N683), .b(N2869), .O(N3069) );
and2 gate859( .a(N687), .b(N2869), .O(N3070) );
and2 gate860( .a(N705), .b(N2869), .O(N3071) );
inv1 gate861( .a(N2874), .O(N3072) );
inv1 gate862( .a(N2877), .O(N3073) );
inv1 gate863( .a(N2882), .O(N3074) );
inv1 gate864( .a(N2885), .O(N3075) );
nand2 gate865( .a(N2881), .b(N2963), .O(N3076) );
inv1 gate866( .a(N2931), .O(N3079) );
inv1 gate867( .a(N2984), .O(N3088) );
inv1 gate868( .a(N2985), .O(N3091) );
inv1 gate869( .a(N3008), .O(N3110) );
inv1 gate870( .a(N3009), .O(N3113) );
and2 gate871( .a(N3055), .b(N1190), .O(N3137) );
and2 gate872( .a(N3056), .b(N1190), .O(N3140) );
and2 gate873( .a(N3057), .b(N2761), .O(N3143) );
and2 gate874( .a(N3058), .b(N2761), .O(N3146) );
and2 gate875( .a(N3059), .b(N2761), .O(N3149) );
and2 gate876( .a(N3060), .b(N2761), .O(N3152) );
and2 gate877( .a(N3066), .b(N1195), .O(N3157) );
and2 gate878( .a(N3067), .b(N1195), .O(N3160) );
and2 gate879( .a(N3068), .b(N2766), .O(N3163) );
and2 gate880( .a(N3069), .b(N2766), .O(N3166) );
and2 gate881( .a(N3070), .b(N2766), .O(N3169) );
and2 gate882( .a(N3071), .b(N2766), .O(N3172) );

  xor2  gate1466(.a(N3072), .b(N2877), .O(gate883inter0));
  nand2 gate1467(.a(gate883inter0), .b(s_28), .O(gate883inter1));
  and2  gate1468(.a(N3072), .b(N2877), .O(gate883inter2));
  inv1  gate1469(.a(s_28), .O(gate883inter3));
  inv1  gate1470(.a(s_29), .O(gate883inter4));
  nand2 gate1471(.a(gate883inter4), .b(gate883inter3), .O(gate883inter5));
  nor2  gate1472(.a(gate883inter5), .b(gate883inter2), .O(gate883inter6));
  inv1  gate1473(.a(N2877), .O(gate883inter7));
  inv1  gate1474(.a(N3072), .O(gate883inter8));
  nand2 gate1475(.a(gate883inter8), .b(gate883inter7), .O(gate883inter9));
  nand2 gate1476(.a(s_29), .b(gate883inter3), .O(gate883inter10));
  nor2  gate1477(.a(gate883inter10), .b(gate883inter9), .O(gate883inter11));
  nor2  gate1478(.a(gate883inter11), .b(gate883inter6), .O(gate883inter12));
  nand2 gate1479(.a(gate883inter12), .b(gate883inter1), .O(N3175));
nand2 gate884( .a(N2874), .b(N3073), .O(N3176) );

  xor2  gate1326(.a(N3074), .b(N2885), .O(gate885inter0));
  nand2 gate1327(.a(gate885inter0), .b(s_8), .O(gate885inter1));
  and2  gate1328(.a(N3074), .b(N2885), .O(gate885inter2));
  inv1  gate1329(.a(s_8), .O(gate885inter3));
  inv1  gate1330(.a(s_9), .O(gate885inter4));
  nand2 gate1331(.a(gate885inter4), .b(gate885inter3), .O(gate885inter5));
  nor2  gate1332(.a(gate885inter5), .b(gate885inter2), .O(gate885inter6));
  inv1  gate1333(.a(N2885), .O(gate885inter7));
  inv1  gate1334(.a(N3074), .O(gate885inter8));
  nand2 gate1335(.a(gate885inter8), .b(gate885inter7), .O(gate885inter9));
  nand2 gate1336(.a(s_9), .b(gate885inter3), .O(gate885inter10));
  nor2  gate1337(.a(gate885inter10), .b(gate885inter9), .O(gate885inter11));
  nor2  gate1338(.a(gate885inter11), .b(gate885inter6), .O(gate885inter12));
  nand2 gate1339(.a(gate885inter12), .b(gate885inter1), .O(N3177));

  xor2  gate1424(.a(N3075), .b(N2882), .O(gate886inter0));
  nand2 gate1425(.a(gate886inter0), .b(s_22), .O(gate886inter1));
  and2  gate1426(.a(N3075), .b(N2882), .O(gate886inter2));
  inv1  gate1427(.a(s_22), .O(gate886inter3));
  inv1  gate1428(.a(s_23), .O(gate886inter4));
  nand2 gate1429(.a(gate886inter4), .b(gate886inter3), .O(gate886inter5));
  nor2  gate1430(.a(gate886inter5), .b(gate886inter2), .O(gate886inter6));
  inv1  gate1431(.a(N2882), .O(gate886inter7));
  inv1  gate1432(.a(N3075), .O(gate886inter8));
  nand2 gate1433(.a(gate886inter8), .b(gate886inter7), .O(gate886inter9));
  nand2 gate1434(.a(s_23), .b(gate886inter3), .O(gate886inter10));
  nor2  gate1435(.a(gate886inter10), .b(gate886inter9), .O(gate886inter11));
  nor2  gate1436(.a(gate886inter11), .b(gate886inter6), .O(gate886inter12));
  nand2 gate1437(.a(gate886inter12), .b(gate886inter1), .O(N3178));

  xor2  gate1634(.a(N3047), .b(N3048), .O(gate887inter0));
  nand2 gate1635(.a(gate887inter0), .b(s_52), .O(gate887inter1));
  and2  gate1636(.a(N3047), .b(N3048), .O(gate887inter2));
  inv1  gate1637(.a(s_52), .O(gate887inter3));
  inv1  gate1638(.a(s_53), .O(gate887inter4));
  nand2 gate1639(.a(gate887inter4), .b(gate887inter3), .O(gate887inter5));
  nor2  gate1640(.a(gate887inter5), .b(gate887inter2), .O(gate887inter6));
  inv1  gate1641(.a(N3048), .O(gate887inter7));
  inv1  gate1642(.a(N3047), .O(gate887inter8));
  nand2 gate1643(.a(gate887inter8), .b(gate887inter7), .O(gate887inter9));
  nand2 gate1644(.a(s_53), .b(gate887inter3), .O(gate887inter10));
  nor2  gate1645(.a(gate887inter10), .b(gate887inter9), .O(gate887inter11));
  nor2  gate1646(.a(gate887inter11), .b(gate887inter6), .O(gate887inter12));
  nand2 gate1647(.a(gate887inter12), .b(gate887inter1), .O(N3180));
inv1 gate888( .a(N2995), .O(N3187) );
inv1 gate889( .a(N2998), .O(N3188) );
inv1 gate890( .a(N3001), .O(N3189) );
inv1 gate891( .a(N3004), .O(N3190) );
and3 gate892( .a(N2796), .b(N2613), .c(N2995), .O(N3191) );
and3 gate893( .a(N2992), .b(N2793), .c(N2998), .O(N3192) );
and3 gate894( .a(N2624), .b(N2368), .c(N3001), .O(N3193) );
and3 gate895( .a(N2803), .b(N2621), .c(N3004), .O(N3194) );

  xor2  gate2964(.a(N2375), .b(N3076), .O(gate896inter0));
  nand2 gate2965(.a(gate896inter0), .b(s_242), .O(gate896inter1));
  and2  gate2966(.a(N2375), .b(N3076), .O(gate896inter2));
  inv1  gate2967(.a(s_242), .O(gate896inter3));
  inv1  gate2968(.a(s_243), .O(gate896inter4));
  nand2 gate2969(.a(gate896inter4), .b(gate896inter3), .O(gate896inter5));
  nor2  gate2970(.a(gate896inter5), .b(gate896inter2), .O(gate896inter6));
  inv1  gate2971(.a(N3076), .O(gate896inter7));
  inv1  gate2972(.a(N2375), .O(gate896inter8));
  nand2 gate2973(.a(gate896inter8), .b(gate896inter7), .O(gate896inter9));
  nand2 gate2974(.a(s_243), .b(gate896inter3), .O(gate896inter10));
  nor2  gate2975(.a(gate896inter10), .b(gate896inter9), .O(gate896inter11));
  nor2  gate2976(.a(gate896inter11), .b(gate896inter6), .O(gate896inter12));
  nand2 gate2977(.a(gate896inter12), .b(gate896inter1), .O(N3195));
inv1 gate897( .a(N3076), .O(N3196) );
and2 gate898( .a(N687), .b(N3030), .O(N3197) );
and2 gate899( .a(N687), .b(N3039), .O(N3208) );
and2 gate900( .a(N705), .b(N3030), .O(N3215) );
and2 gate901( .a(N711), .b(N3030), .O(N3216) );
and2 gate902( .a(N715), .b(N3030), .O(N3217) );
and2 gate903( .a(N705), .b(N3039), .O(N3218) );
and2 gate904( .a(N711), .b(N3039), .O(N3219) );
and2 gate905( .a(N715), .b(N3039), .O(N3220) );
and2 gate906( .a(N719), .b(N3050), .O(N3222) );
and2 gate907( .a(N723), .b(N3050), .O(N3223) );
and2 gate908( .a(N719), .b(N3061), .O(N3230) );
and2 gate909( .a(N723), .b(N3061), .O(N3231) );

  xor2  gate2418(.a(N3176), .b(N3175), .O(gate910inter0));
  nand2 gate2419(.a(gate910inter0), .b(s_164), .O(gate910inter1));
  and2  gate2420(.a(N3176), .b(N3175), .O(gate910inter2));
  inv1  gate2421(.a(s_164), .O(gate910inter3));
  inv1  gate2422(.a(s_165), .O(gate910inter4));
  nand2 gate2423(.a(gate910inter4), .b(gate910inter3), .O(gate910inter5));
  nor2  gate2424(.a(gate910inter5), .b(gate910inter2), .O(gate910inter6));
  inv1  gate2425(.a(N3175), .O(gate910inter7));
  inv1  gate2426(.a(N3176), .O(gate910inter8));
  nand2 gate2427(.a(gate910inter8), .b(gate910inter7), .O(gate910inter9));
  nand2 gate2428(.a(s_165), .b(gate910inter3), .O(gate910inter10));
  nor2  gate2429(.a(gate910inter10), .b(gate910inter9), .O(gate910inter11));
  nor2  gate2430(.a(gate910inter11), .b(gate910inter6), .O(gate910inter12));
  nand2 gate2431(.a(gate910inter12), .b(gate910inter1), .O(N3238));
nand2 gate911( .a(N3177), .b(N3178), .O(N3241) );
buf1 gate912( .a(N2981), .O(N3244) );
buf1 gate913( .a(N2978), .O(N3247) );
buf1 gate914( .a(N2975), .O(N3250) );
buf1 gate915( .a(N2972), .O(N3253) );
buf1 gate916( .a(N2989), .O(N3256) );
buf1 gate917( .a(N2986), .O(N3259) );
buf1 gate918( .a(N3025), .O(N3262) );
buf1 gate919( .a(N3022), .O(N3265) );
buf1 gate920( .a(N3019), .O(N3268) );
buf1 gate921( .a(N3016), .O(N3271) );
buf1 gate922( .a(N3013), .O(N3274) );
buf1 gate923( .a(N3010), .O(N3277) );
and3 gate924( .a(N2793), .b(N2796), .c(N3187), .O(N3281) );
and3 gate925( .a(N2613), .b(N2992), .c(N3188), .O(N3282) );
and3 gate926( .a(N2621), .b(N2624), .c(N3189), .O(N3283) );
and3 gate927( .a(N2368), .b(N2803), .c(N3190), .O(N3284) );

  xor2  gate2838(.a(N3196), .b(N2210), .O(gate928inter0));
  nand2 gate2839(.a(gate928inter0), .b(s_224), .O(gate928inter1));
  and2  gate2840(.a(N3196), .b(N2210), .O(gate928inter2));
  inv1  gate2841(.a(s_224), .O(gate928inter3));
  inv1  gate2842(.a(s_225), .O(gate928inter4));
  nand2 gate2843(.a(gate928inter4), .b(gate928inter3), .O(gate928inter5));
  nor2  gate2844(.a(gate928inter5), .b(gate928inter2), .O(gate928inter6));
  inv1  gate2845(.a(N2210), .O(gate928inter7));
  inv1  gate2846(.a(N3196), .O(gate928inter8));
  nand2 gate2847(.a(gate928inter8), .b(gate928inter7), .O(gate928inter9));
  nand2 gate2848(.a(s_225), .b(gate928inter3), .O(gate928inter10));
  nor2  gate2849(.a(gate928inter10), .b(gate928inter9), .O(gate928inter11));
  nor2  gate2850(.a(gate928inter11), .b(gate928inter6), .O(gate928inter12));
  nand2 gate2851(.a(gate928inter12), .b(gate928inter1), .O(N3286));
or2 gate929( .a(N3197), .b(N3007), .O(N3288) );

  xor2  gate1662(.a(N3049), .b(N3180), .O(gate930inter0));
  nand2 gate1663(.a(gate930inter0), .b(s_56), .O(gate930inter1));
  and2  gate1664(.a(N3049), .b(N3180), .O(gate930inter2));
  inv1  gate1665(.a(s_56), .O(gate930inter3));
  inv1  gate1666(.a(s_57), .O(gate930inter4));
  nand2 gate1667(.a(gate930inter4), .b(gate930inter3), .O(gate930inter5));
  nor2  gate1668(.a(gate930inter5), .b(gate930inter2), .O(gate930inter6));
  inv1  gate1669(.a(N3180), .O(gate930inter7));
  inv1  gate1670(.a(N3049), .O(gate930inter8));
  nand2 gate1671(.a(gate930inter8), .b(gate930inter7), .O(gate930inter9));
  nand2 gate1672(.a(s_57), .b(gate930inter3), .O(gate930inter10));
  nor2  gate1673(.a(gate930inter10), .b(gate930inter9), .O(gate930inter11));
  nor2  gate1674(.a(gate930inter11), .b(gate930inter6), .O(gate930inter12));
  nand2 gate1675(.a(gate930inter12), .b(gate930inter1), .O(N3289));
and2 gate931( .a(N3152), .b(N2981), .O(N3291) );
and2 gate932( .a(N3149), .b(N2978), .O(N3293) );
and2 gate933( .a(N3146), .b(N2975), .O(N3295) );
and2 gate934( .a(N2972), .b(N3143), .O(N3296) );
and2 gate935( .a(N3140), .b(N2989), .O(N3299) );
and2 gate936( .a(N3137), .b(N2986), .O(N3301) );
or2 gate937( .a(N3208), .b(N3029), .O(N3302) );
and2 gate938( .a(N3172), .b(N3025), .O(N3304) );
and2 gate939( .a(N3169), .b(N3022), .O(N3306) );
and2 gate940( .a(N3166), .b(N3019), .O(N3308) );
and2 gate941( .a(N3016), .b(N3163), .O(N3309) );
and2 gate942( .a(N3160), .b(N3013), .O(N3312) );
and2 gate943( .a(N3157), .b(N3010), .O(N3314) );
or2 gate944( .a(N3215), .b(N3035), .O(N3315) );
or2 gate945( .a(N3216), .b(N3036), .O(N3318) );
or2 gate946( .a(N3217), .b(N3037), .O(N3321) );
or2 gate947( .a(N3218), .b(N3044), .O(N3324) );
or2 gate948( .a(N3219), .b(N3045), .O(N3327) );
or2 gate949( .a(N3220), .b(N3046), .O(N3330) );
inv1 gate950( .a(N3180), .O(N3333) );
or2 gate951( .a(N3222), .b(N3053), .O(N3334) );
or2 gate952( .a(N3223), .b(N3054), .O(N3335) );
or2 gate953( .a(N3230), .b(N3064), .O(N3336) );
or2 gate954( .a(N3231), .b(N3065), .O(N3337) );
buf1 gate955( .a(N3152), .O(N3340) );
buf1 gate956( .a(N3149), .O(N3344) );
buf1 gate957( .a(N3146), .O(N3348) );
buf1 gate958( .a(N3143), .O(N3352) );
buf1 gate959( .a(N3140), .O(N3356) );
buf1 gate960( .a(N3137), .O(N3360) );
buf1 gate961( .a(N3091), .O(N3364) );
buf1 gate962( .a(N3088), .O(N3367) );
buf1 gate963( .a(N3172), .O(N3370) );
buf1 gate964( .a(N3169), .O(N3374) );
buf1 gate965( .a(N3166), .O(N3378) );
buf1 gate966( .a(N3163), .O(N3382) );
buf1 gate967( .a(N3160), .O(N3386) );
buf1 gate968( .a(N3157), .O(N3390) );
buf1 gate969( .a(N3113), .O(N3394) );
buf1 gate970( .a(N3110), .O(N3397) );

  xor2  gate2544(.a(N3286), .b(N3195), .O(gate971inter0));
  nand2 gate2545(.a(gate971inter0), .b(s_182), .O(gate971inter1));
  and2  gate2546(.a(N3286), .b(N3195), .O(gate971inter2));
  inv1  gate2547(.a(s_182), .O(gate971inter3));
  inv1  gate2548(.a(s_183), .O(gate971inter4));
  nand2 gate2549(.a(gate971inter4), .b(gate971inter3), .O(gate971inter5));
  nor2  gate2550(.a(gate971inter5), .b(gate971inter2), .O(gate971inter6));
  inv1  gate2551(.a(N3195), .O(gate971inter7));
  inv1  gate2552(.a(N3286), .O(gate971inter8));
  nand2 gate2553(.a(gate971inter8), .b(gate971inter7), .O(gate971inter9));
  nand2 gate2554(.a(s_183), .b(gate971inter3), .O(gate971inter10));
  nor2  gate2555(.a(gate971inter10), .b(gate971inter9), .O(gate971inter11));
  nor2  gate2556(.a(gate971inter11), .b(gate971inter6), .O(gate971inter12));
  nand2 gate2557(.a(gate971inter12), .b(gate971inter1), .O(N3400));
nor2 gate972( .a(N3281), .b(N3191), .O(N3401) );
nor2 gate973( .a(N3282), .b(N3192), .O(N3402) );
nor2 gate974( .a(N3283), .b(N3193), .O(N3403) );

  xor2  gate2586(.a(N3194), .b(N3284), .O(gate975inter0));
  nand2 gate2587(.a(gate975inter0), .b(s_188), .O(gate975inter1));
  and2  gate2588(.a(N3194), .b(N3284), .O(gate975inter2));
  inv1  gate2589(.a(s_188), .O(gate975inter3));
  inv1  gate2590(.a(s_189), .O(gate975inter4));
  nand2 gate2591(.a(gate975inter4), .b(gate975inter3), .O(gate975inter5));
  nor2  gate2592(.a(gate975inter5), .b(gate975inter2), .O(gate975inter6));
  inv1  gate2593(.a(N3284), .O(gate975inter7));
  inv1  gate2594(.a(N3194), .O(gate975inter8));
  nand2 gate2595(.a(gate975inter8), .b(gate975inter7), .O(gate975inter9));
  nand2 gate2596(.a(s_189), .b(gate975inter3), .O(gate975inter10));
  nor2  gate2597(.a(gate975inter10), .b(gate975inter9), .O(gate975inter11));
  nor2  gate2598(.a(gate975inter11), .b(gate975inter6), .O(gate975inter12));
  nand2 gate2599(.a(gate975inter12), .b(gate975inter1), .O(N3404));
inv1 gate976( .a(N3238), .O(N3405) );
inv1 gate977( .a(N3241), .O(N3406) );
and2 gate978( .a(N3288), .b(N1836), .O(N3409) );

  xor2  gate2950(.a(N3333), .b(N2888), .O(gate979inter0));
  nand2 gate2951(.a(gate979inter0), .b(s_240), .O(gate979inter1));
  and2  gate2952(.a(N3333), .b(N2888), .O(gate979inter2));
  inv1  gate2953(.a(s_240), .O(gate979inter3));
  inv1  gate2954(.a(s_241), .O(gate979inter4));
  nand2 gate2955(.a(gate979inter4), .b(gate979inter3), .O(gate979inter5));
  nor2  gate2956(.a(gate979inter5), .b(gate979inter2), .O(gate979inter6));
  inv1  gate2957(.a(N2888), .O(gate979inter7));
  inv1  gate2958(.a(N3333), .O(gate979inter8));
  nand2 gate2959(.a(gate979inter8), .b(gate979inter7), .O(gate979inter9));
  nand2 gate2960(.a(s_241), .b(gate979inter3), .O(gate979inter10));
  nor2  gate2961(.a(gate979inter10), .b(gate979inter9), .O(gate979inter11));
  nor2  gate2962(.a(gate979inter11), .b(gate979inter6), .O(gate979inter12));
  nand2 gate2963(.a(gate979inter12), .b(gate979inter1), .O(N3410));
inv1 gate980( .a(N3244), .O(N3412) );
inv1 gate981( .a(N3247), .O(N3414) );
inv1 gate982( .a(N3250), .O(N3416) );
inv1 gate983( .a(N3253), .O(N3418) );
inv1 gate984( .a(N3256), .O(N3420) );
inv1 gate985( .a(N3259), .O(N3422) );
and2 gate986( .a(N3302), .b(N1836), .O(N3428) );
inv1 gate987( .a(N3262), .O(N3430) );
inv1 gate988( .a(N3265), .O(N3432) );
inv1 gate989( .a(N3268), .O(N3434) );
inv1 gate990( .a(N3271), .O(N3436) );
inv1 gate991( .a(N3274), .O(N3438) );
inv1 gate992( .a(N3277), .O(N3440) );
and2 gate993( .a(N3334), .b(N1190), .O(N3450) );
and2 gate994( .a(N3335), .b(N1190), .O(N3453) );
and2 gate995( .a(N3336), .b(N1195), .O(N3456) );
and2 gate996( .a(N3337), .b(N1195), .O(N3459) );
and2 gate997( .a(N3400), .b(N533), .O(N3478) );
and2 gate998( .a(N3318), .b(N2128), .O(N3479) );
and2 gate999( .a(N3315), .b(N1841), .O(N3480) );
nand2 gate1000( .a(N3410), .b(N3289), .O(N3481) );
inv1 gate1001( .a(N3340), .O(N3482) );

  xor2  gate3020(.a(N3412), .b(N3340), .O(gate1002inter0));
  nand2 gate3021(.a(gate1002inter0), .b(s_250), .O(gate1002inter1));
  and2  gate3022(.a(N3412), .b(N3340), .O(gate1002inter2));
  inv1  gate3023(.a(s_250), .O(gate1002inter3));
  inv1  gate3024(.a(s_251), .O(gate1002inter4));
  nand2 gate3025(.a(gate1002inter4), .b(gate1002inter3), .O(gate1002inter5));
  nor2  gate3026(.a(gate1002inter5), .b(gate1002inter2), .O(gate1002inter6));
  inv1  gate3027(.a(N3340), .O(gate1002inter7));
  inv1  gate3028(.a(N3412), .O(gate1002inter8));
  nand2 gate3029(.a(gate1002inter8), .b(gate1002inter7), .O(gate1002inter9));
  nand2 gate3030(.a(s_251), .b(gate1002inter3), .O(gate1002inter10));
  nor2  gate3031(.a(gate1002inter10), .b(gate1002inter9), .O(gate1002inter11));
  nor2  gate3032(.a(gate1002inter11), .b(gate1002inter6), .O(gate1002inter12));
  nand2 gate3033(.a(gate1002inter12), .b(gate1002inter1), .O(N3483));
inv1 gate1003( .a(N3344), .O(N3484) );

  xor2  gate2138(.a(N3414), .b(N3344), .O(gate1004inter0));
  nand2 gate2139(.a(gate1004inter0), .b(s_124), .O(gate1004inter1));
  and2  gate2140(.a(N3414), .b(N3344), .O(gate1004inter2));
  inv1  gate2141(.a(s_124), .O(gate1004inter3));
  inv1  gate2142(.a(s_125), .O(gate1004inter4));
  nand2 gate2143(.a(gate1004inter4), .b(gate1004inter3), .O(gate1004inter5));
  nor2  gate2144(.a(gate1004inter5), .b(gate1004inter2), .O(gate1004inter6));
  inv1  gate2145(.a(N3344), .O(gate1004inter7));
  inv1  gate2146(.a(N3414), .O(gate1004inter8));
  nand2 gate2147(.a(gate1004inter8), .b(gate1004inter7), .O(gate1004inter9));
  nand2 gate2148(.a(s_125), .b(gate1004inter3), .O(gate1004inter10));
  nor2  gate2149(.a(gate1004inter10), .b(gate1004inter9), .O(gate1004inter11));
  nor2  gate2150(.a(gate1004inter11), .b(gate1004inter6), .O(gate1004inter12));
  nand2 gate2151(.a(gate1004inter12), .b(gate1004inter1), .O(N3485));
inv1 gate1005( .a(N3348), .O(N3486) );
nand2 gate1006( .a(N3348), .b(N3416), .O(N3487) );
inv1 gate1007( .a(N3352), .O(N3488) );
nand2 gate1008( .a(N3352), .b(N3418), .O(N3489) );
inv1 gate1009( .a(N3356), .O(N3490) );
nand2 gate1010( .a(N3356), .b(N3420), .O(N3491) );
inv1 gate1011( .a(N3360), .O(N3492) );

  xor2  gate2880(.a(N3422), .b(N3360), .O(gate1012inter0));
  nand2 gate2881(.a(gate1012inter0), .b(s_230), .O(gate1012inter1));
  and2  gate2882(.a(N3422), .b(N3360), .O(gate1012inter2));
  inv1  gate2883(.a(s_230), .O(gate1012inter3));
  inv1  gate2884(.a(s_231), .O(gate1012inter4));
  nand2 gate2885(.a(gate1012inter4), .b(gate1012inter3), .O(gate1012inter5));
  nor2  gate2886(.a(gate1012inter5), .b(gate1012inter2), .O(gate1012inter6));
  inv1  gate2887(.a(N3360), .O(gate1012inter7));
  inv1  gate2888(.a(N3422), .O(gate1012inter8));
  nand2 gate2889(.a(gate1012inter8), .b(gate1012inter7), .O(gate1012inter9));
  nand2 gate2890(.a(s_231), .b(gate1012inter3), .O(gate1012inter10));
  nor2  gate2891(.a(gate1012inter10), .b(gate1012inter9), .O(gate1012inter11));
  nor2  gate2892(.a(gate1012inter11), .b(gate1012inter6), .O(gate1012inter12));
  nand2 gate2893(.a(gate1012inter12), .b(gate1012inter1), .O(N3493));
inv1 gate1013( .a(N3364), .O(N3494) );
inv1 gate1014( .a(N3367), .O(N3496) );
and2 gate1015( .a(N3321), .b(N2135), .O(N3498) );
and2 gate1016( .a(N3327), .b(N2128), .O(N3499) );
and2 gate1017( .a(N3324), .b(N1841), .O(N3500) );
inv1 gate1018( .a(N3370), .O(N3501) );
nand2 gate1019( .a(N3370), .b(N3430), .O(N3502) );
inv1 gate1020( .a(N3374), .O(N3503) );
nand2 gate1021( .a(N3374), .b(N3432), .O(N3504) );
inv1 gate1022( .a(N3378), .O(N3505) );

  xor2  gate2166(.a(N3434), .b(N3378), .O(gate1023inter0));
  nand2 gate2167(.a(gate1023inter0), .b(s_128), .O(gate1023inter1));
  and2  gate2168(.a(N3434), .b(N3378), .O(gate1023inter2));
  inv1  gate2169(.a(s_128), .O(gate1023inter3));
  inv1  gate2170(.a(s_129), .O(gate1023inter4));
  nand2 gate2171(.a(gate1023inter4), .b(gate1023inter3), .O(gate1023inter5));
  nor2  gate2172(.a(gate1023inter5), .b(gate1023inter2), .O(gate1023inter6));
  inv1  gate2173(.a(N3378), .O(gate1023inter7));
  inv1  gate2174(.a(N3434), .O(gate1023inter8));
  nand2 gate2175(.a(gate1023inter8), .b(gate1023inter7), .O(gate1023inter9));
  nand2 gate2176(.a(s_129), .b(gate1023inter3), .O(gate1023inter10));
  nor2  gate2177(.a(gate1023inter10), .b(gate1023inter9), .O(gate1023inter11));
  nor2  gate2178(.a(gate1023inter11), .b(gate1023inter6), .O(gate1023inter12));
  nand2 gate2179(.a(gate1023inter12), .b(gate1023inter1), .O(N3506));
inv1 gate1024( .a(N3382), .O(N3507) );

  xor2  gate1312(.a(N3436), .b(N3382), .O(gate1025inter0));
  nand2 gate1313(.a(gate1025inter0), .b(s_6), .O(gate1025inter1));
  and2  gate1314(.a(N3436), .b(N3382), .O(gate1025inter2));
  inv1  gate1315(.a(s_6), .O(gate1025inter3));
  inv1  gate1316(.a(s_7), .O(gate1025inter4));
  nand2 gate1317(.a(gate1025inter4), .b(gate1025inter3), .O(gate1025inter5));
  nor2  gate1318(.a(gate1025inter5), .b(gate1025inter2), .O(gate1025inter6));
  inv1  gate1319(.a(N3382), .O(gate1025inter7));
  inv1  gate1320(.a(N3436), .O(gate1025inter8));
  nand2 gate1321(.a(gate1025inter8), .b(gate1025inter7), .O(gate1025inter9));
  nand2 gate1322(.a(s_7), .b(gate1025inter3), .O(gate1025inter10));
  nor2  gate1323(.a(gate1025inter10), .b(gate1025inter9), .O(gate1025inter11));
  nor2  gate1324(.a(gate1025inter11), .b(gate1025inter6), .O(gate1025inter12));
  nand2 gate1325(.a(gate1025inter12), .b(gate1025inter1), .O(N3508));
inv1 gate1026( .a(N3386), .O(N3509) );
nand2 gate1027( .a(N3386), .b(N3438), .O(N3510) );
inv1 gate1028( .a(N3390), .O(N3511) );
nand2 gate1029( .a(N3390), .b(N3440), .O(N3512) );
inv1 gate1030( .a(N3394), .O(N3513) );
inv1 gate1031( .a(N3397), .O(N3515) );
and2 gate1032( .a(N3330), .b(N2135), .O(N3517) );
nand2 gate1033( .a(N3402), .b(N3401), .O(N3522) );

  xor2  gate1396(.a(N3403), .b(N3404), .O(gate1034inter0));
  nand2 gate1397(.a(gate1034inter0), .b(s_18), .O(gate1034inter1));
  and2  gate1398(.a(N3403), .b(N3404), .O(gate1034inter2));
  inv1  gate1399(.a(s_18), .O(gate1034inter3));
  inv1  gate1400(.a(s_19), .O(gate1034inter4));
  nand2 gate1401(.a(gate1034inter4), .b(gate1034inter3), .O(gate1034inter5));
  nor2  gate1402(.a(gate1034inter5), .b(gate1034inter2), .O(gate1034inter6));
  inv1  gate1403(.a(N3404), .O(gate1034inter7));
  inv1  gate1404(.a(N3403), .O(gate1034inter8));
  nand2 gate1405(.a(gate1034inter8), .b(gate1034inter7), .O(gate1034inter9));
  nand2 gate1406(.a(s_19), .b(gate1034inter3), .O(gate1034inter10));
  nor2  gate1407(.a(gate1034inter10), .b(gate1034inter9), .O(gate1034inter11));
  nor2  gate1408(.a(gate1034inter11), .b(gate1034inter6), .O(gate1034inter12));
  nand2 gate1409(.a(gate1034inter12), .b(gate1034inter1), .O(N3525));
buf1 gate1035( .a(N3318), .O(N3528) );
buf1 gate1036( .a(N3315), .O(N3531) );
buf1 gate1037( .a(N3321), .O(N3534) );
buf1 gate1038( .a(N3327), .O(N3537) );
buf1 gate1039( .a(N3324), .O(N3540) );
buf1 gate1040( .a(N3330), .O(N3543) );
or2 gate1041( .a(N3478), .b(N1813), .O(N3546) );
inv1 gate1042( .a(N3481), .O(N3551) );
nand2 gate1043( .a(N3244), .b(N3482), .O(N3552) );

  xor2  gate1270(.a(N3484), .b(N3247), .O(gate1044inter0));
  nand2 gate1271(.a(gate1044inter0), .b(s_0), .O(gate1044inter1));
  and2  gate1272(.a(N3484), .b(N3247), .O(gate1044inter2));
  inv1  gate1273(.a(s_0), .O(gate1044inter3));
  inv1  gate1274(.a(s_1), .O(gate1044inter4));
  nand2 gate1275(.a(gate1044inter4), .b(gate1044inter3), .O(gate1044inter5));
  nor2  gate1276(.a(gate1044inter5), .b(gate1044inter2), .O(gate1044inter6));
  inv1  gate1277(.a(N3247), .O(gate1044inter7));
  inv1  gate1278(.a(N3484), .O(gate1044inter8));
  nand2 gate1279(.a(gate1044inter8), .b(gate1044inter7), .O(gate1044inter9));
  nand2 gate1280(.a(s_1), .b(gate1044inter3), .O(gate1044inter10));
  nor2  gate1281(.a(gate1044inter10), .b(gate1044inter9), .O(gate1044inter11));
  nor2  gate1282(.a(gate1044inter11), .b(gate1044inter6), .O(gate1044inter12));
  nand2 gate1283(.a(gate1044inter12), .b(gate1044inter1), .O(N3553));
nand2 gate1045( .a(N3250), .b(N3486), .O(N3554) );

  xor2  gate1942(.a(N3488), .b(N3253), .O(gate1046inter0));
  nand2 gate1943(.a(gate1046inter0), .b(s_96), .O(gate1046inter1));
  and2  gate1944(.a(N3488), .b(N3253), .O(gate1046inter2));
  inv1  gate1945(.a(s_96), .O(gate1046inter3));
  inv1  gate1946(.a(s_97), .O(gate1046inter4));
  nand2 gate1947(.a(gate1046inter4), .b(gate1046inter3), .O(gate1046inter5));
  nor2  gate1948(.a(gate1046inter5), .b(gate1046inter2), .O(gate1046inter6));
  inv1  gate1949(.a(N3253), .O(gate1046inter7));
  inv1  gate1950(.a(N3488), .O(gate1046inter8));
  nand2 gate1951(.a(gate1046inter8), .b(gate1046inter7), .O(gate1046inter9));
  nand2 gate1952(.a(s_97), .b(gate1046inter3), .O(gate1046inter10));
  nor2  gate1953(.a(gate1046inter10), .b(gate1046inter9), .O(gate1046inter11));
  nor2  gate1954(.a(gate1046inter11), .b(gate1046inter6), .O(gate1046inter12));
  nand2 gate1955(.a(gate1046inter12), .b(gate1046inter1), .O(N3555));
nand2 gate1047( .a(N3256), .b(N3490), .O(N3556) );

  xor2  gate2180(.a(N3492), .b(N3259), .O(gate1048inter0));
  nand2 gate2181(.a(gate1048inter0), .b(s_130), .O(gate1048inter1));
  and2  gate2182(.a(N3492), .b(N3259), .O(gate1048inter2));
  inv1  gate2183(.a(s_130), .O(gate1048inter3));
  inv1  gate2184(.a(s_131), .O(gate1048inter4));
  nand2 gate2185(.a(gate1048inter4), .b(gate1048inter3), .O(gate1048inter5));
  nor2  gate2186(.a(gate1048inter5), .b(gate1048inter2), .O(gate1048inter6));
  inv1  gate2187(.a(N3259), .O(gate1048inter7));
  inv1  gate2188(.a(N3492), .O(gate1048inter8));
  nand2 gate2189(.a(gate1048inter8), .b(gate1048inter7), .O(gate1048inter9));
  nand2 gate2190(.a(s_131), .b(gate1048inter3), .O(gate1048inter10));
  nor2  gate2191(.a(gate1048inter10), .b(gate1048inter9), .O(gate1048inter11));
  nor2  gate2192(.a(gate1048inter11), .b(gate1048inter6), .O(gate1048inter12));
  nand2 gate2193(.a(gate1048inter12), .b(gate1048inter1), .O(N3557));
and2 gate1049( .a(N3453), .b(N3091), .O(N3558) );
and2 gate1050( .a(N3450), .b(N3088), .O(N3559) );

  xor2  gate2726(.a(N3501), .b(N3262), .O(gate1051inter0));
  nand2 gate2727(.a(gate1051inter0), .b(s_208), .O(gate1051inter1));
  and2  gate2728(.a(N3501), .b(N3262), .O(gate1051inter2));
  inv1  gate2729(.a(s_208), .O(gate1051inter3));
  inv1  gate2730(.a(s_209), .O(gate1051inter4));
  nand2 gate2731(.a(gate1051inter4), .b(gate1051inter3), .O(gate1051inter5));
  nor2  gate2732(.a(gate1051inter5), .b(gate1051inter2), .O(gate1051inter6));
  inv1  gate2733(.a(N3262), .O(gate1051inter7));
  inv1  gate2734(.a(N3501), .O(gate1051inter8));
  nand2 gate2735(.a(gate1051inter8), .b(gate1051inter7), .O(gate1051inter9));
  nand2 gate2736(.a(s_209), .b(gate1051inter3), .O(gate1051inter10));
  nor2  gate2737(.a(gate1051inter10), .b(gate1051inter9), .O(gate1051inter11));
  nor2  gate2738(.a(gate1051inter11), .b(gate1051inter6), .O(gate1051inter12));
  nand2 gate2739(.a(gate1051inter12), .b(gate1051inter1), .O(N3563));
nand2 gate1052( .a(N3265), .b(N3503), .O(N3564) );
nand2 gate1053( .a(N3268), .b(N3505), .O(N3565) );
nand2 gate1054( .a(N3271), .b(N3507), .O(N3566) );

  xor2  gate2110(.a(N3509), .b(N3274), .O(gate1055inter0));
  nand2 gate2111(.a(gate1055inter0), .b(s_120), .O(gate1055inter1));
  and2  gate2112(.a(N3509), .b(N3274), .O(gate1055inter2));
  inv1  gate2113(.a(s_120), .O(gate1055inter3));
  inv1  gate2114(.a(s_121), .O(gate1055inter4));
  nand2 gate2115(.a(gate1055inter4), .b(gate1055inter3), .O(gate1055inter5));
  nor2  gate2116(.a(gate1055inter5), .b(gate1055inter2), .O(gate1055inter6));
  inv1  gate2117(.a(N3274), .O(gate1055inter7));
  inv1  gate2118(.a(N3509), .O(gate1055inter8));
  nand2 gate2119(.a(gate1055inter8), .b(gate1055inter7), .O(gate1055inter9));
  nand2 gate2120(.a(s_121), .b(gate1055inter3), .O(gate1055inter10));
  nor2  gate2121(.a(gate1055inter10), .b(gate1055inter9), .O(gate1055inter11));
  nor2  gate2122(.a(gate1055inter11), .b(gate1055inter6), .O(gate1055inter12));
  nand2 gate2123(.a(gate1055inter12), .b(gate1055inter1), .O(N3567));
nand2 gate1056( .a(N3277), .b(N3511), .O(N3568) );
and2 gate1057( .a(N3459), .b(N3113), .O(N3569) );
and2 gate1058( .a(N3456), .b(N3110), .O(N3570) );
buf1 gate1059( .a(N3453), .O(N3576) );
buf1 gate1060( .a(N3450), .O(N3579) );
buf1 gate1061( .a(N3459), .O(N3585) );
buf1 gate1062( .a(N3456), .O(N3588) );
inv1 gate1063( .a(N3522), .O(N3592) );

  xor2  gate1690(.a(N3405), .b(N3522), .O(gate1064inter0));
  nand2 gate1691(.a(gate1064inter0), .b(s_60), .O(gate1064inter1));
  and2  gate1692(.a(N3405), .b(N3522), .O(gate1064inter2));
  inv1  gate1693(.a(s_60), .O(gate1064inter3));
  inv1  gate1694(.a(s_61), .O(gate1064inter4));
  nand2 gate1695(.a(gate1064inter4), .b(gate1064inter3), .O(gate1064inter5));
  nor2  gate1696(.a(gate1064inter5), .b(gate1064inter2), .O(gate1064inter6));
  inv1  gate1697(.a(N3522), .O(gate1064inter7));
  inv1  gate1698(.a(N3405), .O(gate1064inter8));
  nand2 gate1699(.a(gate1064inter8), .b(gate1064inter7), .O(gate1064inter9));
  nand2 gate1700(.a(s_61), .b(gate1064inter3), .O(gate1064inter10));
  nor2  gate1701(.a(gate1064inter10), .b(gate1064inter9), .O(gate1064inter11));
  nor2  gate1702(.a(gate1064inter11), .b(gate1064inter6), .O(gate1064inter12));
  nand2 gate1703(.a(gate1064inter12), .b(gate1064inter1), .O(N3593));
inv1 gate1065( .a(N3525), .O(N3594) );

  xor2  gate1704(.a(N3406), .b(N3525), .O(gate1066inter0));
  nand2 gate1705(.a(gate1066inter0), .b(s_62), .O(gate1066inter1));
  and2  gate1706(.a(N3406), .b(N3525), .O(gate1066inter2));
  inv1  gate1707(.a(s_62), .O(gate1066inter3));
  inv1  gate1708(.a(s_63), .O(gate1066inter4));
  nand2 gate1709(.a(gate1066inter4), .b(gate1066inter3), .O(gate1066inter5));
  nor2  gate1710(.a(gate1066inter5), .b(gate1066inter2), .O(gate1066inter6));
  inv1  gate1711(.a(N3525), .O(gate1066inter7));
  inv1  gate1712(.a(N3406), .O(gate1066inter8));
  nand2 gate1713(.a(gate1066inter8), .b(gate1066inter7), .O(gate1066inter9));
  nand2 gate1714(.a(s_63), .b(gate1066inter3), .O(gate1066inter10));
  nor2  gate1715(.a(gate1066inter10), .b(gate1066inter9), .O(gate1066inter11));
  nor2  gate1716(.a(gate1066inter11), .b(gate1066inter6), .O(gate1066inter12));
  nand2 gate1717(.a(gate1066inter12), .b(gate1066inter1), .O(N3595));
inv1 gate1067( .a(N3528), .O(N3596) );
nand2 gate1068( .a(N3528), .b(N2630), .O(N3597) );
nand2 gate1069( .a(N3531), .b(N2376), .O(N3598) );
inv1 gate1070( .a(N3531), .O(N3599) );
and2 gate1071( .a(N3551), .b(N800), .O(N3600) );

  xor2  gate2264(.a(N3483), .b(N3552), .O(gate1072inter0));
  nand2 gate2265(.a(gate1072inter0), .b(s_142), .O(gate1072inter1));
  and2  gate2266(.a(N3483), .b(N3552), .O(gate1072inter2));
  inv1  gate2267(.a(s_142), .O(gate1072inter3));
  inv1  gate2268(.a(s_143), .O(gate1072inter4));
  nand2 gate2269(.a(gate1072inter4), .b(gate1072inter3), .O(gate1072inter5));
  nor2  gate2270(.a(gate1072inter5), .b(gate1072inter2), .O(gate1072inter6));
  inv1  gate2271(.a(N3552), .O(gate1072inter7));
  inv1  gate2272(.a(N3483), .O(gate1072inter8));
  nand2 gate2273(.a(gate1072inter8), .b(gate1072inter7), .O(gate1072inter9));
  nand2 gate2274(.a(s_143), .b(gate1072inter3), .O(gate1072inter10));
  nor2  gate2275(.a(gate1072inter10), .b(gate1072inter9), .O(gate1072inter11));
  nor2  gate2276(.a(gate1072inter11), .b(gate1072inter6), .O(gate1072inter12));
  nand2 gate2277(.a(gate1072inter12), .b(gate1072inter1), .O(N3603));

  xor2  gate1788(.a(N3485), .b(N3553), .O(gate1073inter0));
  nand2 gate1789(.a(gate1073inter0), .b(s_74), .O(gate1073inter1));
  and2  gate1790(.a(N3485), .b(N3553), .O(gate1073inter2));
  inv1  gate1791(.a(s_74), .O(gate1073inter3));
  inv1  gate1792(.a(s_75), .O(gate1073inter4));
  nand2 gate1793(.a(gate1073inter4), .b(gate1073inter3), .O(gate1073inter5));
  nor2  gate1794(.a(gate1073inter5), .b(gate1073inter2), .O(gate1073inter6));
  inv1  gate1795(.a(N3553), .O(gate1073inter7));
  inv1  gate1796(.a(N3485), .O(gate1073inter8));
  nand2 gate1797(.a(gate1073inter8), .b(gate1073inter7), .O(gate1073inter9));
  nand2 gate1798(.a(s_75), .b(gate1073inter3), .O(gate1073inter10));
  nor2  gate1799(.a(gate1073inter10), .b(gate1073inter9), .O(gate1073inter11));
  nor2  gate1800(.a(gate1073inter11), .b(gate1073inter6), .O(gate1073inter12));
  nand2 gate1801(.a(gate1073inter12), .b(gate1073inter1), .O(N3608));
nand2 gate1074( .a(N3554), .b(N3487), .O(N3612) );
nand2 gate1075( .a(N3555), .b(N3489), .O(N3615) );
nand2 gate1076( .a(N3556), .b(N3491), .O(N3616) );

  xor2  gate2026(.a(N3493), .b(N3557), .O(gate1077inter0));
  nand2 gate2027(.a(gate1077inter0), .b(s_108), .O(gate1077inter1));
  and2  gate2028(.a(N3493), .b(N3557), .O(gate1077inter2));
  inv1  gate2029(.a(s_108), .O(gate1077inter3));
  inv1  gate2030(.a(s_109), .O(gate1077inter4));
  nand2 gate2031(.a(gate1077inter4), .b(gate1077inter3), .O(gate1077inter5));
  nor2  gate2032(.a(gate1077inter5), .b(gate1077inter2), .O(gate1077inter6));
  inv1  gate2033(.a(N3557), .O(gate1077inter7));
  inv1  gate2034(.a(N3493), .O(gate1077inter8));
  nand2 gate2035(.a(gate1077inter8), .b(gate1077inter7), .O(gate1077inter9));
  nand2 gate2036(.a(s_109), .b(gate1077inter3), .O(gate1077inter10));
  nor2  gate2037(.a(gate1077inter10), .b(gate1077inter9), .O(gate1077inter11));
  nor2  gate2038(.a(gate1077inter11), .b(gate1077inter6), .O(gate1077inter12));
  nand2 gate2039(.a(gate1077inter12), .b(gate1077inter1), .O(N3622));
inv1 gate1078( .a(N3534), .O(N3629) );
nand2 gate1079( .a(N3534), .b(N2645), .O(N3630) );
inv1 gate1080( .a(N3537), .O(N3631) );
nand2 gate1081( .a(N3537), .b(N2655), .O(N3632) );

  xor2  gate1452(.a(N2403), .b(N3540), .O(gate1082inter0));
  nand2 gate1453(.a(gate1082inter0), .b(s_26), .O(gate1082inter1));
  and2  gate1454(.a(N2403), .b(N3540), .O(gate1082inter2));
  inv1  gate1455(.a(s_26), .O(gate1082inter3));
  inv1  gate1456(.a(s_27), .O(gate1082inter4));
  nand2 gate1457(.a(gate1082inter4), .b(gate1082inter3), .O(gate1082inter5));
  nor2  gate1458(.a(gate1082inter5), .b(gate1082inter2), .O(gate1082inter6));
  inv1  gate1459(.a(N3540), .O(gate1082inter7));
  inv1  gate1460(.a(N2403), .O(gate1082inter8));
  nand2 gate1461(.a(gate1082inter8), .b(gate1082inter7), .O(gate1082inter9));
  nand2 gate1462(.a(s_27), .b(gate1082inter3), .O(gate1082inter10));
  nor2  gate1463(.a(gate1082inter10), .b(gate1082inter9), .O(gate1082inter11));
  nor2  gate1464(.a(gate1082inter11), .b(gate1082inter6), .O(gate1082inter12));
  nand2 gate1465(.a(gate1082inter12), .b(gate1082inter1), .O(N3633));
inv1 gate1083( .a(N3540), .O(N3634) );
nand2 gate1084( .a(N3563), .b(N3502), .O(N3635) );

  xor2  gate2446(.a(N3504), .b(N3564), .O(gate1085inter0));
  nand2 gate2447(.a(gate1085inter0), .b(s_168), .O(gate1085inter1));
  and2  gate2448(.a(N3504), .b(N3564), .O(gate1085inter2));
  inv1  gate2449(.a(s_168), .O(gate1085inter3));
  inv1  gate2450(.a(s_169), .O(gate1085inter4));
  nand2 gate2451(.a(gate1085inter4), .b(gate1085inter3), .O(gate1085inter5));
  nor2  gate2452(.a(gate1085inter5), .b(gate1085inter2), .O(gate1085inter6));
  inv1  gate2453(.a(N3564), .O(gate1085inter7));
  inv1  gate2454(.a(N3504), .O(gate1085inter8));
  nand2 gate2455(.a(gate1085inter8), .b(gate1085inter7), .O(gate1085inter9));
  nand2 gate2456(.a(s_169), .b(gate1085inter3), .O(gate1085inter10));
  nor2  gate2457(.a(gate1085inter10), .b(gate1085inter9), .O(gate1085inter11));
  nor2  gate2458(.a(gate1085inter11), .b(gate1085inter6), .O(gate1085inter12));
  nand2 gate2459(.a(gate1085inter12), .b(gate1085inter1), .O(N3640));
nand2 gate1086( .a(N3565), .b(N3506), .O(N3644) );

  xor2  gate2684(.a(N3508), .b(N3566), .O(gate1087inter0));
  nand2 gate2685(.a(gate1087inter0), .b(s_202), .O(gate1087inter1));
  and2  gate2686(.a(N3508), .b(N3566), .O(gate1087inter2));
  inv1  gate2687(.a(s_202), .O(gate1087inter3));
  inv1  gate2688(.a(s_203), .O(gate1087inter4));
  nand2 gate2689(.a(gate1087inter4), .b(gate1087inter3), .O(gate1087inter5));
  nor2  gate2690(.a(gate1087inter5), .b(gate1087inter2), .O(gate1087inter6));
  inv1  gate2691(.a(N3566), .O(gate1087inter7));
  inv1  gate2692(.a(N3508), .O(gate1087inter8));
  nand2 gate2693(.a(gate1087inter8), .b(gate1087inter7), .O(gate1087inter9));
  nand2 gate2694(.a(s_203), .b(gate1087inter3), .O(gate1087inter10));
  nor2  gate2695(.a(gate1087inter10), .b(gate1087inter9), .O(gate1087inter11));
  nor2  gate2696(.a(gate1087inter11), .b(gate1087inter6), .O(gate1087inter12));
  nand2 gate2697(.a(gate1087inter12), .b(gate1087inter1), .O(N3647));
nand2 gate1088( .a(N3567), .b(N3510), .O(N3648) );
nand2 gate1089( .a(N3568), .b(N3512), .O(N3654) );
inv1 gate1090( .a(N3543), .O(N3661) );
nand2 gate1091( .a(N3543), .b(N2656), .O(N3662) );

  xor2  gate2404(.a(N3592), .b(N3238), .O(gate1092inter0));
  nand2 gate2405(.a(gate1092inter0), .b(s_162), .O(gate1092inter1));
  and2  gate2406(.a(N3592), .b(N3238), .O(gate1092inter2));
  inv1  gate2407(.a(s_162), .O(gate1092inter3));
  inv1  gate2408(.a(s_163), .O(gate1092inter4));
  nand2 gate2409(.a(gate1092inter4), .b(gate1092inter3), .O(gate1092inter5));
  nor2  gate2410(.a(gate1092inter5), .b(gate1092inter2), .O(gate1092inter6));
  inv1  gate2411(.a(N3238), .O(gate1092inter7));
  inv1  gate2412(.a(N3592), .O(gate1092inter8));
  nand2 gate2413(.a(gate1092inter8), .b(gate1092inter7), .O(gate1092inter9));
  nand2 gate2414(.a(s_163), .b(gate1092inter3), .O(gate1092inter10));
  nor2  gate2415(.a(gate1092inter10), .b(gate1092inter9), .O(gate1092inter11));
  nor2  gate2416(.a(gate1092inter11), .b(gate1092inter6), .O(gate1092inter12));
  nand2 gate2417(.a(gate1092inter12), .b(gate1092inter1), .O(N3667));

  xor2  gate1382(.a(N3594), .b(N3241), .O(gate1093inter0));
  nand2 gate1383(.a(gate1093inter0), .b(s_16), .O(gate1093inter1));
  and2  gate1384(.a(N3594), .b(N3241), .O(gate1093inter2));
  inv1  gate1385(.a(s_16), .O(gate1093inter3));
  inv1  gate1386(.a(s_17), .O(gate1093inter4));
  nand2 gate1387(.a(gate1093inter4), .b(gate1093inter3), .O(gate1093inter5));
  nor2  gate1388(.a(gate1093inter5), .b(gate1093inter2), .O(gate1093inter6));
  inv1  gate1389(.a(N3241), .O(gate1093inter7));
  inv1  gate1390(.a(N3594), .O(gate1093inter8));
  nand2 gate1391(.a(gate1093inter8), .b(gate1093inter7), .O(gate1093inter9));
  nand2 gate1392(.a(s_17), .b(gate1093inter3), .O(gate1093inter10));
  nor2  gate1393(.a(gate1093inter10), .b(gate1093inter9), .O(gate1093inter11));
  nor2  gate1394(.a(gate1093inter11), .b(gate1093inter6), .O(gate1093inter12));
  nand2 gate1395(.a(gate1093inter12), .b(gate1093inter1), .O(N3668));

  xor2  gate1606(.a(N3596), .b(N2472), .O(gate1094inter0));
  nand2 gate1607(.a(gate1094inter0), .b(s_48), .O(gate1094inter1));
  and2  gate1608(.a(N3596), .b(N2472), .O(gate1094inter2));
  inv1  gate1609(.a(s_48), .O(gate1094inter3));
  inv1  gate1610(.a(s_49), .O(gate1094inter4));
  nand2 gate1611(.a(gate1094inter4), .b(gate1094inter3), .O(gate1094inter5));
  nor2  gate1612(.a(gate1094inter5), .b(gate1094inter2), .O(gate1094inter6));
  inv1  gate1613(.a(N2472), .O(gate1094inter7));
  inv1  gate1614(.a(N3596), .O(gate1094inter8));
  nand2 gate1615(.a(gate1094inter8), .b(gate1094inter7), .O(gate1094inter9));
  nand2 gate1616(.a(s_49), .b(gate1094inter3), .O(gate1094inter10));
  nor2  gate1617(.a(gate1094inter10), .b(gate1094inter9), .O(gate1094inter11));
  nor2  gate1618(.a(gate1094inter11), .b(gate1094inter6), .O(gate1094inter12));
  nand2 gate1619(.a(gate1094inter12), .b(gate1094inter1), .O(N3669));
nand2 gate1095( .a(N2213), .b(N3599), .O(N3670) );
buf1 gate1096( .a(N3600), .O(N3671) );
inv1 gate1097( .a(N3576), .O(N3691) );

  xor2  gate2054(.a(N3494), .b(N3576), .O(gate1098inter0));
  nand2 gate2055(.a(gate1098inter0), .b(s_112), .O(gate1098inter1));
  and2  gate2056(.a(N3494), .b(N3576), .O(gate1098inter2));
  inv1  gate2057(.a(s_112), .O(gate1098inter3));
  inv1  gate2058(.a(s_113), .O(gate1098inter4));
  nand2 gate2059(.a(gate1098inter4), .b(gate1098inter3), .O(gate1098inter5));
  nor2  gate2060(.a(gate1098inter5), .b(gate1098inter2), .O(gate1098inter6));
  inv1  gate2061(.a(N3576), .O(gate1098inter7));
  inv1  gate2062(.a(N3494), .O(gate1098inter8));
  nand2 gate2063(.a(gate1098inter8), .b(gate1098inter7), .O(gate1098inter9));
  nand2 gate2064(.a(s_113), .b(gate1098inter3), .O(gate1098inter10));
  nor2  gate2065(.a(gate1098inter10), .b(gate1098inter9), .O(gate1098inter11));
  nor2  gate2066(.a(gate1098inter11), .b(gate1098inter6), .O(gate1098inter12));
  nand2 gate2067(.a(gate1098inter12), .b(gate1098inter1), .O(N3692));
inv1 gate1099( .a(N3579), .O(N3693) );

  xor2  gate2768(.a(N3496), .b(N3579), .O(gate1100inter0));
  nand2 gate2769(.a(gate1100inter0), .b(s_214), .O(gate1100inter1));
  and2  gate2770(.a(N3496), .b(N3579), .O(gate1100inter2));
  inv1  gate2771(.a(s_214), .O(gate1100inter3));
  inv1  gate2772(.a(s_215), .O(gate1100inter4));
  nand2 gate2773(.a(gate1100inter4), .b(gate1100inter3), .O(gate1100inter5));
  nor2  gate2774(.a(gate1100inter5), .b(gate1100inter2), .O(gate1100inter6));
  inv1  gate2775(.a(N3579), .O(gate1100inter7));
  inv1  gate2776(.a(N3496), .O(gate1100inter8));
  nand2 gate2777(.a(gate1100inter8), .b(gate1100inter7), .O(gate1100inter9));
  nand2 gate2778(.a(s_215), .b(gate1100inter3), .O(gate1100inter10));
  nor2  gate2779(.a(gate1100inter10), .b(gate1100inter9), .O(gate1100inter11));
  nor2  gate2780(.a(gate1100inter11), .b(gate1100inter6), .O(gate1100inter12));
  nand2 gate2781(.a(gate1100inter12), .b(gate1100inter1), .O(N3694));

  xor2  gate1760(.a(N3629), .b(N2475), .O(gate1101inter0));
  nand2 gate1761(.a(gate1101inter0), .b(s_70), .O(gate1101inter1));
  and2  gate1762(.a(N3629), .b(N2475), .O(gate1101inter2));
  inv1  gate1763(.a(s_70), .O(gate1101inter3));
  inv1  gate1764(.a(s_71), .O(gate1101inter4));
  nand2 gate1765(.a(gate1101inter4), .b(gate1101inter3), .O(gate1101inter5));
  nor2  gate1766(.a(gate1101inter5), .b(gate1101inter2), .O(gate1101inter6));
  inv1  gate1767(.a(N2475), .O(gate1101inter7));
  inv1  gate1768(.a(N3629), .O(gate1101inter8));
  nand2 gate1769(.a(gate1101inter8), .b(gate1101inter7), .O(gate1101inter9));
  nand2 gate1770(.a(s_71), .b(gate1101inter3), .O(gate1101inter10));
  nor2  gate1771(.a(gate1101inter10), .b(gate1101inter9), .O(gate1101inter11));
  nor2  gate1772(.a(gate1101inter11), .b(gate1101inter6), .O(gate1101inter12));
  nand2 gate1773(.a(gate1101inter12), .b(gate1101inter1), .O(N3695));
nand2 gate1102( .a(N2478), .b(N3631), .O(N3696) );
nand2 gate1103( .a(N2216), .b(N3634), .O(N3697) );
inv1 gate1104( .a(N3585), .O(N3716) );

  xor2  gate2376(.a(N3513), .b(N3585), .O(gate1105inter0));
  nand2 gate2377(.a(gate1105inter0), .b(s_158), .O(gate1105inter1));
  and2  gate2378(.a(N3513), .b(N3585), .O(gate1105inter2));
  inv1  gate2379(.a(s_158), .O(gate1105inter3));
  inv1  gate2380(.a(s_159), .O(gate1105inter4));
  nand2 gate2381(.a(gate1105inter4), .b(gate1105inter3), .O(gate1105inter5));
  nor2  gate2382(.a(gate1105inter5), .b(gate1105inter2), .O(gate1105inter6));
  inv1  gate2383(.a(N3585), .O(gate1105inter7));
  inv1  gate2384(.a(N3513), .O(gate1105inter8));
  nand2 gate2385(.a(gate1105inter8), .b(gate1105inter7), .O(gate1105inter9));
  nand2 gate2386(.a(s_159), .b(gate1105inter3), .O(gate1105inter10));
  nor2  gate2387(.a(gate1105inter10), .b(gate1105inter9), .O(gate1105inter11));
  nor2  gate2388(.a(gate1105inter11), .b(gate1105inter6), .O(gate1105inter12));
  nand2 gate2389(.a(gate1105inter12), .b(gate1105inter1), .O(N3717));
inv1 gate1106( .a(N3588), .O(N3718) );

  xor2  gate2936(.a(N3515), .b(N3588), .O(gate1107inter0));
  nand2 gate2937(.a(gate1107inter0), .b(s_238), .O(gate1107inter1));
  and2  gate2938(.a(N3515), .b(N3588), .O(gate1107inter2));
  inv1  gate2939(.a(s_238), .O(gate1107inter3));
  inv1  gate2940(.a(s_239), .O(gate1107inter4));
  nand2 gate2941(.a(gate1107inter4), .b(gate1107inter3), .O(gate1107inter5));
  nor2  gate2942(.a(gate1107inter5), .b(gate1107inter2), .O(gate1107inter6));
  inv1  gate2943(.a(N3588), .O(gate1107inter7));
  inv1  gate2944(.a(N3515), .O(gate1107inter8));
  nand2 gate2945(.a(gate1107inter8), .b(gate1107inter7), .O(gate1107inter9));
  nand2 gate2946(.a(s_239), .b(gate1107inter3), .O(gate1107inter10));
  nor2  gate2947(.a(gate1107inter10), .b(gate1107inter9), .O(gate1107inter11));
  nor2  gate2948(.a(gate1107inter11), .b(gate1107inter6), .O(gate1107inter12));
  nand2 gate2949(.a(gate1107inter12), .b(gate1107inter1), .O(N3719));

  xor2  gate1494(.a(N3661), .b(N2481), .O(gate1108inter0));
  nand2 gate1495(.a(gate1108inter0), .b(s_32), .O(gate1108inter1));
  and2  gate1496(.a(N3661), .b(N2481), .O(gate1108inter2));
  inv1  gate1497(.a(s_32), .O(gate1108inter3));
  inv1  gate1498(.a(s_33), .O(gate1108inter4));
  nand2 gate1499(.a(gate1108inter4), .b(gate1108inter3), .O(gate1108inter5));
  nor2  gate1500(.a(gate1108inter5), .b(gate1108inter2), .O(gate1108inter6));
  inv1  gate1501(.a(N2481), .O(gate1108inter7));
  inv1  gate1502(.a(N3661), .O(gate1108inter8));
  nand2 gate1503(.a(gate1108inter8), .b(gate1108inter7), .O(gate1108inter9));
  nand2 gate1504(.a(s_33), .b(gate1108inter3), .O(gate1108inter10));
  nor2  gate1505(.a(gate1108inter10), .b(gate1108inter9), .O(gate1108inter11));
  nor2  gate1506(.a(gate1108inter11), .b(gate1108inter6), .O(gate1108inter12));
  nand2 gate1507(.a(gate1108inter12), .b(gate1108inter1), .O(N3720));
nand2 gate1109( .a(N3667), .b(N3593), .O(N3721) );
nand2 gate1110( .a(N3668), .b(N3595), .O(N3722) );
nand2 gate1111( .a(N3669), .b(N3597), .O(N3723) );
nand2 gate1112( .a(N3670), .b(N3598), .O(N3726) );
inv1 gate1113( .a(N3600), .O(N3727) );
nand2 gate1114( .a(N3364), .b(N3691), .O(N3728) );

  xor2  gate1354(.a(N3693), .b(N3367), .O(gate1115inter0));
  nand2 gate1355(.a(gate1115inter0), .b(s_12), .O(gate1115inter1));
  and2  gate1356(.a(N3693), .b(N3367), .O(gate1115inter2));
  inv1  gate1357(.a(s_12), .O(gate1115inter3));
  inv1  gate1358(.a(s_13), .O(gate1115inter4));
  nand2 gate1359(.a(gate1115inter4), .b(gate1115inter3), .O(gate1115inter5));
  nor2  gate1360(.a(gate1115inter5), .b(gate1115inter2), .O(gate1115inter6));
  inv1  gate1361(.a(N3367), .O(gate1115inter7));
  inv1  gate1362(.a(N3693), .O(gate1115inter8));
  nand2 gate1363(.a(gate1115inter8), .b(gate1115inter7), .O(gate1115inter9));
  nand2 gate1364(.a(s_13), .b(gate1115inter3), .O(gate1115inter10));
  nor2  gate1365(.a(gate1115inter10), .b(gate1115inter9), .O(gate1115inter11));
  nor2  gate1366(.a(gate1115inter11), .b(gate1115inter6), .O(gate1115inter12));
  nand2 gate1367(.a(gate1115inter12), .b(gate1115inter1), .O(N3729));

  xor2  gate2628(.a(N3630), .b(N3695), .O(gate1116inter0));
  nand2 gate2629(.a(gate1116inter0), .b(s_194), .O(gate1116inter1));
  and2  gate2630(.a(N3630), .b(N3695), .O(gate1116inter2));
  inv1  gate2631(.a(s_194), .O(gate1116inter3));
  inv1  gate2632(.a(s_195), .O(gate1116inter4));
  nand2 gate2633(.a(gate1116inter4), .b(gate1116inter3), .O(gate1116inter5));
  nor2  gate2634(.a(gate1116inter5), .b(gate1116inter2), .O(gate1116inter6));
  inv1  gate2635(.a(N3695), .O(gate1116inter7));
  inv1  gate2636(.a(N3630), .O(gate1116inter8));
  nand2 gate2637(.a(gate1116inter8), .b(gate1116inter7), .O(gate1116inter9));
  nand2 gate2638(.a(s_195), .b(gate1116inter3), .O(gate1116inter10));
  nor2  gate2639(.a(gate1116inter10), .b(gate1116inter9), .O(gate1116inter11));
  nor2  gate2640(.a(gate1116inter11), .b(gate1116inter6), .O(gate1116inter12));
  nand2 gate2641(.a(gate1116inter12), .b(gate1116inter1), .O(N3730));
and4 gate1117( .a(N3608), .b(N3615), .c(N3612), .d(N3603), .O(N3731) );
and2 gate1118( .a(N3603), .b(N3293), .O(N3732) );
and3 gate1119( .a(N3608), .b(N3603), .c(N3295), .O(N3733) );
and4 gate1120( .a(N3612), .b(N3603), .c(N3296), .d(N3608), .O(N3734) );
and2 gate1121( .a(N3616), .b(N3301), .O(N3735) );
and3 gate1122( .a(N3622), .b(N3616), .c(N3558), .O(N3736) );

  xor2  gate1676(.a(N3632), .b(N3696), .O(gate1123inter0));
  nand2 gate1677(.a(gate1123inter0), .b(s_58), .O(gate1123inter1));
  and2  gate1678(.a(N3632), .b(N3696), .O(gate1123inter2));
  inv1  gate1679(.a(s_58), .O(gate1123inter3));
  inv1  gate1680(.a(s_59), .O(gate1123inter4));
  nand2 gate1681(.a(gate1123inter4), .b(gate1123inter3), .O(gate1123inter5));
  nor2  gate1682(.a(gate1123inter5), .b(gate1123inter2), .O(gate1123inter6));
  inv1  gate1683(.a(N3696), .O(gate1123inter7));
  inv1  gate1684(.a(N3632), .O(gate1123inter8));
  nand2 gate1685(.a(gate1123inter8), .b(gate1123inter7), .O(gate1123inter9));
  nand2 gate1686(.a(s_59), .b(gate1123inter3), .O(gate1123inter10));
  nor2  gate1687(.a(gate1123inter10), .b(gate1123inter9), .O(gate1123inter11));
  nor2  gate1688(.a(gate1123inter11), .b(gate1123inter6), .O(gate1123inter12));
  nand2 gate1689(.a(gate1123inter12), .b(gate1123inter1), .O(N3737));

  xor2  gate1578(.a(N3633), .b(N3697), .O(gate1124inter0));
  nand2 gate1579(.a(gate1124inter0), .b(s_44), .O(gate1124inter1));
  and2  gate1580(.a(N3633), .b(N3697), .O(gate1124inter2));
  inv1  gate1581(.a(s_44), .O(gate1124inter3));
  inv1  gate1582(.a(s_45), .O(gate1124inter4));
  nand2 gate1583(.a(gate1124inter4), .b(gate1124inter3), .O(gate1124inter5));
  nor2  gate1584(.a(gate1124inter5), .b(gate1124inter2), .O(gate1124inter6));
  inv1  gate1585(.a(N3697), .O(gate1124inter7));
  inv1  gate1586(.a(N3633), .O(gate1124inter8));
  nand2 gate1587(.a(gate1124inter8), .b(gate1124inter7), .O(gate1124inter9));
  nand2 gate1588(.a(s_45), .b(gate1124inter3), .O(gate1124inter10));
  nor2  gate1589(.a(gate1124inter10), .b(gate1124inter9), .O(gate1124inter11));
  nor2  gate1590(.a(gate1124inter11), .b(gate1124inter6), .O(gate1124inter12));
  nand2 gate1591(.a(gate1124inter12), .b(gate1124inter1), .O(N3740));

  xor2  gate1648(.a(N3716), .b(N3394), .O(gate1125inter0));
  nand2 gate1649(.a(gate1125inter0), .b(s_54), .O(gate1125inter1));
  and2  gate1650(.a(N3716), .b(N3394), .O(gate1125inter2));
  inv1  gate1651(.a(s_54), .O(gate1125inter3));
  inv1  gate1652(.a(s_55), .O(gate1125inter4));
  nand2 gate1653(.a(gate1125inter4), .b(gate1125inter3), .O(gate1125inter5));
  nor2  gate1654(.a(gate1125inter5), .b(gate1125inter2), .O(gate1125inter6));
  inv1  gate1655(.a(N3394), .O(gate1125inter7));
  inv1  gate1656(.a(N3716), .O(gate1125inter8));
  nand2 gate1657(.a(gate1125inter8), .b(gate1125inter7), .O(gate1125inter9));
  nand2 gate1658(.a(s_55), .b(gate1125inter3), .O(gate1125inter10));
  nor2  gate1659(.a(gate1125inter10), .b(gate1125inter9), .O(gate1125inter11));
  nor2  gate1660(.a(gate1125inter11), .b(gate1125inter6), .O(gate1125inter12));
  nand2 gate1661(.a(gate1125inter12), .b(gate1125inter1), .O(N3741));
nand2 gate1126( .a(N3397), .b(N3718), .O(N3742) );
nand2 gate1127( .a(N3720), .b(N3662), .O(N3743) );
and4 gate1128( .a(N3640), .b(N3647), .c(N3644), .d(N3635), .O(N3744) );
and2 gate1129( .a(N3635), .b(N3306), .O(N3745) );
and3 gate1130( .a(N3640), .b(N3635), .c(N3308), .O(N3746) );
and4 gate1131( .a(N3644), .b(N3635), .c(N3309), .d(N3640), .O(N3747) );
and2 gate1132( .a(N3648), .b(N3314), .O(N3748) );
and3 gate1133( .a(N3654), .b(N3648), .c(N3569), .O(N3749) );
inv1 gate1134( .a(N3721), .O(N3750) );
and2 gate1135( .a(N3722), .b(N246), .O(N3753) );

  xor2  gate2278(.a(N3692), .b(N3728), .O(gate1136inter0));
  nand2 gate2279(.a(gate1136inter0), .b(s_144), .O(gate1136inter1));
  and2  gate2280(.a(N3692), .b(N3728), .O(gate1136inter2));
  inv1  gate2281(.a(s_144), .O(gate1136inter3));
  inv1  gate2282(.a(s_145), .O(gate1136inter4));
  nand2 gate2283(.a(gate1136inter4), .b(gate1136inter3), .O(gate1136inter5));
  nor2  gate2284(.a(gate1136inter5), .b(gate1136inter2), .O(gate1136inter6));
  inv1  gate2285(.a(N3728), .O(gate1136inter7));
  inv1  gate2286(.a(N3692), .O(gate1136inter8));
  nand2 gate2287(.a(gate1136inter8), .b(gate1136inter7), .O(gate1136inter9));
  nand2 gate2288(.a(s_145), .b(gate1136inter3), .O(gate1136inter10));
  nor2  gate2289(.a(gate1136inter10), .b(gate1136inter9), .O(gate1136inter11));
  nor2  gate2290(.a(gate1136inter11), .b(gate1136inter6), .O(gate1136inter12));
  nand2 gate2291(.a(gate1136inter12), .b(gate1136inter1), .O(N3754));
nand2 gate1137( .a(N3729), .b(N3694), .O(N3758) );
inv1 gate1138( .a(N3731), .O(N3761) );
or4 gate1139( .a(N3291), .b(N3732), .c(N3733), .d(N3734), .O(N3762) );

  xor2  gate2040(.a(N3717), .b(N3741), .O(gate1140inter0));
  nand2 gate2041(.a(gate1140inter0), .b(s_110), .O(gate1140inter1));
  and2  gate2042(.a(N3717), .b(N3741), .O(gate1140inter2));
  inv1  gate2043(.a(s_110), .O(gate1140inter3));
  inv1  gate2044(.a(s_111), .O(gate1140inter4));
  nand2 gate2045(.a(gate1140inter4), .b(gate1140inter3), .O(gate1140inter5));
  nor2  gate2046(.a(gate1140inter5), .b(gate1140inter2), .O(gate1140inter6));
  inv1  gate2047(.a(N3741), .O(gate1140inter7));
  inv1  gate2048(.a(N3717), .O(gate1140inter8));
  nand2 gate2049(.a(gate1140inter8), .b(gate1140inter7), .O(gate1140inter9));
  nand2 gate2050(.a(s_111), .b(gate1140inter3), .O(gate1140inter10));
  nor2  gate2051(.a(gate1140inter10), .b(gate1140inter9), .O(gate1140inter11));
  nor2  gate2052(.a(gate1140inter11), .b(gate1140inter6), .O(gate1140inter12));
  nand2 gate2053(.a(gate1140inter12), .b(gate1140inter1), .O(N3767));
nand2 gate1141( .a(N3742), .b(N3719), .O(N3771) );
inv1 gate1142( .a(N3744), .O(N3774) );
or4 gate1143( .a(N3304), .b(N3745), .c(N3746), .d(N3747), .O(N3775) );
and2 gate1144( .a(N3723), .b(N3480), .O(N3778) );
and3 gate1145( .a(N3726), .b(N3723), .c(N3409), .O(N3779) );
or2 gate1146( .a(N2125), .b(N3753), .O(N3780) );
and2 gate1147( .a(N3750), .b(N800), .O(N3790) );
and2 gate1148( .a(N3737), .b(N3500), .O(N3793) );
and3 gate1149( .a(N3740), .b(N3737), .c(N3428), .O(N3794) );
or3 gate1150( .a(N3479), .b(N3778), .c(N3779), .O(N3802) );
buf1 gate1151( .a(N3780), .O(N3803) );
buf1 gate1152( .a(N3780), .O(N3804) );
inv1 gate1153( .a(N3762), .O(N3805) );
and5 gate1154( .a(N3622), .b(N3730), .c(N3754), .d(N3616), .e(N3758), .O(N3806) );
and4 gate1155( .a(N3754), .b(N3616), .c(N3559), .d(N3622), .O(N3807) );
and5 gate1156( .a(N3758), .b(N3754), .c(N3616), .d(N3498), .e(N3622), .O(N3808) );
buf1 gate1157( .a(N3790), .O(N3809) );
or3 gate1158( .a(N3499), .b(N3793), .c(N3794), .O(N3811) );
inv1 gate1159( .a(N3775), .O(N3812) );
and5 gate1160( .a(N3654), .b(N3743), .c(N3767), .d(N3648), .e(N3771), .O(N3813) );
and4 gate1161( .a(N3767), .b(N3648), .c(N3570), .d(N3654), .O(N3814) );
and5 gate1162( .a(N3771), .b(N3767), .c(N3648), .d(N3517), .e(N3654), .O(N3815) );
or5 gate1163( .a(N3299), .b(N3735), .c(N3736), .d(N3807), .e(N3808), .O(N3816) );
and2 gate1164( .a(N3806), .b(N3802), .O(N3817) );
nand2 gate1165( .a(N3805), .b(N3761), .O(N3818) );
inv1 gate1166( .a(N3790), .O(N3819) );
or5 gate1167( .a(N3312), .b(N3748), .c(N3749), .d(N3814), .e(N3815), .O(N3820) );
and2 gate1168( .a(N3813), .b(N3811), .O(N3821) );
nand2 gate1169( .a(N3812), .b(N3774), .O(N3822) );
or2 gate1170( .a(N3816), .b(N3817), .O(N3823) );
and3 gate1171( .a(N3727), .b(N3819), .c(N2841), .O(N3826) );
or2 gate1172( .a(N3820), .b(N3821), .O(N3827) );
inv1 gate1173( .a(N3823), .O(N3834) );
and2 gate1174( .a(N3818), .b(N3823), .O(N3835) );
inv1 gate1175( .a(N3827), .O(N3836) );
and2 gate1176( .a(N3822), .b(N3827), .O(N3837) );
and2 gate1177( .a(N3762), .b(N3834), .O(N3838) );
and2 gate1178( .a(N3775), .b(N3836), .O(N3839) );
or2 gate1179( .a(N3838), .b(N3835), .O(N3840) );
or2 gate1180( .a(N3839), .b(N3837), .O(N3843) );
buf1 gate1181( .a(N3843), .O(N3851) );

  xor2  gate1886(.a(N3840), .b(N3843), .O(gate1182inter0));
  nand2 gate1887(.a(gate1182inter0), .b(s_88), .O(gate1182inter1));
  and2  gate1888(.a(N3840), .b(N3843), .O(gate1182inter2));
  inv1  gate1889(.a(s_88), .O(gate1182inter3));
  inv1  gate1890(.a(s_89), .O(gate1182inter4));
  nand2 gate1891(.a(gate1182inter4), .b(gate1182inter3), .O(gate1182inter5));
  nor2  gate1892(.a(gate1182inter5), .b(gate1182inter2), .O(gate1182inter6));
  inv1  gate1893(.a(N3843), .O(gate1182inter7));
  inv1  gate1894(.a(N3840), .O(gate1182inter8));
  nand2 gate1895(.a(gate1182inter8), .b(gate1182inter7), .O(gate1182inter9));
  nand2 gate1896(.a(s_89), .b(gate1182inter3), .O(gate1182inter10));
  nor2  gate1897(.a(gate1182inter10), .b(gate1182inter9), .O(gate1182inter11));
  nor2  gate1898(.a(gate1182inter11), .b(gate1182inter6), .O(gate1182inter12));
  nand2 gate1899(.a(gate1182inter12), .b(gate1182inter1), .O(N3852));
and2 gate1183( .a(N3843), .b(N3852), .O(N3857) );
and2 gate1184( .a(N3852), .b(N3840), .O(N3858) );
or2 gate1185( .a(N3857), .b(N3858), .O(N3859) );
inv1 gate1186( .a(N3859), .O(N3864) );
and2 gate1187( .a(N3859), .b(N3864), .O(N3869) );
or2 gate1188( .a(N3869), .b(N3864), .O(N3870) );
inv1 gate1189( .a(N3870), .O(N3875) );
and3 gate1190( .a(N2826), .b(N3028), .c(N3870), .O(N3876) );
and3 gate1191( .a(N3826), .b(N3876), .c(N1591), .O(N3877) );
buf1 gate1192( .a(N3877), .O(N3881) );
inv1 gate1193( .a(N3877), .O(N3882) );
buf1 gate1194( .a(N143_I), .O(N143_O) );
buf1 gate1195( .a(N144_I), .O(N144_O) );
buf1 gate1196( .a(N145_I), .O(N145_O) );
buf1 gate1197( .a(N146_I), .O(N146_O) );
buf1 gate1198( .a(N147_I), .O(N147_O) );
buf1 gate1199( .a(N148_I), .O(N148_O) );
buf1 gate1200( .a(N149_I), .O(N149_O) );
buf1 gate1201( .a(N150_I), .O(N150_O) );
buf1 gate1202( .a(N151_I), .O(N151_O) );
buf1 gate1203( .a(N152_I), .O(N152_O) );
buf1 gate1204( .a(N153_I), .O(N153_O) );
buf1 gate1205( .a(N154_I), .O(N154_O) );
buf1 gate1206( .a(N155_I), .O(N155_O) );
buf1 gate1207( .a(N156_I), .O(N156_O) );
buf1 gate1208( .a(N157_I), .O(N157_O) );
buf1 gate1209( .a(N158_I), .O(N158_O) );
buf1 gate1210( .a(N159_I), .O(N159_O) );
buf1 gate1211( .a(N160_I), .O(N160_O) );
buf1 gate1212( .a(N161_I), .O(N161_O) );
buf1 gate1213( .a(N162_I), .O(N162_O) );
buf1 gate1214( .a(N163_I), .O(N163_O) );
buf1 gate1215( .a(N164_I), .O(N164_O) );
buf1 gate1216( .a(N165_I), .O(N165_O) );
buf1 gate1217( .a(N166_I), .O(N166_O) );
buf1 gate1218( .a(N167_I), .O(N167_O) );
buf1 gate1219( .a(N168_I), .O(N168_O) );
buf1 gate1220( .a(N169_I), .O(N169_O) );
buf1 gate1221( .a(N170_I), .O(N170_O) );
buf1 gate1222( .a(N171_I), .O(N171_O) );
buf1 gate1223( .a(N172_I), .O(N172_O) );
buf1 gate1224( .a(N173_I), .O(N173_O) );
buf1 gate1225( .a(N174_I), .O(N174_O) );
buf1 gate1226( .a(N175_I), .O(N175_O) );
buf1 gate1227( .a(N176_I), .O(N176_O) );
buf1 gate1228( .a(N177_I), .O(N177_O) );
buf1 gate1229( .a(N178_I), .O(N178_O) );
buf1 gate1230( .a(N179_I), .O(N179_O) );
buf1 gate1231( .a(N180_I), .O(N180_O) );
buf1 gate1232( .a(N181_I), .O(N181_O) );
buf1 gate1233( .a(N182_I), .O(N182_O) );
buf1 gate1234( .a(N183_I), .O(N183_O) );
buf1 gate1235( .a(N184_I), .O(N184_O) );
buf1 gate1236( .a(N185_I), .O(N185_O) );
buf1 gate1237( .a(N186_I), .O(N186_O) );
buf1 gate1238( .a(N187_I), .O(N187_O) );
buf1 gate1239( .a(N188_I), .O(N188_O) );
buf1 gate1240( .a(N189_I), .O(N189_O) );
buf1 gate1241( .a(N190_I), .O(N190_O) );
buf1 gate1242( .a(N191_I), .O(N191_O) );
buf1 gate1243( .a(N192_I), .O(N192_O) );
buf1 gate1244( .a(N193_I), .O(N193_O) );
buf1 gate1245( .a(N194_I), .O(N194_O) );
buf1 gate1246( .a(N195_I), .O(N195_O) );
buf1 gate1247( .a(N196_I), .O(N196_O) );
buf1 gate1248( .a(N197_I), .O(N197_O) );
buf1 gate1249( .a(N198_I), .O(N198_O) );
buf1 gate1250( .a(N199_I), .O(N199_O) );
buf1 gate1251( .a(N200_I), .O(N200_O) );
buf1 gate1252( .a(N201_I), .O(N201_O) );
buf1 gate1253( .a(N202_I), .O(N202_O) );
buf1 gate1254( .a(N203_I), .O(N203_O) );
buf1 gate1255( .a(N204_I), .O(N204_O) );
buf1 gate1256( .a(N205_I), .O(N205_O) );
buf1 gate1257( .a(N206_I), .O(N206_O) );
buf1 gate1258( .a(N207_I), .O(N207_O) );
buf1 gate1259( .a(N208_I), .O(N208_O) );
buf1 gate1260( .a(N209_I), .O(N209_O) );
buf1 gate1261( .a(N210_I), .O(N210_O) );
buf1 gate1262( .a(N211_I), .O(N211_O) );
buf1 gate1263( .a(N212_I), .O(N212_O) );
buf1 gate1264( .a(N213_I), .O(N213_O) );
buf1 gate1265( .a(N214_I), .O(N214_O) );
buf1 gate1266( .a(N215_I), .O(N215_O) );
buf1 gate1267( .a(N216_I), .O(N216_O) );
buf1 gate1268( .a(N217_I), .O(N217_O) );
buf1 gate1269( .a(N218_I), .O(N218_O) );

endmodule