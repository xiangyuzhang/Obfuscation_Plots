module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate1387(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate1388(.a(gate13inter0), .b(s_120), .O(gate13inter1));
  and2  gate1389(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate1390(.a(s_120), .O(gate13inter3));
  inv1  gate1391(.a(s_121), .O(gate13inter4));
  nand2 gate1392(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate1393(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate1394(.a(G9), .O(gate13inter7));
  inv1  gate1395(.a(G10), .O(gate13inter8));
  nand2 gate1396(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate1397(.a(s_121), .b(gate13inter3), .O(gate13inter10));
  nor2  gate1398(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate1399(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate1400(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate1093(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate1094(.a(gate18inter0), .b(s_78), .O(gate18inter1));
  and2  gate1095(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate1096(.a(s_78), .O(gate18inter3));
  inv1  gate1097(.a(s_79), .O(gate18inter4));
  nand2 gate1098(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate1099(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate1100(.a(G19), .O(gate18inter7));
  inv1  gate1101(.a(G20), .O(gate18inter8));
  nand2 gate1102(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate1103(.a(s_79), .b(gate18inter3), .O(gate18inter10));
  nor2  gate1104(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate1105(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate1106(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate2241(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate2242(.a(gate27inter0), .b(s_242), .O(gate27inter1));
  and2  gate2243(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate2244(.a(s_242), .O(gate27inter3));
  inv1  gate2245(.a(s_243), .O(gate27inter4));
  nand2 gate2246(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate2247(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate2248(.a(G2), .O(gate27inter7));
  inv1  gate2249(.a(G6), .O(gate27inter8));
  nand2 gate2250(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate2251(.a(s_243), .b(gate27inter3), .O(gate27inter10));
  nor2  gate2252(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate2253(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate2254(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );

  xor2  gate1905(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate1906(.a(gate30inter0), .b(s_194), .O(gate30inter1));
  and2  gate1907(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate1908(.a(s_194), .O(gate30inter3));
  inv1  gate1909(.a(s_195), .O(gate30inter4));
  nand2 gate1910(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate1911(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate1912(.a(G11), .O(gate30inter7));
  inv1  gate1913(.a(G15), .O(gate30inter8));
  nand2 gate1914(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate1915(.a(s_195), .b(gate30inter3), .O(gate30inter10));
  nor2  gate1916(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate1917(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate1918(.a(gate30inter12), .b(gate30inter1), .O(G329));

  xor2  gate575(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate576(.a(gate31inter0), .b(s_4), .O(gate31inter1));
  and2  gate577(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate578(.a(s_4), .O(gate31inter3));
  inv1  gate579(.a(s_5), .O(gate31inter4));
  nand2 gate580(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate581(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate582(.a(G4), .O(gate31inter7));
  inv1  gate583(.a(G8), .O(gate31inter8));
  nand2 gate584(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate585(.a(s_5), .b(gate31inter3), .O(gate31inter10));
  nor2  gate586(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate587(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate588(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate2339(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate2340(.a(gate33inter0), .b(s_256), .O(gate33inter1));
  and2  gate2341(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate2342(.a(s_256), .O(gate33inter3));
  inv1  gate2343(.a(s_257), .O(gate33inter4));
  nand2 gate2344(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate2345(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate2346(.a(G17), .O(gate33inter7));
  inv1  gate2347(.a(G21), .O(gate33inter8));
  nand2 gate2348(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate2349(.a(s_257), .b(gate33inter3), .O(gate33inter10));
  nor2  gate2350(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate2351(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate2352(.a(gate33inter12), .b(gate33inter1), .O(G338));
nand2 gate34( .a(G25), .b(G29), .O(G341) );

  xor2  gate603(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate604(.a(gate35inter0), .b(s_8), .O(gate35inter1));
  and2  gate605(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate606(.a(s_8), .O(gate35inter3));
  inv1  gate607(.a(s_9), .O(gate35inter4));
  nand2 gate608(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate609(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate610(.a(G18), .O(gate35inter7));
  inv1  gate611(.a(G22), .O(gate35inter8));
  nand2 gate612(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate613(.a(s_9), .b(gate35inter3), .O(gate35inter10));
  nor2  gate614(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate615(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate616(.a(gate35inter12), .b(gate35inter1), .O(G344));
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate2283(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate2284(.a(gate39inter0), .b(s_248), .O(gate39inter1));
  and2  gate2285(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate2286(.a(s_248), .O(gate39inter3));
  inv1  gate2287(.a(s_249), .O(gate39inter4));
  nand2 gate2288(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate2289(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate2290(.a(G20), .O(gate39inter7));
  inv1  gate2291(.a(G24), .O(gate39inter8));
  nand2 gate2292(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate2293(.a(s_249), .b(gate39inter3), .O(gate39inter10));
  nor2  gate2294(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate2295(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate2296(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate631(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate632(.a(gate44inter0), .b(s_12), .O(gate44inter1));
  and2  gate633(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate634(.a(s_12), .O(gate44inter3));
  inv1  gate635(.a(s_13), .O(gate44inter4));
  nand2 gate636(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate637(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate638(.a(G4), .O(gate44inter7));
  inv1  gate639(.a(G269), .O(gate44inter8));
  nand2 gate640(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate641(.a(s_13), .b(gate44inter3), .O(gate44inter10));
  nor2  gate642(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate643(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate644(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate995(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate996(.a(gate46inter0), .b(s_64), .O(gate46inter1));
  and2  gate997(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate998(.a(s_64), .O(gate46inter3));
  inv1  gate999(.a(s_65), .O(gate46inter4));
  nand2 gate1000(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate1001(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate1002(.a(G6), .O(gate46inter7));
  inv1  gate1003(.a(G272), .O(gate46inter8));
  nand2 gate1004(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate1005(.a(s_65), .b(gate46inter3), .O(gate46inter10));
  nor2  gate1006(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate1007(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate1008(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate939(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate940(.a(gate58inter0), .b(s_56), .O(gate58inter1));
  and2  gate941(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate942(.a(s_56), .O(gate58inter3));
  inv1  gate943(.a(s_57), .O(gate58inter4));
  nand2 gate944(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate945(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate946(.a(G18), .O(gate58inter7));
  inv1  gate947(.a(G290), .O(gate58inter8));
  nand2 gate948(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate949(.a(s_57), .b(gate58inter3), .O(gate58inter10));
  nor2  gate950(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate951(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate952(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate1765(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate1766(.a(gate60inter0), .b(s_174), .O(gate60inter1));
  and2  gate1767(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate1768(.a(s_174), .O(gate60inter3));
  inv1  gate1769(.a(s_175), .O(gate60inter4));
  nand2 gate1770(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate1771(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate1772(.a(G20), .O(gate60inter7));
  inv1  gate1773(.a(G293), .O(gate60inter8));
  nand2 gate1774(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate1775(.a(s_175), .b(gate60inter3), .O(gate60inter10));
  nor2  gate1776(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate1777(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate1778(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate1821(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate1822(.a(gate63inter0), .b(s_182), .O(gate63inter1));
  and2  gate1823(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate1824(.a(s_182), .O(gate63inter3));
  inv1  gate1825(.a(s_183), .O(gate63inter4));
  nand2 gate1826(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate1827(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate1828(.a(G23), .O(gate63inter7));
  inv1  gate1829(.a(G299), .O(gate63inter8));
  nand2 gate1830(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate1831(.a(s_183), .b(gate63inter3), .O(gate63inter10));
  nor2  gate1832(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate1833(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate1834(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate1919(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate1920(.a(gate65inter0), .b(s_196), .O(gate65inter1));
  and2  gate1921(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate1922(.a(s_196), .O(gate65inter3));
  inv1  gate1923(.a(s_197), .O(gate65inter4));
  nand2 gate1924(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate1925(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate1926(.a(G25), .O(gate65inter7));
  inv1  gate1927(.a(G302), .O(gate65inter8));
  nand2 gate1928(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate1929(.a(s_197), .b(gate65inter3), .O(gate65inter10));
  nor2  gate1930(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate1931(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate1932(.a(gate65inter12), .b(gate65inter1), .O(G386));

  xor2  gate617(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate618(.a(gate66inter0), .b(s_10), .O(gate66inter1));
  and2  gate619(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate620(.a(s_10), .O(gate66inter3));
  inv1  gate621(.a(s_11), .O(gate66inter4));
  nand2 gate622(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate623(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate624(.a(G26), .O(gate66inter7));
  inv1  gate625(.a(G302), .O(gate66inter8));
  nand2 gate626(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate627(.a(s_11), .b(gate66inter3), .O(gate66inter10));
  nor2  gate628(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate629(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate630(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );

  xor2  gate1121(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate1122(.a(gate68inter0), .b(s_82), .O(gate68inter1));
  and2  gate1123(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate1124(.a(s_82), .O(gate68inter3));
  inv1  gate1125(.a(s_83), .O(gate68inter4));
  nand2 gate1126(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate1127(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate1128(.a(G28), .O(gate68inter7));
  inv1  gate1129(.a(G305), .O(gate68inter8));
  nand2 gate1130(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate1131(.a(s_83), .b(gate68inter3), .O(gate68inter10));
  nor2  gate1132(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate1133(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate1134(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate2185(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate2186(.a(gate70inter0), .b(s_234), .O(gate70inter1));
  and2  gate2187(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate2188(.a(s_234), .O(gate70inter3));
  inv1  gate2189(.a(s_235), .O(gate70inter4));
  nand2 gate2190(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate2191(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate2192(.a(G30), .O(gate70inter7));
  inv1  gate2193(.a(G308), .O(gate70inter8));
  nand2 gate2194(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate2195(.a(s_235), .b(gate70inter3), .O(gate70inter10));
  nor2  gate2196(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate2197(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate2198(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );

  xor2  gate1975(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate1976(.a(gate79inter0), .b(s_204), .O(gate79inter1));
  and2  gate1977(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate1978(.a(s_204), .O(gate79inter3));
  inv1  gate1979(.a(s_205), .O(gate79inter4));
  nand2 gate1980(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate1981(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate1982(.a(G10), .O(gate79inter7));
  inv1  gate1983(.a(G323), .O(gate79inter8));
  nand2 gate1984(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate1985(.a(s_205), .b(gate79inter3), .O(gate79inter10));
  nor2  gate1986(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate1987(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate1988(.a(gate79inter12), .b(gate79inter1), .O(G400));

  xor2  gate589(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate590(.a(gate80inter0), .b(s_6), .O(gate80inter1));
  and2  gate591(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate592(.a(s_6), .O(gate80inter3));
  inv1  gate593(.a(s_7), .O(gate80inter4));
  nand2 gate594(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate595(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate596(.a(G14), .O(gate80inter7));
  inv1  gate597(.a(G323), .O(gate80inter8));
  nand2 gate598(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate599(.a(s_7), .b(gate80inter3), .O(gate80inter10));
  nor2  gate600(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate601(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate602(.a(gate80inter12), .b(gate80inter1), .O(G401));

  xor2  gate1149(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate1150(.a(gate81inter0), .b(s_86), .O(gate81inter1));
  and2  gate1151(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate1152(.a(s_86), .O(gate81inter3));
  inv1  gate1153(.a(s_87), .O(gate81inter4));
  nand2 gate1154(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate1155(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate1156(.a(G3), .O(gate81inter7));
  inv1  gate1157(.a(G326), .O(gate81inter8));
  nand2 gate1158(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate1159(.a(s_87), .b(gate81inter3), .O(gate81inter10));
  nor2  gate1160(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate1161(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate1162(.a(gate81inter12), .b(gate81inter1), .O(G402));

  xor2  gate1681(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate1682(.a(gate82inter0), .b(s_162), .O(gate82inter1));
  and2  gate1683(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate1684(.a(s_162), .O(gate82inter3));
  inv1  gate1685(.a(s_163), .O(gate82inter4));
  nand2 gate1686(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate1687(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate1688(.a(G7), .O(gate82inter7));
  inv1  gate1689(.a(G326), .O(gate82inter8));
  nand2 gate1690(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate1691(.a(s_163), .b(gate82inter3), .O(gate82inter10));
  nor2  gate1692(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate1693(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate1694(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate1135(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate1136(.a(gate86inter0), .b(s_84), .O(gate86inter1));
  and2  gate1137(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate1138(.a(s_84), .O(gate86inter3));
  inv1  gate1139(.a(s_85), .O(gate86inter4));
  nand2 gate1140(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate1141(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate1142(.a(G8), .O(gate86inter7));
  inv1  gate1143(.a(G332), .O(gate86inter8));
  nand2 gate1144(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate1145(.a(s_85), .b(gate86inter3), .O(gate86inter10));
  nor2  gate1146(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate1147(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate1148(.a(gate86inter12), .b(gate86inter1), .O(G407));

  xor2  gate1457(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate1458(.a(gate87inter0), .b(s_130), .O(gate87inter1));
  and2  gate1459(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate1460(.a(s_130), .O(gate87inter3));
  inv1  gate1461(.a(s_131), .O(gate87inter4));
  nand2 gate1462(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate1463(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate1464(.a(G12), .O(gate87inter7));
  inv1  gate1465(.a(G335), .O(gate87inter8));
  nand2 gate1466(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate1467(.a(s_131), .b(gate87inter3), .O(gate87inter10));
  nor2  gate1468(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate1469(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate1470(.a(gate87inter12), .b(gate87inter1), .O(G408));

  xor2  gate547(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate548(.a(gate88inter0), .b(s_0), .O(gate88inter1));
  and2  gate549(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate550(.a(s_0), .O(gate88inter3));
  inv1  gate551(.a(s_1), .O(gate88inter4));
  nand2 gate552(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate553(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate554(.a(G16), .O(gate88inter7));
  inv1  gate555(.a(G335), .O(gate88inter8));
  nand2 gate556(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate557(.a(s_1), .b(gate88inter3), .O(gate88inter10));
  nor2  gate558(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate559(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate560(.a(gate88inter12), .b(gate88inter1), .O(G409));

  xor2  gate2437(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate2438(.a(gate89inter0), .b(s_270), .O(gate89inter1));
  and2  gate2439(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate2440(.a(s_270), .O(gate89inter3));
  inv1  gate2441(.a(s_271), .O(gate89inter4));
  nand2 gate2442(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate2443(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate2444(.a(G17), .O(gate89inter7));
  inv1  gate2445(.a(G338), .O(gate89inter8));
  nand2 gate2446(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate2447(.a(s_271), .b(gate89inter3), .O(gate89inter10));
  nor2  gate2448(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate2449(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate2450(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );

  xor2  gate1303(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate1304(.a(gate92inter0), .b(s_108), .O(gate92inter1));
  and2  gate1305(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate1306(.a(s_108), .O(gate92inter3));
  inv1  gate1307(.a(s_109), .O(gate92inter4));
  nand2 gate1308(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate1309(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate1310(.a(G29), .O(gate92inter7));
  inv1  gate1311(.a(G341), .O(gate92inter8));
  nand2 gate1312(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate1313(.a(s_109), .b(gate92inter3), .O(gate92inter10));
  nor2  gate1314(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate1315(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate1316(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate2157(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate2158(.a(gate99inter0), .b(s_230), .O(gate99inter1));
  and2  gate2159(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate2160(.a(s_230), .O(gate99inter3));
  inv1  gate2161(.a(s_231), .O(gate99inter4));
  nand2 gate2162(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate2163(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate2164(.a(G27), .O(gate99inter7));
  inv1  gate2165(.a(G353), .O(gate99inter8));
  nand2 gate2166(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate2167(.a(s_231), .b(gate99inter3), .O(gate99inter10));
  nor2  gate2168(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate2169(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate2170(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );

  xor2  gate1037(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate1038(.a(gate103inter0), .b(s_70), .O(gate103inter1));
  and2  gate1039(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate1040(.a(s_70), .O(gate103inter3));
  inv1  gate1041(.a(s_71), .O(gate103inter4));
  nand2 gate1042(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate1043(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate1044(.a(G28), .O(gate103inter7));
  inv1  gate1045(.a(G359), .O(gate103inter8));
  nand2 gate1046(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate1047(.a(s_71), .b(gate103inter3), .O(gate103inter10));
  nor2  gate1048(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate1049(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate1050(.a(gate103inter12), .b(gate103inter1), .O(G424));

  xor2  gate2409(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate2410(.a(gate104inter0), .b(s_266), .O(gate104inter1));
  and2  gate2411(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate2412(.a(s_266), .O(gate104inter3));
  inv1  gate2413(.a(s_267), .O(gate104inter4));
  nand2 gate2414(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate2415(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate2416(.a(G32), .O(gate104inter7));
  inv1  gate2417(.a(G359), .O(gate104inter8));
  nand2 gate2418(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate2419(.a(s_267), .b(gate104inter3), .O(gate104inter10));
  nor2  gate2420(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate2421(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate2422(.a(gate104inter12), .b(gate104inter1), .O(G425));

  xor2  gate1555(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate1556(.a(gate105inter0), .b(s_144), .O(gate105inter1));
  and2  gate1557(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate1558(.a(s_144), .O(gate105inter3));
  inv1  gate1559(.a(s_145), .O(gate105inter4));
  nand2 gate1560(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate1561(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate1562(.a(G362), .O(gate105inter7));
  inv1  gate1563(.a(G363), .O(gate105inter8));
  nand2 gate1564(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate1565(.a(s_145), .b(gate105inter3), .O(gate105inter10));
  nor2  gate1566(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate1567(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate1568(.a(gate105inter12), .b(gate105inter1), .O(G426));

  xor2  gate1177(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate1178(.a(gate106inter0), .b(s_90), .O(gate106inter1));
  and2  gate1179(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate1180(.a(s_90), .O(gate106inter3));
  inv1  gate1181(.a(s_91), .O(gate106inter4));
  nand2 gate1182(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate1183(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate1184(.a(G364), .O(gate106inter7));
  inv1  gate1185(.a(G365), .O(gate106inter8));
  nand2 gate1186(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate1187(.a(s_91), .b(gate106inter3), .O(gate106inter10));
  nor2  gate1188(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate1189(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate1190(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );

  xor2  gate2087(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate2088(.a(gate111inter0), .b(s_220), .O(gate111inter1));
  and2  gate2089(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate2090(.a(s_220), .O(gate111inter3));
  inv1  gate2091(.a(s_221), .O(gate111inter4));
  nand2 gate2092(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate2093(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate2094(.a(G374), .O(gate111inter7));
  inv1  gate2095(.a(G375), .O(gate111inter8));
  nand2 gate2096(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate2097(.a(s_221), .b(gate111inter3), .O(gate111inter10));
  nor2  gate2098(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate2099(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate2100(.a(gate111inter12), .b(gate111inter1), .O(G444));

  xor2  gate1737(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate1738(.a(gate112inter0), .b(s_170), .O(gate112inter1));
  and2  gate1739(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate1740(.a(s_170), .O(gate112inter3));
  inv1  gate1741(.a(s_171), .O(gate112inter4));
  nand2 gate1742(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate1743(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate1744(.a(G376), .O(gate112inter7));
  inv1  gate1745(.a(G377), .O(gate112inter8));
  nand2 gate1746(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate1747(.a(s_171), .b(gate112inter3), .O(gate112inter10));
  nor2  gate1748(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate1749(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate1750(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate1835(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate1836(.a(gate115inter0), .b(s_184), .O(gate115inter1));
  and2  gate1837(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate1838(.a(s_184), .O(gate115inter3));
  inv1  gate1839(.a(s_185), .O(gate115inter4));
  nand2 gate1840(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate1841(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate1842(.a(G382), .O(gate115inter7));
  inv1  gate1843(.a(G383), .O(gate115inter8));
  nand2 gate1844(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate1845(.a(s_185), .b(gate115inter3), .O(gate115inter10));
  nor2  gate1846(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate1847(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate1848(.a(gate115inter12), .b(gate115inter1), .O(G456));

  xor2  gate1513(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate1514(.a(gate116inter0), .b(s_138), .O(gate116inter1));
  and2  gate1515(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate1516(.a(s_138), .O(gate116inter3));
  inv1  gate1517(.a(s_139), .O(gate116inter4));
  nand2 gate1518(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate1519(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate1520(.a(G384), .O(gate116inter7));
  inv1  gate1521(.a(G385), .O(gate116inter8));
  nand2 gate1522(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate1523(.a(s_139), .b(gate116inter3), .O(gate116inter10));
  nor2  gate1524(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate1525(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate1526(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate1023(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate1024(.a(gate123inter0), .b(s_68), .O(gate123inter1));
  and2  gate1025(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate1026(.a(s_68), .O(gate123inter3));
  inv1  gate1027(.a(s_69), .O(gate123inter4));
  nand2 gate1028(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate1029(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate1030(.a(G398), .O(gate123inter7));
  inv1  gate1031(.a(G399), .O(gate123inter8));
  nand2 gate1032(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate1033(.a(s_69), .b(gate123inter3), .O(gate123inter10));
  nor2  gate1034(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate1035(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate1036(.a(gate123inter12), .b(gate123inter1), .O(G480));

  xor2  gate1569(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate1570(.a(gate124inter0), .b(s_146), .O(gate124inter1));
  and2  gate1571(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate1572(.a(s_146), .O(gate124inter3));
  inv1  gate1573(.a(s_147), .O(gate124inter4));
  nand2 gate1574(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate1575(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate1576(.a(G400), .O(gate124inter7));
  inv1  gate1577(.a(G401), .O(gate124inter8));
  nand2 gate1578(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate1579(.a(s_147), .b(gate124inter3), .O(gate124inter10));
  nor2  gate1580(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate1581(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate1582(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate953(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate954(.a(gate128inter0), .b(s_58), .O(gate128inter1));
  and2  gate955(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate956(.a(s_58), .O(gate128inter3));
  inv1  gate957(.a(s_59), .O(gate128inter4));
  nand2 gate958(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate959(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate960(.a(G408), .O(gate128inter7));
  inv1  gate961(.a(G409), .O(gate128inter8));
  nand2 gate962(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate963(.a(s_59), .b(gate128inter3), .O(gate128inter10));
  nor2  gate964(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate965(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate966(.a(gate128inter12), .b(gate128inter1), .O(G495));
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate1219(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate1220(.a(gate130inter0), .b(s_96), .O(gate130inter1));
  and2  gate1221(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate1222(.a(s_96), .O(gate130inter3));
  inv1  gate1223(.a(s_97), .O(gate130inter4));
  nand2 gate1224(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate1225(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate1226(.a(G412), .O(gate130inter7));
  inv1  gate1227(.a(G413), .O(gate130inter8));
  nand2 gate1228(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate1229(.a(s_97), .b(gate130inter3), .O(gate130inter10));
  nor2  gate1230(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate1231(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate1232(.a(gate130inter12), .b(gate130inter1), .O(G501));

  xor2  gate1695(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate1696(.a(gate131inter0), .b(s_164), .O(gate131inter1));
  and2  gate1697(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate1698(.a(s_164), .O(gate131inter3));
  inv1  gate1699(.a(s_165), .O(gate131inter4));
  nand2 gate1700(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate1701(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate1702(.a(G414), .O(gate131inter7));
  inv1  gate1703(.a(G415), .O(gate131inter8));
  nand2 gate1704(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate1705(.a(s_165), .b(gate131inter3), .O(gate131inter10));
  nor2  gate1706(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate1707(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate1708(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );

  xor2  gate2003(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate2004(.a(gate134inter0), .b(s_208), .O(gate134inter1));
  and2  gate2005(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate2006(.a(s_208), .O(gate134inter3));
  inv1  gate2007(.a(s_209), .O(gate134inter4));
  nand2 gate2008(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate2009(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate2010(.a(G420), .O(gate134inter7));
  inv1  gate2011(.a(G421), .O(gate134inter8));
  nand2 gate2012(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate2013(.a(s_209), .b(gate134inter3), .O(gate134inter10));
  nor2  gate2014(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate2015(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate2016(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate1051(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate1052(.a(gate137inter0), .b(s_72), .O(gate137inter1));
  and2  gate1053(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate1054(.a(s_72), .O(gate137inter3));
  inv1  gate1055(.a(s_73), .O(gate137inter4));
  nand2 gate1056(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate1057(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate1058(.a(G426), .O(gate137inter7));
  inv1  gate1059(.a(G429), .O(gate137inter8));
  nand2 gate1060(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate1061(.a(s_73), .b(gate137inter3), .O(gate137inter10));
  nor2  gate1062(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate1063(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate1064(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate1709(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate1710(.a(gate143inter0), .b(s_166), .O(gate143inter1));
  and2  gate1711(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate1712(.a(s_166), .O(gate143inter3));
  inv1  gate1713(.a(s_167), .O(gate143inter4));
  nand2 gate1714(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate1715(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate1716(.a(G462), .O(gate143inter7));
  inv1  gate1717(.a(G465), .O(gate143inter8));
  nand2 gate1718(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate1719(.a(s_167), .b(gate143inter3), .O(gate143inter10));
  nor2  gate1720(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate1721(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate1722(.a(gate143inter12), .b(gate143inter1), .O(G540));

  xor2  gate743(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate744(.a(gate144inter0), .b(s_28), .O(gate144inter1));
  and2  gate745(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate746(.a(s_28), .O(gate144inter3));
  inv1  gate747(.a(s_29), .O(gate144inter4));
  nand2 gate748(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate749(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate750(.a(G468), .O(gate144inter7));
  inv1  gate751(.a(G471), .O(gate144inter8));
  nand2 gate752(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate753(.a(s_29), .b(gate144inter3), .O(gate144inter10));
  nor2  gate754(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate755(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate756(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate1401(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate1402(.a(gate150inter0), .b(s_122), .O(gate150inter1));
  and2  gate1403(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate1404(.a(s_122), .O(gate150inter3));
  inv1  gate1405(.a(s_123), .O(gate150inter4));
  nand2 gate1406(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate1407(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate1408(.a(G504), .O(gate150inter7));
  inv1  gate1409(.a(G507), .O(gate150inter8));
  nand2 gate1410(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate1411(.a(s_123), .b(gate150inter3), .O(gate150inter10));
  nor2  gate1412(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate1413(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate1414(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate1107(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate1108(.a(gate154inter0), .b(s_80), .O(gate154inter1));
  and2  gate1109(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate1110(.a(s_80), .O(gate154inter3));
  inv1  gate1111(.a(s_81), .O(gate154inter4));
  nand2 gate1112(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate1113(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate1114(.a(G429), .O(gate154inter7));
  inv1  gate1115(.a(G522), .O(gate154inter8));
  nand2 gate1116(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate1117(.a(s_81), .b(gate154inter3), .O(gate154inter10));
  nor2  gate1118(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate1119(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate1120(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate771(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate772(.a(gate156inter0), .b(s_32), .O(gate156inter1));
  and2  gate773(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate774(.a(s_32), .O(gate156inter3));
  inv1  gate775(.a(s_33), .O(gate156inter4));
  nand2 gate776(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate777(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate778(.a(G435), .O(gate156inter7));
  inv1  gate779(.a(G525), .O(gate156inter8));
  nand2 gate780(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate781(.a(s_33), .b(gate156inter3), .O(gate156inter10));
  nor2  gate782(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate783(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate784(.a(gate156inter12), .b(gate156inter1), .O(G573));

  xor2  gate2101(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate2102(.a(gate157inter0), .b(s_222), .O(gate157inter1));
  and2  gate2103(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate2104(.a(s_222), .O(gate157inter3));
  inv1  gate2105(.a(s_223), .O(gate157inter4));
  nand2 gate2106(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate2107(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate2108(.a(G438), .O(gate157inter7));
  inv1  gate2109(.a(G528), .O(gate157inter8));
  nand2 gate2110(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate2111(.a(s_223), .b(gate157inter3), .O(gate157inter10));
  nor2  gate2112(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate2113(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate2114(.a(gate157inter12), .b(gate157inter1), .O(G574));

  xor2  gate841(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate842(.a(gate158inter0), .b(s_42), .O(gate158inter1));
  and2  gate843(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate844(.a(s_42), .O(gate158inter3));
  inv1  gate845(.a(s_43), .O(gate158inter4));
  nand2 gate846(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate847(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate848(.a(G441), .O(gate158inter7));
  inv1  gate849(.a(G528), .O(gate158inter8));
  nand2 gate850(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate851(.a(s_43), .b(gate158inter3), .O(gate158inter10));
  nor2  gate852(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate853(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate854(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate659(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate660(.a(gate173inter0), .b(s_16), .O(gate173inter1));
  and2  gate661(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate662(.a(s_16), .O(gate173inter3));
  inv1  gate663(.a(s_17), .O(gate173inter4));
  nand2 gate664(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate665(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate666(.a(G486), .O(gate173inter7));
  inv1  gate667(.a(G552), .O(gate173inter8));
  nand2 gate668(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate669(.a(s_17), .b(gate173inter3), .O(gate173inter10));
  nor2  gate670(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate671(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate672(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );

  xor2  gate1443(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate1444(.a(gate177inter0), .b(s_128), .O(gate177inter1));
  and2  gate1445(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate1446(.a(s_128), .O(gate177inter3));
  inv1  gate1447(.a(s_129), .O(gate177inter4));
  nand2 gate1448(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate1449(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate1450(.a(G498), .O(gate177inter7));
  inv1  gate1451(.a(G558), .O(gate177inter8));
  nand2 gate1452(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate1453(.a(s_129), .b(gate177inter3), .O(gate177inter10));
  nor2  gate1454(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate1455(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate1456(.a(gate177inter12), .b(gate177inter1), .O(G594));

  xor2  gate2143(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate2144(.a(gate178inter0), .b(s_228), .O(gate178inter1));
  and2  gate2145(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate2146(.a(s_228), .O(gate178inter3));
  inv1  gate2147(.a(s_229), .O(gate178inter4));
  nand2 gate2148(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate2149(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate2150(.a(G501), .O(gate178inter7));
  inv1  gate2151(.a(G558), .O(gate178inter8));
  nand2 gate2152(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate2153(.a(s_229), .b(gate178inter3), .O(gate178inter10));
  nor2  gate2154(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate2155(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate2156(.a(gate178inter12), .b(gate178inter1), .O(G595));
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate2311(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate2312(.a(gate183inter0), .b(s_252), .O(gate183inter1));
  and2  gate2313(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate2314(.a(s_252), .O(gate183inter3));
  inv1  gate2315(.a(s_253), .O(gate183inter4));
  nand2 gate2316(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate2317(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate2318(.a(G516), .O(gate183inter7));
  inv1  gate2319(.a(G567), .O(gate183inter8));
  nand2 gate2320(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate2321(.a(s_253), .b(gate183inter3), .O(gate183inter10));
  nor2  gate2322(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate2323(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate2324(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate2115(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate2116(.a(gate188inter0), .b(s_224), .O(gate188inter1));
  and2  gate2117(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate2118(.a(s_224), .O(gate188inter3));
  inv1  gate2119(.a(s_225), .O(gate188inter4));
  nand2 gate2120(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate2121(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate2122(.a(G576), .O(gate188inter7));
  inv1  gate2123(.a(G577), .O(gate188inter8));
  nand2 gate2124(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate2125(.a(s_225), .b(gate188inter3), .O(gate188inter10));
  nor2  gate2126(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate2127(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate2128(.a(gate188inter12), .b(gate188inter1), .O(G617));

  xor2  gate1877(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate1878(.a(gate189inter0), .b(s_190), .O(gate189inter1));
  and2  gate1879(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate1880(.a(s_190), .O(gate189inter3));
  inv1  gate1881(.a(s_191), .O(gate189inter4));
  nand2 gate1882(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate1883(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate1884(.a(G578), .O(gate189inter7));
  inv1  gate1885(.a(G579), .O(gate189inter8));
  nand2 gate1886(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate1887(.a(s_191), .b(gate189inter3), .O(gate189inter10));
  nor2  gate1888(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate1889(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate1890(.a(gate189inter12), .b(gate189inter1), .O(G622));

  xor2  gate2199(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate2200(.a(gate190inter0), .b(s_236), .O(gate190inter1));
  and2  gate2201(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate2202(.a(s_236), .O(gate190inter3));
  inv1  gate2203(.a(s_237), .O(gate190inter4));
  nand2 gate2204(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate2205(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate2206(.a(G580), .O(gate190inter7));
  inv1  gate2207(.a(G581), .O(gate190inter8));
  nand2 gate2208(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate2209(.a(s_237), .b(gate190inter3), .O(gate190inter10));
  nor2  gate2210(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate2211(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate2212(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate2031(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate2032(.a(gate197inter0), .b(s_212), .O(gate197inter1));
  and2  gate2033(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate2034(.a(s_212), .O(gate197inter3));
  inv1  gate2035(.a(s_213), .O(gate197inter4));
  nand2 gate2036(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate2037(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate2038(.a(G594), .O(gate197inter7));
  inv1  gate2039(.a(G595), .O(gate197inter8));
  nand2 gate2040(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate2041(.a(s_213), .b(gate197inter3), .O(gate197inter10));
  nor2  gate2042(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate2043(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate2044(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate2227(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate2228(.a(gate200inter0), .b(s_240), .O(gate200inter1));
  and2  gate2229(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate2230(.a(s_240), .O(gate200inter3));
  inv1  gate2231(.a(s_241), .O(gate200inter4));
  nand2 gate2232(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate2233(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate2234(.a(G600), .O(gate200inter7));
  inv1  gate2235(.a(G601), .O(gate200inter8));
  nand2 gate2236(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate2237(.a(s_241), .b(gate200inter3), .O(gate200inter10));
  nor2  gate2238(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate2239(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate2240(.a(gate200inter12), .b(gate200inter1), .O(G663));

  xor2  gate855(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate856(.a(gate201inter0), .b(s_44), .O(gate201inter1));
  and2  gate857(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate858(.a(s_44), .O(gate201inter3));
  inv1  gate859(.a(s_45), .O(gate201inter4));
  nand2 gate860(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate861(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate862(.a(G602), .O(gate201inter7));
  inv1  gate863(.a(G607), .O(gate201inter8));
  nand2 gate864(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate865(.a(s_45), .b(gate201inter3), .O(gate201inter10));
  nor2  gate866(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate867(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate868(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate1541(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate1542(.a(gate206inter0), .b(s_142), .O(gate206inter1));
  and2  gate1543(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate1544(.a(s_142), .O(gate206inter3));
  inv1  gate1545(.a(s_143), .O(gate206inter4));
  nand2 gate1546(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate1547(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate1548(.a(G632), .O(gate206inter7));
  inv1  gate1549(.a(G637), .O(gate206inter8));
  nand2 gate1550(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate1551(.a(s_143), .b(gate206inter3), .O(gate206inter10));
  nor2  gate1552(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate1553(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate1554(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate729(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate730(.a(gate213inter0), .b(s_26), .O(gate213inter1));
  and2  gate731(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate732(.a(s_26), .O(gate213inter3));
  inv1  gate733(.a(s_27), .O(gate213inter4));
  nand2 gate734(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate735(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate736(.a(G602), .O(gate213inter7));
  inv1  gate737(.a(G672), .O(gate213inter8));
  nand2 gate738(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate739(.a(s_27), .b(gate213inter3), .O(gate213inter10));
  nor2  gate740(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate741(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate742(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate1261(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate1262(.a(gate216inter0), .b(s_102), .O(gate216inter1));
  and2  gate1263(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate1264(.a(s_102), .O(gate216inter3));
  inv1  gate1265(.a(s_103), .O(gate216inter4));
  nand2 gate1266(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate1267(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate1268(.a(G617), .O(gate216inter7));
  inv1  gate1269(.a(G675), .O(gate216inter8));
  nand2 gate1270(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate1271(.a(s_103), .b(gate216inter3), .O(gate216inter10));
  nor2  gate1272(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate1273(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate1274(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );

  xor2  gate1625(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate1626(.a(gate221inter0), .b(s_154), .O(gate221inter1));
  and2  gate1627(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate1628(.a(s_154), .O(gate221inter3));
  inv1  gate1629(.a(s_155), .O(gate221inter4));
  nand2 gate1630(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate1631(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate1632(.a(G622), .O(gate221inter7));
  inv1  gate1633(.a(G684), .O(gate221inter8));
  nand2 gate1634(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate1635(.a(s_155), .b(gate221inter3), .O(gate221inter10));
  nor2  gate1636(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate1637(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate1638(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate1779(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate1780(.a(gate224inter0), .b(s_176), .O(gate224inter1));
  and2  gate1781(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate1782(.a(s_176), .O(gate224inter3));
  inv1  gate1783(.a(s_177), .O(gate224inter4));
  nand2 gate1784(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate1785(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate1786(.a(G637), .O(gate224inter7));
  inv1  gate1787(.a(G687), .O(gate224inter8));
  nand2 gate1788(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate1789(.a(s_177), .b(gate224inter3), .O(gate224inter10));
  nor2  gate1790(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate1791(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate1792(.a(gate224inter12), .b(gate224inter1), .O(G705));

  xor2  gate1597(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate1598(.a(gate225inter0), .b(s_150), .O(gate225inter1));
  and2  gate1599(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate1600(.a(s_150), .O(gate225inter3));
  inv1  gate1601(.a(s_151), .O(gate225inter4));
  nand2 gate1602(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate1603(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate1604(.a(G690), .O(gate225inter7));
  inv1  gate1605(.a(G691), .O(gate225inter8));
  nand2 gate1606(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate1607(.a(s_151), .b(gate225inter3), .O(gate225inter10));
  nor2  gate1608(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate1609(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate1610(.a(gate225inter12), .b(gate225inter1), .O(G706));
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate2325(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate2326(.a(gate228inter0), .b(s_254), .O(gate228inter1));
  and2  gate2327(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate2328(.a(s_254), .O(gate228inter3));
  inv1  gate2329(.a(s_255), .O(gate228inter4));
  nand2 gate2330(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate2331(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate2332(.a(G696), .O(gate228inter7));
  inv1  gate2333(.a(G697), .O(gate228inter8));
  nand2 gate2334(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate2335(.a(s_255), .b(gate228inter3), .O(gate228inter10));
  nor2  gate2336(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate2337(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate2338(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate1793(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate1794(.a(gate231inter0), .b(s_178), .O(gate231inter1));
  and2  gate1795(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate1796(.a(s_178), .O(gate231inter3));
  inv1  gate1797(.a(s_179), .O(gate231inter4));
  nand2 gate1798(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate1799(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate1800(.a(G702), .O(gate231inter7));
  inv1  gate1801(.a(G703), .O(gate231inter8));
  nand2 gate1802(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate1803(.a(s_179), .b(gate231inter3), .O(gate231inter10));
  nor2  gate1804(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate1805(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate1806(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate1751(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate1752(.a(gate234inter0), .b(s_172), .O(gate234inter1));
  and2  gate1753(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate1754(.a(s_172), .O(gate234inter3));
  inv1  gate1755(.a(s_173), .O(gate234inter4));
  nand2 gate1756(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1757(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1758(.a(G245), .O(gate234inter7));
  inv1  gate1759(.a(G721), .O(gate234inter8));
  nand2 gate1760(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1761(.a(s_173), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1762(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1763(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1764(.a(gate234inter12), .b(gate234inter1), .O(G733));

  xor2  gate2255(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate2256(.a(gate235inter0), .b(s_244), .O(gate235inter1));
  and2  gate2257(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate2258(.a(s_244), .O(gate235inter3));
  inv1  gate2259(.a(s_245), .O(gate235inter4));
  nand2 gate2260(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate2261(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate2262(.a(G248), .O(gate235inter7));
  inv1  gate2263(.a(G724), .O(gate235inter8));
  nand2 gate2264(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate2265(.a(s_245), .b(gate235inter3), .O(gate235inter10));
  nor2  gate2266(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate2267(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate2268(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );

  xor2  gate715(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate716(.a(gate238inter0), .b(s_24), .O(gate238inter1));
  and2  gate717(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate718(.a(s_24), .O(gate238inter3));
  inv1  gate719(.a(s_25), .O(gate238inter4));
  nand2 gate720(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate721(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate722(.a(G257), .O(gate238inter7));
  inv1  gate723(.a(G709), .O(gate238inter8));
  nand2 gate724(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate725(.a(s_25), .b(gate238inter3), .O(gate238inter10));
  nor2  gate726(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate727(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate728(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate1485(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate1486(.a(gate240inter0), .b(s_134), .O(gate240inter1));
  and2  gate1487(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate1488(.a(s_134), .O(gate240inter3));
  inv1  gate1489(.a(s_135), .O(gate240inter4));
  nand2 gate1490(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate1491(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate1492(.a(G263), .O(gate240inter7));
  inv1  gate1493(.a(G715), .O(gate240inter8));
  nand2 gate1494(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate1495(.a(s_135), .b(gate240inter3), .O(gate240inter10));
  nor2  gate1496(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate1497(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate1498(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate2171(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate2172(.a(gate243inter0), .b(s_232), .O(gate243inter1));
  and2  gate2173(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate2174(.a(s_232), .O(gate243inter3));
  inv1  gate2175(.a(s_233), .O(gate243inter4));
  nand2 gate2176(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate2177(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate2178(.a(G245), .O(gate243inter7));
  inv1  gate2179(.a(G733), .O(gate243inter8));
  nand2 gate2180(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate2181(.a(s_233), .b(gate243inter3), .O(gate243inter10));
  nor2  gate2182(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate2183(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate2184(.a(gate243inter12), .b(gate243inter1), .O(G756));

  xor2  gate1415(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate1416(.a(gate244inter0), .b(s_124), .O(gate244inter1));
  and2  gate1417(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate1418(.a(s_124), .O(gate244inter3));
  inv1  gate1419(.a(s_125), .O(gate244inter4));
  nand2 gate1420(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate1421(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate1422(.a(G721), .O(gate244inter7));
  inv1  gate1423(.a(G733), .O(gate244inter8));
  nand2 gate1424(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate1425(.a(s_125), .b(gate244inter3), .O(gate244inter10));
  nor2  gate1426(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate1427(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate1428(.a(gate244inter12), .b(gate244inter1), .O(G757));

  xor2  gate2213(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate2214(.a(gate245inter0), .b(s_238), .O(gate245inter1));
  and2  gate2215(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate2216(.a(s_238), .O(gate245inter3));
  inv1  gate2217(.a(s_239), .O(gate245inter4));
  nand2 gate2218(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate2219(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate2220(.a(G248), .O(gate245inter7));
  inv1  gate2221(.a(G736), .O(gate245inter8));
  nand2 gate2222(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate2223(.a(s_239), .b(gate245inter3), .O(gate245inter10));
  nor2  gate2224(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate2225(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate2226(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );

  xor2  gate1807(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate1808(.a(gate251inter0), .b(s_180), .O(gate251inter1));
  and2  gate1809(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate1810(.a(s_180), .O(gate251inter3));
  inv1  gate1811(.a(s_181), .O(gate251inter4));
  nand2 gate1812(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate1813(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate1814(.a(G257), .O(gate251inter7));
  inv1  gate1815(.a(G745), .O(gate251inter8));
  nand2 gate1816(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate1817(.a(s_181), .b(gate251inter3), .O(gate251inter10));
  nor2  gate1818(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate1819(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate1820(.a(gate251inter12), .b(gate251inter1), .O(G764));
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );

  xor2  gate1009(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate1010(.a(gate254inter0), .b(s_66), .O(gate254inter1));
  and2  gate1011(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate1012(.a(s_66), .O(gate254inter3));
  inv1  gate1013(.a(s_67), .O(gate254inter4));
  nand2 gate1014(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate1015(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate1016(.a(G712), .O(gate254inter7));
  inv1  gate1017(.a(G748), .O(gate254inter8));
  nand2 gate1018(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate1019(.a(s_67), .b(gate254inter3), .O(gate254inter10));
  nor2  gate1020(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate1021(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate1022(.a(gate254inter12), .b(gate254inter1), .O(G767));
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate799(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate800(.a(gate258inter0), .b(s_36), .O(gate258inter1));
  and2  gate801(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate802(.a(s_36), .O(gate258inter3));
  inv1  gate803(.a(s_37), .O(gate258inter4));
  nand2 gate804(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate805(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate806(.a(G756), .O(gate258inter7));
  inv1  gate807(.a(G757), .O(gate258inter8));
  nand2 gate808(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate809(.a(s_37), .b(gate258inter3), .O(gate258inter10));
  nor2  gate810(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate811(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate812(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );

  xor2  gate2381(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate2382(.a(gate260inter0), .b(s_262), .O(gate260inter1));
  and2  gate2383(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate2384(.a(s_262), .O(gate260inter3));
  inv1  gate2385(.a(s_263), .O(gate260inter4));
  nand2 gate2386(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate2387(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate2388(.a(G760), .O(gate260inter7));
  inv1  gate2389(.a(G761), .O(gate260inter8));
  nand2 gate2390(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate2391(.a(s_263), .b(gate260inter3), .O(gate260inter10));
  nor2  gate2392(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate2393(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate2394(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate813(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate814(.a(gate266inter0), .b(s_38), .O(gate266inter1));
  and2  gate815(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate816(.a(s_38), .O(gate266inter3));
  inv1  gate817(.a(s_39), .O(gate266inter4));
  nand2 gate818(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate819(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate820(.a(G645), .O(gate266inter7));
  inv1  gate821(.a(G773), .O(gate266inter8));
  nand2 gate822(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate823(.a(s_39), .b(gate266inter3), .O(gate266inter10));
  nor2  gate824(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate825(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate826(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate1247(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate1248(.a(gate268inter0), .b(s_100), .O(gate268inter1));
  and2  gate1249(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate1250(.a(s_100), .O(gate268inter3));
  inv1  gate1251(.a(s_101), .O(gate268inter4));
  nand2 gate1252(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1253(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1254(.a(G651), .O(gate268inter7));
  inv1  gate1255(.a(G779), .O(gate268inter8));
  nand2 gate1256(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1257(.a(s_101), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1258(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1259(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1260(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate1947(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate1948(.a(gate271inter0), .b(s_200), .O(gate271inter1));
  and2  gate1949(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate1950(.a(s_200), .O(gate271inter3));
  inv1  gate1951(.a(s_201), .O(gate271inter4));
  nand2 gate1952(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate1953(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate1954(.a(G660), .O(gate271inter7));
  inv1  gate1955(.a(G788), .O(gate271inter8));
  nand2 gate1956(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate1957(.a(s_201), .b(gate271inter3), .O(gate271inter10));
  nor2  gate1958(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate1959(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate1960(.a(gate271inter12), .b(gate271inter1), .O(G812));

  xor2  gate1583(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate1584(.a(gate272inter0), .b(s_148), .O(gate272inter1));
  and2  gate1585(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate1586(.a(s_148), .O(gate272inter3));
  inv1  gate1587(.a(s_149), .O(gate272inter4));
  nand2 gate1588(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate1589(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate1590(.a(G663), .O(gate272inter7));
  inv1  gate1591(.a(G791), .O(gate272inter8));
  nand2 gate1592(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate1593(.a(s_149), .b(gate272inter3), .O(gate272inter10));
  nor2  gate1594(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate1595(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate1596(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate1961(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate1962(.a(gate274inter0), .b(s_202), .O(gate274inter1));
  and2  gate1963(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate1964(.a(s_202), .O(gate274inter3));
  inv1  gate1965(.a(s_203), .O(gate274inter4));
  nand2 gate1966(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate1967(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate1968(.a(G770), .O(gate274inter7));
  inv1  gate1969(.a(G794), .O(gate274inter8));
  nand2 gate1970(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate1971(.a(s_203), .b(gate274inter3), .O(gate274inter10));
  nor2  gate1972(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate1973(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate1974(.a(gate274inter12), .b(gate274inter1), .O(G819));

  xor2  gate1989(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate1990(.a(gate275inter0), .b(s_206), .O(gate275inter1));
  and2  gate1991(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate1992(.a(s_206), .O(gate275inter3));
  inv1  gate1993(.a(s_207), .O(gate275inter4));
  nand2 gate1994(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate1995(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate1996(.a(G645), .O(gate275inter7));
  inv1  gate1997(.a(G797), .O(gate275inter8));
  nand2 gate1998(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate1999(.a(s_207), .b(gate275inter3), .O(gate275inter10));
  nor2  gate2000(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate2001(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate2002(.a(gate275inter12), .b(gate275inter1), .O(G820));

  xor2  gate757(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate758(.a(gate276inter0), .b(s_30), .O(gate276inter1));
  and2  gate759(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate760(.a(s_30), .O(gate276inter3));
  inv1  gate761(.a(s_31), .O(gate276inter4));
  nand2 gate762(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate763(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate764(.a(G773), .O(gate276inter7));
  inv1  gate765(.a(G797), .O(gate276inter8));
  nand2 gate766(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate767(.a(s_31), .b(gate276inter3), .O(gate276inter10));
  nor2  gate768(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate769(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate770(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate2395(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate2396(.a(gate279inter0), .b(s_264), .O(gate279inter1));
  and2  gate2397(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate2398(.a(s_264), .O(gate279inter3));
  inv1  gate2399(.a(s_265), .O(gate279inter4));
  nand2 gate2400(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate2401(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate2402(.a(G651), .O(gate279inter7));
  inv1  gate2403(.a(G803), .O(gate279inter8));
  nand2 gate2404(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate2405(.a(s_265), .b(gate279inter3), .O(gate279inter10));
  nor2  gate2406(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate2407(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate2408(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );

  xor2  gate1667(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate1668(.a(gate281inter0), .b(s_160), .O(gate281inter1));
  and2  gate1669(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate1670(.a(s_160), .O(gate281inter3));
  inv1  gate1671(.a(s_161), .O(gate281inter4));
  nand2 gate1672(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate1673(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate1674(.a(G654), .O(gate281inter7));
  inv1  gate1675(.a(G806), .O(gate281inter8));
  nand2 gate1676(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate1677(.a(s_161), .b(gate281inter3), .O(gate281inter10));
  nor2  gate1678(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate1679(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate1680(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate1359(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate1360(.a(gate283inter0), .b(s_116), .O(gate283inter1));
  and2  gate1361(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate1362(.a(s_116), .O(gate283inter3));
  inv1  gate1363(.a(s_117), .O(gate283inter4));
  nand2 gate1364(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate1365(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate1366(.a(G657), .O(gate283inter7));
  inv1  gate1367(.a(G809), .O(gate283inter8));
  nand2 gate1368(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate1369(.a(s_117), .b(gate283inter3), .O(gate283inter10));
  nor2  gate1370(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate1371(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate1372(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate1205(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate1206(.a(gate286inter0), .b(s_94), .O(gate286inter1));
  and2  gate1207(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate1208(.a(s_94), .O(gate286inter3));
  inv1  gate1209(.a(s_95), .O(gate286inter4));
  nand2 gate1210(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate1211(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate1212(.a(G788), .O(gate286inter7));
  inv1  gate1213(.a(G812), .O(gate286inter8));
  nand2 gate1214(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate1215(.a(s_95), .b(gate286inter3), .O(gate286inter10));
  nor2  gate1216(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate1217(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate1218(.a(gate286inter12), .b(gate286inter1), .O(G831));
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate1191(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate1192(.a(gate288inter0), .b(s_92), .O(gate288inter1));
  and2  gate1193(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate1194(.a(s_92), .O(gate288inter3));
  inv1  gate1195(.a(s_93), .O(gate288inter4));
  nand2 gate1196(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate1197(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate1198(.a(G791), .O(gate288inter7));
  inv1  gate1199(.a(G815), .O(gate288inter8));
  nand2 gate1200(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate1201(.a(s_93), .b(gate288inter3), .O(gate288inter10));
  nor2  gate1202(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate1203(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate1204(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate1891(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate1892(.a(gate290inter0), .b(s_192), .O(gate290inter1));
  and2  gate1893(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate1894(.a(s_192), .O(gate290inter3));
  inv1  gate1895(.a(s_193), .O(gate290inter4));
  nand2 gate1896(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate1897(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate1898(.a(G820), .O(gate290inter7));
  inv1  gate1899(.a(G821), .O(gate290inter8));
  nand2 gate1900(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate1901(.a(s_193), .b(gate290inter3), .O(gate290inter10));
  nor2  gate1902(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate1903(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate1904(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate2353(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate2354(.a(gate293inter0), .b(s_258), .O(gate293inter1));
  and2  gate2355(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate2356(.a(s_258), .O(gate293inter3));
  inv1  gate2357(.a(s_259), .O(gate293inter4));
  nand2 gate2358(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate2359(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate2360(.a(G828), .O(gate293inter7));
  inv1  gate2361(.a(G829), .O(gate293inter8));
  nand2 gate2362(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate2363(.a(s_259), .b(gate293inter3), .O(gate293inter10));
  nor2  gate2364(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate2365(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate2366(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate897(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate898(.a(gate296inter0), .b(s_50), .O(gate296inter1));
  and2  gate899(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate900(.a(s_50), .O(gate296inter3));
  inv1  gate901(.a(s_51), .O(gate296inter4));
  nand2 gate902(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate903(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate904(.a(G826), .O(gate296inter7));
  inv1  gate905(.a(G827), .O(gate296inter8));
  nand2 gate906(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate907(.a(s_51), .b(gate296inter3), .O(gate296inter10));
  nor2  gate908(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate909(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate910(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate673(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate674(.a(gate393inter0), .b(s_18), .O(gate393inter1));
  and2  gate675(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate676(.a(s_18), .O(gate393inter3));
  inv1  gate677(.a(s_19), .O(gate393inter4));
  nand2 gate678(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate679(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate680(.a(G7), .O(gate393inter7));
  inv1  gate681(.a(G1054), .O(gate393inter8));
  nand2 gate682(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate683(.a(s_19), .b(gate393inter3), .O(gate393inter10));
  nor2  gate684(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate685(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate686(.a(gate393inter12), .b(gate393inter1), .O(G1150));

  xor2  gate925(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate926(.a(gate394inter0), .b(s_54), .O(gate394inter1));
  and2  gate927(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate928(.a(s_54), .O(gate394inter3));
  inv1  gate929(.a(s_55), .O(gate394inter4));
  nand2 gate930(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate931(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate932(.a(G8), .O(gate394inter7));
  inv1  gate933(.a(G1057), .O(gate394inter8));
  nand2 gate934(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate935(.a(s_55), .b(gate394inter3), .O(gate394inter10));
  nor2  gate936(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate937(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate938(.a(gate394inter12), .b(gate394inter1), .O(G1153));

  xor2  gate1499(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1500(.a(gate395inter0), .b(s_136), .O(gate395inter1));
  and2  gate1501(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1502(.a(s_136), .O(gate395inter3));
  inv1  gate1503(.a(s_137), .O(gate395inter4));
  nand2 gate1504(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1505(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1506(.a(G9), .O(gate395inter7));
  inv1  gate1507(.a(G1060), .O(gate395inter8));
  nand2 gate1508(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1509(.a(s_137), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1510(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1511(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1512(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate1611(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate1612(.a(gate400inter0), .b(s_152), .O(gate400inter1));
  and2  gate1613(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate1614(.a(s_152), .O(gate400inter3));
  inv1  gate1615(.a(s_153), .O(gate400inter4));
  nand2 gate1616(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate1617(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate1618(.a(G14), .O(gate400inter7));
  inv1  gate1619(.a(G1075), .O(gate400inter8));
  nand2 gate1620(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate1621(.a(s_153), .b(gate400inter3), .O(gate400inter10));
  nor2  gate1622(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate1623(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate1624(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate785(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate786(.a(gate402inter0), .b(s_34), .O(gate402inter1));
  and2  gate787(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate788(.a(s_34), .O(gate402inter3));
  inv1  gate789(.a(s_35), .O(gate402inter4));
  nand2 gate790(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate791(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate792(.a(G16), .O(gate402inter7));
  inv1  gate793(.a(G1081), .O(gate402inter8));
  nand2 gate794(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate795(.a(s_35), .b(gate402inter3), .O(gate402inter10));
  nor2  gate796(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate797(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate798(.a(gate402inter12), .b(gate402inter1), .O(G1177));
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );

  xor2  gate1317(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate1318(.a(gate405inter0), .b(s_110), .O(gate405inter1));
  and2  gate1319(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate1320(.a(s_110), .O(gate405inter3));
  inv1  gate1321(.a(s_111), .O(gate405inter4));
  nand2 gate1322(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate1323(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate1324(.a(G19), .O(gate405inter7));
  inv1  gate1325(.a(G1090), .O(gate405inter8));
  nand2 gate1326(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate1327(.a(s_111), .b(gate405inter3), .O(gate405inter10));
  nor2  gate1328(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate1329(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate1330(.a(gate405inter12), .b(gate405inter1), .O(G1186));
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate701(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate702(.a(gate407inter0), .b(s_22), .O(gate407inter1));
  and2  gate703(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate704(.a(s_22), .O(gate407inter3));
  inv1  gate705(.a(s_23), .O(gate407inter4));
  nand2 gate706(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate707(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate708(.a(G21), .O(gate407inter7));
  inv1  gate709(.a(G1096), .O(gate407inter8));
  nand2 gate710(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate711(.a(s_23), .b(gate407inter3), .O(gate407inter10));
  nor2  gate712(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate713(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate714(.a(gate407inter12), .b(gate407inter1), .O(G1192));

  xor2  gate1065(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate1066(.a(gate408inter0), .b(s_74), .O(gate408inter1));
  and2  gate1067(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate1068(.a(s_74), .O(gate408inter3));
  inv1  gate1069(.a(s_75), .O(gate408inter4));
  nand2 gate1070(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate1071(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate1072(.a(G22), .O(gate408inter7));
  inv1  gate1073(.a(G1099), .O(gate408inter8));
  nand2 gate1074(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate1075(.a(s_75), .b(gate408inter3), .O(gate408inter10));
  nor2  gate1076(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate1077(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate1078(.a(gate408inter12), .b(gate408inter1), .O(G1195));
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate1863(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate1864(.a(gate410inter0), .b(s_188), .O(gate410inter1));
  and2  gate1865(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate1866(.a(s_188), .O(gate410inter3));
  inv1  gate1867(.a(s_189), .O(gate410inter4));
  nand2 gate1868(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate1869(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate1870(.a(G24), .O(gate410inter7));
  inv1  gate1871(.a(G1105), .O(gate410inter8));
  nand2 gate1872(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate1873(.a(s_189), .b(gate410inter3), .O(gate410inter10));
  nor2  gate1874(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate1875(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate1876(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate1723(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate1724(.a(gate413inter0), .b(s_168), .O(gate413inter1));
  and2  gate1725(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate1726(.a(s_168), .O(gate413inter3));
  inv1  gate1727(.a(s_169), .O(gate413inter4));
  nand2 gate1728(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1729(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1730(.a(G27), .O(gate413inter7));
  inv1  gate1731(.a(G1114), .O(gate413inter8));
  nand2 gate1732(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1733(.a(s_169), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1734(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1735(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1736(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate1079(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate1080(.a(gate421inter0), .b(s_76), .O(gate421inter1));
  and2  gate1081(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate1082(.a(s_76), .O(gate421inter3));
  inv1  gate1083(.a(s_77), .O(gate421inter4));
  nand2 gate1084(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate1085(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate1086(.a(G2), .O(gate421inter7));
  inv1  gate1087(.a(G1135), .O(gate421inter8));
  nand2 gate1088(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate1089(.a(s_77), .b(gate421inter3), .O(gate421inter10));
  nor2  gate1090(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate1091(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate1092(.a(gate421inter12), .b(gate421inter1), .O(G1230));
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );

  xor2  gate561(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate562(.a(gate423inter0), .b(s_2), .O(gate423inter1));
  and2  gate563(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate564(.a(s_2), .O(gate423inter3));
  inv1  gate565(.a(s_3), .O(gate423inter4));
  nand2 gate566(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate567(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate568(.a(G3), .O(gate423inter7));
  inv1  gate569(.a(G1138), .O(gate423inter8));
  nand2 gate570(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate571(.a(s_3), .b(gate423inter3), .O(gate423inter10));
  nor2  gate572(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate573(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate574(.a(gate423inter12), .b(gate423inter1), .O(G1232));
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate645(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate646(.a(gate428inter0), .b(s_14), .O(gate428inter1));
  and2  gate647(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate648(.a(s_14), .O(gate428inter3));
  inv1  gate649(.a(s_15), .O(gate428inter4));
  nand2 gate650(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate651(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate652(.a(G1048), .O(gate428inter7));
  inv1  gate653(.a(G1144), .O(gate428inter8));
  nand2 gate654(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate655(.a(s_15), .b(gate428inter3), .O(gate428inter10));
  nor2  gate656(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate657(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate658(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate1849(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate1850(.a(gate431inter0), .b(s_186), .O(gate431inter1));
  and2  gate1851(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate1852(.a(s_186), .O(gate431inter3));
  inv1  gate1853(.a(s_187), .O(gate431inter4));
  nand2 gate1854(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate1855(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate1856(.a(G7), .O(gate431inter7));
  inv1  gate1857(.a(G1150), .O(gate431inter8));
  nand2 gate1858(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate1859(.a(s_187), .b(gate431inter3), .O(gate431inter10));
  nor2  gate1860(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate1861(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate1862(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );

  xor2  gate883(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate884(.a(gate436inter0), .b(s_48), .O(gate436inter1));
  and2  gate885(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate886(.a(s_48), .O(gate436inter3));
  inv1  gate887(.a(s_49), .O(gate436inter4));
  nand2 gate888(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate889(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate890(.a(G1060), .O(gate436inter7));
  inv1  gate891(.a(G1156), .O(gate436inter8));
  nand2 gate892(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate893(.a(s_49), .b(gate436inter3), .O(gate436inter10));
  nor2  gate894(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate895(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate896(.a(gate436inter12), .b(gate436inter1), .O(G1245));
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate1289(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate1290(.a(gate438inter0), .b(s_106), .O(gate438inter1));
  and2  gate1291(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate1292(.a(s_106), .O(gate438inter3));
  inv1  gate1293(.a(s_107), .O(gate438inter4));
  nand2 gate1294(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate1295(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate1296(.a(G1063), .O(gate438inter7));
  inv1  gate1297(.a(G1159), .O(gate438inter8));
  nand2 gate1298(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate1299(.a(s_107), .b(gate438inter3), .O(gate438inter10));
  nor2  gate1300(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate1301(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate1302(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate2297(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate2298(.a(gate441inter0), .b(s_250), .O(gate441inter1));
  and2  gate2299(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate2300(.a(s_250), .O(gate441inter3));
  inv1  gate2301(.a(s_251), .O(gate441inter4));
  nand2 gate2302(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate2303(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate2304(.a(G12), .O(gate441inter7));
  inv1  gate2305(.a(G1165), .O(gate441inter8));
  nand2 gate2306(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate2307(.a(s_251), .b(gate441inter3), .O(gate441inter10));
  nor2  gate2308(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate2309(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate2310(.a(gate441inter12), .b(gate441inter1), .O(G1250));

  xor2  gate2073(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate2074(.a(gate442inter0), .b(s_218), .O(gate442inter1));
  and2  gate2075(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate2076(.a(s_218), .O(gate442inter3));
  inv1  gate2077(.a(s_219), .O(gate442inter4));
  nand2 gate2078(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate2079(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate2080(.a(G1069), .O(gate442inter7));
  inv1  gate2081(.a(G1165), .O(gate442inter8));
  nand2 gate2082(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate2083(.a(s_219), .b(gate442inter3), .O(gate442inter10));
  nor2  gate2084(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate2085(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate2086(.a(gate442inter12), .b(gate442inter1), .O(G1251));

  xor2  gate1345(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate1346(.a(gate443inter0), .b(s_114), .O(gate443inter1));
  and2  gate1347(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate1348(.a(s_114), .O(gate443inter3));
  inv1  gate1349(.a(s_115), .O(gate443inter4));
  nand2 gate1350(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate1351(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate1352(.a(G13), .O(gate443inter7));
  inv1  gate1353(.a(G1168), .O(gate443inter8));
  nand2 gate1354(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate1355(.a(s_115), .b(gate443inter3), .O(gate443inter10));
  nor2  gate1356(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate1357(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate1358(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate1933(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate1934(.a(gate456inter0), .b(s_198), .O(gate456inter1));
  and2  gate1935(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate1936(.a(s_198), .O(gate456inter3));
  inv1  gate1937(.a(s_199), .O(gate456inter4));
  nand2 gate1938(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate1939(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate1940(.a(G1090), .O(gate456inter7));
  inv1  gate1941(.a(G1186), .O(gate456inter8));
  nand2 gate1942(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate1943(.a(s_199), .b(gate456inter3), .O(gate456inter10));
  nor2  gate1944(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate1945(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate1946(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate1331(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate1332(.a(gate459inter0), .b(s_112), .O(gate459inter1));
  and2  gate1333(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate1334(.a(s_112), .O(gate459inter3));
  inv1  gate1335(.a(s_113), .O(gate459inter4));
  nand2 gate1336(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate1337(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate1338(.a(G21), .O(gate459inter7));
  inv1  gate1339(.a(G1192), .O(gate459inter8));
  nand2 gate1340(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate1341(.a(s_113), .b(gate459inter3), .O(gate459inter10));
  nor2  gate1342(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate1343(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate1344(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate2059(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate2060(.a(gate461inter0), .b(s_216), .O(gate461inter1));
  and2  gate2061(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate2062(.a(s_216), .O(gate461inter3));
  inv1  gate2063(.a(s_217), .O(gate461inter4));
  nand2 gate2064(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate2065(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate2066(.a(G22), .O(gate461inter7));
  inv1  gate2067(.a(G1195), .O(gate461inter8));
  nand2 gate2068(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate2069(.a(s_217), .b(gate461inter3), .O(gate461inter10));
  nor2  gate2070(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate2071(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate2072(.a(gate461inter12), .b(gate461inter1), .O(G1270));

  xor2  gate2367(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate2368(.a(gate462inter0), .b(s_260), .O(gate462inter1));
  and2  gate2369(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate2370(.a(s_260), .O(gate462inter3));
  inv1  gate2371(.a(s_261), .O(gate462inter4));
  nand2 gate2372(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate2373(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate2374(.a(G1099), .O(gate462inter7));
  inv1  gate2375(.a(G1195), .O(gate462inter8));
  nand2 gate2376(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate2377(.a(s_261), .b(gate462inter3), .O(gate462inter10));
  nor2  gate2378(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate2379(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate2380(.a(gate462inter12), .b(gate462inter1), .O(G1271));

  xor2  gate981(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate982(.a(gate463inter0), .b(s_62), .O(gate463inter1));
  and2  gate983(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate984(.a(s_62), .O(gate463inter3));
  inv1  gate985(.a(s_63), .O(gate463inter4));
  nand2 gate986(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate987(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate988(.a(G23), .O(gate463inter7));
  inv1  gate989(.a(G1198), .O(gate463inter8));
  nand2 gate990(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate991(.a(s_63), .b(gate463inter3), .O(gate463inter10));
  nor2  gate992(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate993(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate994(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate1653(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate1654(.a(gate466inter0), .b(s_158), .O(gate466inter1));
  and2  gate1655(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate1656(.a(s_158), .O(gate466inter3));
  inv1  gate1657(.a(s_159), .O(gate466inter4));
  nand2 gate1658(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate1659(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate1660(.a(G1105), .O(gate466inter7));
  inv1  gate1661(.a(G1201), .O(gate466inter8));
  nand2 gate1662(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate1663(.a(s_159), .b(gate466inter3), .O(gate466inter10));
  nor2  gate1664(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate1665(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate1666(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );

  xor2  gate687(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate688(.a(gate468inter0), .b(s_20), .O(gate468inter1));
  and2  gate689(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate690(.a(s_20), .O(gate468inter3));
  inv1  gate691(.a(s_21), .O(gate468inter4));
  nand2 gate692(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate693(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate694(.a(G1108), .O(gate468inter7));
  inv1  gate695(.a(G1204), .O(gate468inter8));
  nand2 gate696(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate697(.a(s_21), .b(gate468inter3), .O(gate468inter10));
  nor2  gate698(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate699(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate700(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );

  xor2  gate967(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate968(.a(gate473inter0), .b(s_60), .O(gate473inter1));
  and2  gate969(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate970(.a(s_60), .O(gate473inter3));
  inv1  gate971(.a(s_61), .O(gate473inter4));
  nand2 gate972(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate973(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate974(.a(G28), .O(gate473inter7));
  inv1  gate975(.a(G1213), .O(gate473inter8));
  nand2 gate976(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate977(.a(s_61), .b(gate473inter3), .O(gate473inter10));
  nor2  gate978(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate979(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate980(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate1639(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate1640(.a(gate476inter0), .b(s_156), .O(gate476inter1));
  and2  gate1641(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate1642(.a(s_156), .O(gate476inter3));
  inv1  gate1643(.a(s_157), .O(gate476inter4));
  nand2 gate1644(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate1645(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate1646(.a(G1120), .O(gate476inter7));
  inv1  gate1647(.a(G1216), .O(gate476inter8));
  nand2 gate1648(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate1649(.a(s_157), .b(gate476inter3), .O(gate476inter10));
  nor2  gate1650(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate1651(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate1652(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );

  xor2  gate1233(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate1234(.a(gate478inter0), .b(s_98), .O(gate478inter1));
  and2  gate1235(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate1236(.a(s_98), .O(gate478inter3));
  inv1  gate1237(.a(s_99), .O(gate478inter4));
  nand2 gate1238(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate1239(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate1240(.a(G1123), .O(gate478inter7));
  inv1  gate1241(.a(G1219), .O(gate478inter8));
  nand2 gate1242(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate1243(.a(s_99), .b(gate478inter3), .O(gate478inter10));
  nor2  gate1244(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate1245(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate1246(.a(gate478inter12), .b(gate478inter1), .O(G1287));

  xor2  gate1275(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate1276(.a(gate479inter0), .b(s_104), .O(gate479inter1));
  and2  gate1277(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate1278(.a(s_104), .O(gate479inter3));
  inv1  gate1279(.a(s_105), .O(gate479inter4));
  nand2 gate1280(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate1281(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate1282(.a(G31), .O(gate479inter7));
  inv1  gate1283(.a(G1222), .O(gate479inter8));
  nand2 gate1284(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate1285(.a(s_105), .b(gate479inter3), .O(gate479inter10));
  nor2  gate1286(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate1287(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate1288(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate1471(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate1472(.a(gate481inter0), .b(s_132), .O(gate481inter1));
  and2  gate1473(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate1474(.a(s_132), .O(gate481inter3));
  inv1  gate1475(.a(s_133), .O(gate481inter4));
  nand2 gate1476(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate1477(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate1478(.a(G32), .O(gate481inter7));
  inv1  gate1479(.a(G1225), .O(gate481inter8));
  nand2 gate1480(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate1481(.a(s_133), .b(gate481inter3), .O(gate481inter10));
  nor2  gate1482(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate1483(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate1484(.a(gate481inter12), .b(gate481inter1), .O(G1290));
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate1527(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate1528(.a(gate486inter0), .b(s_140), .O(gate486inter1));
  and2  gate1529(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate1530(.a(s_140), .O(gate486inter3));
  inv1  gate1531(.a(s_141), .O(gate486inter4));
  nand2 gate1532(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate1533(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate1534(.a(G1234), .O(gate486inter7));
  inv1  gate1535(.a(G1235), .O(gate486inter8));
  nand2 gate1536(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate1537(.a(s_141), .b(gate486inter3), .O(gate486inter10));
  nor2  gate1538(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate1539(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate1540(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate911(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate912(.a(gate488inter0), .b(s_52), .O(gate488inter1));
  and2  gate913(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate914(.a(s_52), .O(gate488inter3));
  inv1  gate915(.a(s_53), .O(gate488inter4));
  nand2 gate916(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate917(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate918(.a(G1238), .O(gate488inter7));
  inv1  gate919(.a(G1239), .O(gate488inter8));
  nand2 gate920(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate921(.a(s_53), .b(gate488inter3), .O(gate488inter10));
  nor2  gate922(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate923(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate924(.a(gate488inter12), .b(gate488inter1), .O(G1297));

  xor2  gate869(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate870(.a(gate489inter0), .b(s_46), .O(gate489inter1));
  and2  gate871(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate872(.a(s_46), .O(gate489inter3));
  inv1  gate873(.a(s_47), .O(gate489inter4));
  nand2 gate874(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate875(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate876(.a(G1240), .O(gate489inter7));
  inv1  gate877(.a(G1241), .O(gate489inter8));
  nand2 gate878(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate879(.a(s_47), .b(gate489inter3), .O(gate489inter10));
  nor2  gate880(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate881(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate882(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate2129(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate2130(.a(gate492inter0), .b(s_226), .O(gate492inter1));
  and2  gate2131(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate2132(.a(s_226), .O(gate492inter3));
  inv1  gate2133(.a(s_227), .O(gate492inter4));
  nand2 gate2134(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate2135(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate2136(.a(G1246), .O(gate492inter7));
  inv1  gate2137(.a(G1247), .O(gate492inter8));
  nand2 gate2138(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate2139(.a(s_227), .b(gate492inter3), .O(gate492inter10));
  nor2  gate2140(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate2141(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate2142(.a(gate492inter12), .b(gate492inter1), .O(G1301));
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate1163(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1164(.a(gate494inter0), .b(s_88), .O(gate494inter1));
  and2  gate1165(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1166(.a(s_88), .O(gate494inter3));
  inv1  gate1167(.a(s_89), .O(gate494inter4));
  nand2 gate1168(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1169(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1170(.a(G1250), .O(gate494inter7));
  inv1  gate1171(.a(G1251), .O(gate494inter8));
  nand2 gate1172(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1173(.a(s_89), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1174(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1175(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1176(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate827(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate828(.a(gate499inter0), .b(s_40), .O(gate499inter1));
  and2  gate829(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate830(.a(s_40), .O(gate499inter3));
  inv1  gate831(.a(s_41), .O(gate499inter4));
  nand2 gate832(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate833(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate834(.a(G1260), .O(gate499inter7));
  inv1  gate835(.a(G1261), .O(gate499inter8));
  nand2 gate836(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate837(.a(s_41), .b(gate499inter3), .O(gate499inter10));
  nor2  gate838(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate839(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate840(.a(gate499inter12), .b(gate499inter1), .O(G1308));

  xor2  gate1429(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate1430(.a(gate500inter0), .b(s_126), .O(gate500inter1));
  and2  gate1431(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate1432(.a(s_126), .O(gate500inter3));
  inv1  gate1433(.a(s_127), .O(gate500inter4));
  nand2 gate1434(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate1435(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate1436(.a(G1262), .O(gate500inter7));
  inv1  gate1437(.a(G1263), .O(gate500inter8));
  nand2 gate1438(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate1439(.a(s_127), .b(gate500inter3), .O(gate500inter10));
  nor2  gate1440(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate1441(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate1442(.a(gate500inter12), .b(gate500inter1), .O(G1309));

  xor2  gate1373(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate1374(.a(gate501inter0), .b(s_118), .O(gate501inter1));
  and2  gate1375(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate1376(.a(s_118), .O(gate501inter3));
  inv1  gate1377(.a(s_119), .O(gate501inter4));
  nand2 gate1378(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1379(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1380(.a(G1264), .O(gate501inter7));
  inv1  gate1381(.a(G1265), .O(gate501inter8));
  nand2 gate1382(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1383(.a(s_119), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1384(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1385(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1386(.a(gate501inter12), .b(gate501inter1), .O(G1310));

  xor2  gate2017(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate2018(.a(gate502inter0), .b(s_210), .O(gate502inter1));
  and2  gate2019(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate2020(.a(s_210), .O(gate502inter3));
  inv1  gate2021(.a(s_211), .O(gate502inter4));
  nand2 gate2022(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate2023(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate2024(.a(G1266), .O(gate502inter7));
  inv1  gate2025(.a(G1267), .O(gate502inter8));
  nand2 gate2026(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate2027(.a(s_211), .b(gate502inter3), .O(gate502inter10));
  nor2  gate2028(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate2029(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate2030(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate2269(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate2270(.a(gate504inter0), .b(s_246), .O(gate504inter1));
  and2  gate2271(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate2272(.a(s_246), .O(gate504inter3));
  inv1  gate2273(.a(s_247), .O(gate504inter4));
  nand2 gate2274(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate2275(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate2276(.a(G1270), .O(gate504inter7));
  inv1  gate2277(.a(G1271), .O(gate504inter8));
  nand2 gate2278(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate2279(.a(s_247), .b(gate504inter3), .O(gate504inter10));
  nor2  gate2280(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate2281(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate2282(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate2045(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate2046(.a(gate509inter0), .b(s_214), .O(gate509inter1));
  and2  gate2047(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate2048(.a(s_214), .O(gate509inter3));
  inv1  gate2049(.a(s_215), .O(gate509inter4));
  nand2 gate2050(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate2051(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate2052(.a(G1280), .O(gate509inter7));
  inv1  gate2053(.a(G1281), .O(gate509inter8));
  nand2 gate2054(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate2055(.a(s_215), .b(gate509inter3), .O(gate509inter10));
  nor2  gate2056(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate2057(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate2058(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );

  xor2  gate2423(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate2424(.a(gate512inter0), .b(s_268), .O(gate512inter1));
  and2  gate2425(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate2426(.a(s_268), .O(gate512inter3));
  inv1  gate2427(.a(s_269), .O(gate512inter4));
  nand2 gate2428(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate2429(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate2430(.a(G1286), .O(gate512inter7));
  inv1  gate2431(.a(G1287), .O(gate512inter8));
  nand2 gate2432(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate2433(.a(s_269), .b(gate512inter3), .O(gate512inter10));
  nor2  gate2434(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate2435(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate2436(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule