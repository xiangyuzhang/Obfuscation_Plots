module c499 (N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
             N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
             N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
             N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
             N137,N724,N725,N726,N727,N728,N729,N730,N731,N732,
             N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,
             N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,
             N753,N754,N755);
input N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
      N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
      N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
      N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
      N137;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61;
output N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,
       N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
       N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
       N754,N755;
wire N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
     N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
     N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,
     N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,
     N290,N293,N296,N299,N302,N305,N308,N311,N314,N315,
     N316,N317,N318,N319,N320,N321,N338,N339,N340,N341,
     N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,
     N352,N353,N354,N367,N380,N393,N406,N419,N432,N445,
     N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
     N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,
     N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,
     N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,
     N594,N595,N596,N597,N598,N599,N600,N601,N602,N607,
     N620,N625,N630,N635,N640,N645,N650,N655,N692,N693,
     N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,
     N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,
     N714,N715,N716,N717,N718,N719,N720,N721,N722,N723, gate2inter0, gate2inter1, gate2inter2, gate2inter3, gate2inter4, gate2inter5, gate2inter6, gate2inter7, gate2inter8, gate2inter9, gate2inter10, gate2inter11, gate2inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate8inter0, gate8inter1, gate8inter2, gate8inter3, gate8inter4, gate8inter5, gate8inter6, gate8inter7, gate8inter8, gate8inter9, gate8inter10, gate8inter11, gate8inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12;


xor2 gate1( .a(N1), .b(N5), .O(N250) );

  xor2  gate203(.a(N13), .b(N9), .O(gate2inter0));
  nand2 gate204(.a(gate2inter0), .b(s_0), .O(gate2inter1));
  and2  gate205(.a(N13), .b(N9), .O(gate2inter2));
  inv1  gate206(.a(s_0), .O(gate2inter3));
  inv1  gate207(.a(s_1), .O(gate2inter4));
  nand2 gate208(.a(gate2inter4), .b(gate2inter3), .O(gate2inter5));
  nor2  gate209(.a(gate2inter5), .b(gate2inter2), .O(gate2inter6));
  inv1  gate210(.a(N9), .O(gate2inter7));
  inv1  gate211(.a(N13), .O(gate2inter8));
  nand2 gate212(.a(gate2inter8), .b(gate2inter7), .O(gate2inter9));
  nand2 gate213(.a(s_1), .b(gate2inter3), .O(gate2inter10));
  nor2  gate214(.a(gate2inter10), .b(gate2inter9), .O(gate2inter11));
  nor2  gate215(.a(gate2inter11), .b(gate2inter6), .O(gate2inter12));
  nand2 gate216(.a(gate2inter12), .b(gate2inter1), .O(N251));
xor2 gate3( .a(N17), .b(N21), .O(N252) );
xor2 gate4( .a(N25), .b(N29), .O(N253) );
xor2 gate5( .a(N33), .b(N37), .O(N254) );
xor2 gate6( .a(N41), .b(N45), .O(N255) );
xor2 gate7( .a(N49), .b(N53), .O(N256) );

  xor2  gate483(.a(N61), .b(N57), .O(gate8inter0));
  nand2 gate484(.a(gate8inter0), .b(s_40), .O(gate8inter1));
  and2  gate485(.a(N61), .b(N57), .O(gate8inter2));
  inv1  gate486(.a(s_40), .O(gate8inter3));
  inv1  gate487(.a(s_41), .O(gate8inter4));
  nand2 gate488(.a(gate8inter4), .b(gate8inter3), .O(gate8inter5));
  nor2  gate489(.a(gate8inter5), .b(gate8inter2), .O(gate8inter6));
  inv1  gate490(.a(N57), .O(gate8inter7));
  inv1  gate491(.a(N61), .O(gate8inter8));
  nand2 gate492(.a(gate8inter8), .b(gate8inter7), .O(gate8inter9));
  nand2 gate493(.a(s_41), .b(gate8inter3), .O(gate8inter10));
  nor2  gate494(.a(gate8inter10), .b(gate8inter9), .O(gate8inter11));
  nor2  gate495(.a(gate8inter11), .b(gate8inter6), .O(gate8inter12));
  nand2 gate496(.a(gate8inter12), .b(gate8inter1), .O(N257));

  xor2  gate273(.a(N69), .b(N65), .O(gate9inter0));
  nand2 gate274(.a(gate9inter0), .b(s_10), .O(gate9inter1));
  and2  gate275(.a(N69), .b(N65), .O(gate9inter2));
  inv1  gate276(.a(s_10), .O(gate9inter3));
  inv1  gate277(.a(s_11), .O(gate9inter4));
  nand2 gate278(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate279(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate280(.a(N65), .O(gate9inter7));
  inv1  gate281(.a(N69), .O(gate9inter8));
  nand2 gate282(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate283(.a(s_11), .b(gate9inter3), .O(gate9inter10));
  nor2  gate284(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate285(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate286(.a(gate9inter12), .b(gate9inter1), .O(N258));
xor2 gate10( .a(N73), .b(N77), .O(N259) );
xor2 gate11( .a(N81), .b(N85), .O(N260) );
xor2 gate12( .a(N89), .b(N93), .O(N261) );
xor2 gate13( .a(N97), .b(N101), .O(N262) );

  xor2  gate525(.a(N109), .b(N105), .O(gate14inter0));
  nand2 gate526(.a(gate14inter0), .b(s_46), .O(gate14inter1));
  and2  gate527(.a(N109), .b(N105), .O(gate14inter2));
  inv1  gate528(.a(s_46), .O(gate14inter3));
  inv1  gate529(.a(s_47), .O(gate14inter4));
  nand2 gate530(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate531(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate532(.a(N105), .O(gate14inter7));
  inv1  gate533(.a(N109), .O(gate14inter8));
  nand2 gate534(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate535(.a(s_47), .b(gate14inter3), .O(gate14inter10));
  nor2  gate536(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate537(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate538(.a(gate14inter12), .b(gate14inter1), .O(N263));
xor2 gate15( .a(N113), .b(N117), .O(N264) );
xor2 gate16( .a(N121), .b(N125), .O(N265) );
and2 gate17( .a(N129), .b(N137), .O(N266) );
and2 gate18( .a(N130), .b(N137), .O(N267) );
and2 gate19( .a(N131), .b(N137), .O(N268) );
and2 gate20( .a(N132), .b(N137), .O(N269) );
and2 gate21( .a(N133), .b(N137), .O(N270) );
and2 gate22( .a(N134), .b(N137), .O(N271) );
and2 gate23( .a(N135), .b(N137), .O(N272) );
and2 gate24( .a(N136), .b(N137), .O(N273) );
xor2 gate25( .a(N1), .b(N17), .O(N274) );

  xor2  gate399(.a(N49), .b(N33), .O(gate26inter0));
  nand2 gate400(.a(gate26inter0), .b(s_28), .O(gate26inter1));
  and2  gate401(.a(N49), .b(N33), .O(gate26inter2));
  inv1  gate402(.a(s_28), .O(gate26inter3));
  inv1  gate403(.a(s_29), .O(gate26inter4));
  nand2 gate404(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate405(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate406(.a(N33), .O(gate26inter7));
  inv1  gate407(.a(N49), .O(gate26inter8));
  nand2 gate408(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate409(.a(s_29), .b(gate26inter3), .O(gate26inter10));
  nor2  gate410(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate411(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate412(.a(gate26inter12), .b(gate26inter1), .O(N275));
xor2 gate27( .a(N5), .b(N21), .O(N276) );

  xor2  gate581(.a(N53), .b(N37), .O(gate28inter0));
  nand2 gate582(.a(gate28inter0), .b(s_54), .O(gate28inter1));
  and2  gate583(.a(N53), .b(N37), .O(gate28inter2));
  inv1  gate584(.a(s_54), .O(gate28inter3));
  inv1  gate585(.a(s_55), .O(gate28inter4));
  nand2 gate586(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate587(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate588(.a(N37), .O(gate28inter7));
  inv1  gate589(.a(N53), .O(gate28inter8));
  nand2 gate590(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate591(.a(s_55), .b(gate28inter3), .O(gate28inter10));
  nor2  gate592(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate593(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate594(.a(gate28inter12), .b(gate28inter1), .O(N277));
xor2 gate29( .a(N9), .b(N25), .O(N278) );

  xor2  gate301(.a(N57), .b(N41), .O(gate30inter0));
  nand2 gate302(.a(gate30inter0), .b(s_14), .O(gate30inter1));
  and2  gate303(.a(N57), .b(N41), .O(gate30inter2));
  inv1  gate304(.a(s_14), .O(gate30inter3));
  inv1  gate305(.a(s_15), .O(gate30inter4));
  nand2 gate306(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate307(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate308(.a(N41), .O(gate30inter7));
  inv1  gate309(.a(N57), .O(gate30inter8));
  nand2 gate310(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate311(.a(s_15), .b(gate30inter3), .O(gate30inter10));
  nor2  gate312(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate313(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate314(.a(gate30inter12), .b(gate30inter1), .O(N279));
xor2 gate31( .a(N13), .b(N29), .O(N280) );
xor2 gate32( .a(N45), .b(N61), .O(N281) );
xor2 gate33( .a(N65), .b(N81), .O(N282) );
xor2 gate34( .a(N97), .b(N113), .O(N283) );

  xor2  gate567(.a(N85), .b(N69), .O(gate35inter0));
  nand2 gate568(.a(gate35inter0), .b(s_52), .O(gate35inter1));
  and2  gate569(.a(N85), .b(N69), .O(gate35inter2));
  inv1  gate570(.a(s_52), .O(gate35inter3));
  inv1  gate571(.a(s_53), .O(gate35inter4));
  nand2 gate572(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate573(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate574(.a(N69), .O(gate35inter7));
  inv1  gate575(.a(N85), .O(gate35inter8));
  nand2 gate576(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate577(.a(s_53), .b(gate35inter3), .O(gate35inter10));
  nor2  gate578(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate579(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate580(.a(gate35inter12), .b(gate35inter1), .O(N284));
xor2 gate36( .a(N101), .b(N117), .O(N285) );

  xor2  gate469(.a(N89), .b(N73), .O(gate37inter0));
  nand2 gate470(.a(gate37inter0), .b(s_38), .O(gate37inter1));
  and2  gate471(.a(N89), .b(N73), .O(gate37inter2));
  inv1  gate472(.a(s_38), .O(gate37inter3));
  inv1  gate473(.a(s_39), .O(gate37inter4));
  nand2 gate474(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate475(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate476(.a(N73), .O(gate37inter7));
  inv1  gate477(.a(N89), .O(gate37inter8));
  nand2 gate478(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate479(.a(s_39), .b(gate37inter3), .O(gate37inter10));
  nor2  gate480(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate481(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate482(.a(gate37inter12), .b(gate37inter1), .O(N286));
xor2 gate38( .a(N105), .b(N121), .O(N287) );
xor2 gate39( .a(N77), .b(N93), .O(N288) );
xor2 gate40( .a(N109), .b(N125), .O(N289) );
xor2 gate41( .a(N250), .b(N251), .O(N290) );

  xor2  gate329(.a(N253), .b(N252), .O(gate42inter0));
  nand2 gate330(.a(gate42inter0), .b(s_18), .O(gate42inter1));
  and2  gate331(.a(N253), .b(N252), .O(gate42inter2));
  inv1  gate332(.a(s_18), .O(gate42inter3));
  inv1  gate333(.a(s_19), .O(gate42inter4));
  nand2 gate334(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate335(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate336(.a(N252), .O(gate42inter7));
  inv1  gate337(.a(N253), .O(gate42inter8));
  nand2 gate338(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate339(.a(s_19), .b(gate42inter3), .O(gate42inter10));
  nor2  gate340(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate341(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate342(.a(gate42inter12), .b(gate42inter1), .O(N293));

  xor2  gate231(.a(N255), .b(N254), .O(gate43inter0));
  nand2 gate232(.a(gate43inter0), .b(s_4), .O(gate43inter1));
  and2  gate233(.a(N255), .b(N254), .O(gate43inter2));
  inv1  gate234(.a(s_4), .O(gate43inter3));
  inv1  gate235(.a(s_5), .O(gate43inter4));
  nand2 gate236(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate237(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate238(.a(N254), .O(gate43inter7));
  inv1  gate239(.a(N255), .O(gate43inter8));
  nand2 gate240(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate241(.a(s_5), .b(gate43inter3), .O(gate43inter10));
  nor2  gate242(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate243(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate244(.a(gate43inter12), .b(gate43inter1), .O(N296));
xor2 gate44( .a(N256), .b(N257), .O(N299) );
xor2 gate45( .a(N258), .b(N259), .O(N302) );

  xor2  gate553(.a(N261), .b(N260), .O(gate46inter0));
  nand2 gate554(.a(gate46inter0), .b(s_50), .O(gate46inter1));
  and2  gate555(.a(N261), .b(N260), .O(gate46inter2));
  inv1  gate556(.a(s_50), .O(gate46inter3));
  inv1  gate557(.a(s_51), .O(gate46inter4));
  nand2 gate558(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate559(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate560(.a(N260), .O(gate46inter7));
  inv1  gate561(.a(N261), .O(gate46inter8));
  nand2 gate562(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate563(.a(s_51), .b(gate46inter3), .O(gate46inter10));
  nor2  gate564(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate565(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate566(.a(gate46inter12), .b(gate46inter1), .O(N305));
xor2 gate47( .a(N262), .b(N263), .O(N308) );
xor2 gate48( .a(N264), .b(N265), .O(N311) );
xor2 gate49( .a(N274), .b(N275), .O(N314) );

  xor2  gate245(.a(N277), .b(N276), .O(gate50inter0));
  nand2 gate246(.a(gate50inter0), .b(s_6), .O(gate50inter1));
  and2  gate247(.a(N277), .b(N276), .O(gate50inter2));
  inv1  gate248(.a(s_6), .O(gate50inter3));
  inv1  gate249(.a(s_7), .O(gate50inter4));
  nand2 gate250(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate251(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate252(.a(N276), .O(gate50inter7));
  inv1  gate253(.a(N277), .O(gate50inter8));
  nand2 gate254(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate255(.a(s_7), .b(gate50inter3), .O(gate50inter10));
  nor2  gate256(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate257(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate258(.a(gate50inter12), .b(gate50inter1), .O(N315));
xor2 gate51( .a(N278), .b(N279), .O(N316) );
xor2 gate52( .a(N280), .b(N281), .O(N317) );
xor2 gate53( .a(N282), .b(N283), .O(N318) );

  xor2  gate315(.a(N285), .b(N284), .O(gate54inter0));
  nand2 gate316(.a(gate54inter0), .b(s_16), .O(gate54inter1));
  and2  gate317(.a(N285), .b(N284), .O(gate54inter2));
  inv1  gate318(.a(s_16), .O(gate54inter3));
  inv1  gate319(.a(s_17), .O(gate54inter4));
  nand2 gate320(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate321(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate322(.a(N284), .O(gate54inter7));
  inv1  gate323(.a(N285), .O(gate54inter8));
  nand2 gate324(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate325(.a(s_17), .b(gate54inter3), .O(gate54inter10));
  nor2  gate326(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate327(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate328(.a(gate54inter12), .b(gate54inter1), .O(N319));

  xor2  gate609(.a(N287), .b(N286), .O(gate55inter0));
  nand2 gate610(.a(gate55inter0), .b(s_58), .O(gate55inter1));
  and2  gate611(.a(N287), .b(N286), .O(gate55inter2));
  inv1  gate612(.a(s_58), .O(gate55inter3));
  inv1  gate613(.a(s_59), .O(gate55inter4));
  nand2 gate614(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate615(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate616(.a(N286), .O(gate55inter7));
  inv1  gate617(.a(N287), .O(gate55inter8));
  nand2 gate618(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate619(.a(s_59), .b(gate55inter3), .O(gate55inter10));
  nor2  gate620(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate621(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate622(.a(gate55inter12), .b(gate55inter1), .O(N320));
xor2 gate56( .a(N288), .b(N289), .O(N321) );

  xor2  gate413(.a(N293), .b(N290), .O(gate57inter0));
  nand2 gate414(.a(gate57inter0), .b(s_30), .O(gate57inter1));
  and2  gate415(.a(N293), .b(N290), .O(gate57inter2));
  inv1  gate416(.a(s_30), .O(gate57inter3));
  inv1  gate417(.a(s_31), .O(gate57inter4));
  nand2 gate418(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate419(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate420(.a(N290), .O(gate57inter7));
  inv1  gate421(.a(N293), .O(gate57inter8));
  nand2 gate422(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate423(.a(s_31), .b(gate57inter3), .O(gate57inter10));
  nor2  gate424(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate425(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate426(.a(gate57inter12), .b(gate57inter1), .O(N338));
xor2 gate58( .a(N296), .b(N299), .O(N339) );
xor2 gate59( .a(N290), .b(N296), .O(N340) );
xor2 gate60( .a(N293), .b(N299), .O(N341) );
xor2 gate61( .a(N302), .b(N305), .O(N342) );

  xor2  gate217(.a(N311), .b(N308), .O(gate62inter0));
  nand2 gate218(.a(gate62inter0), .b(s_2), .O(gate62inter1));
  and2  gate219(.a(N311), .b(N308), .O(gate62inter2));
  inv1  gate220(.a(s_2), .O(gate62inter3));
  inv1  gate221(.a(s_3), .O(gate62inter4));
  nand2 gate222(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate223(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate224(.a(N308), .O(gate62inter7));
  inv1  gate225(.a(N311), .O(gate62inter8));
  nand2 gate226(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate227(.a(s_3), .b(gate62inter3), .O(gate62inter10));
  nor2  gate228(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate229(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate230(.a(gate62inter12), .b(gate62inter1), .O(N343));
xor2 gate63( .a(N302), .b(N308), .O(N344) );
xor2 gate64( .a(N305), .b(N311), .O(N345) );

  xor2  gate427(.a(N342), .b(N266), .O(gate65inter0));
  nand2 gate428(.a(gate65inter0), .b(s_32), .O(gate65inter1));
  and2  gate429(.a(N342), .b(N266), .O(gate65inter2));
  inv1  gate430(.a(s_32), .O(gate65inter3));
  inv1  gate431(.a(s_33), .O(gate65inter4));
  nand2 gate432(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate433(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate434(.a(N266), .O(gate65inter7));
  inv1  gate435(.a(N342), .O(gate65inter8));
  nand2 gate436(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate437(.a(s_33), .b(gate65inter3), .O(gate65inter10));
  nor2  gate438(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate439(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate440(.a(gate65inter12), .b(gate65inter1), .O(N346));
xor2 gate66( .a(N267), .b(N343), .O(N347) );
xor2 gate67( .a(N268), .b(N344), .O(N348) );
xor2 gate68( .a(N269), .b(N345), .O(N349) );
xor2 gate69( .a(N270), .b(N338), .O(N350) );

  xor2  gate595(.a(N339), .b(N271), .O(gate70inter0));
  nand2 gate596(.a(gate70inter0), .b(s_56), .O(gate70inter1));
  and2  gate597(.a(N339), .b(N271), .O(gate70inter2));
  inv1  gate598(.a(s_56), .O(gate70inter3));
  inv1  gate599(.a(s_57), .O(gate70inter4));
  nand2 gate600(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate601(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate602(.a(N271), .O(gate70inter7));
  inv1  gate603(.a(N339), .O(gate70inter8));
  nand2 gate604(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate605(.a(s_57), .b(gate70inter3), .O(gate70inter10));
  nor2  gate606(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate607(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate608(.a(gate70inter12), .b(gate70inter1), .O(N351));
xor2 gate71( .a(N272), .b(N340), .O(N352) );

  xor2  gate287(.a(N341), .b(N273), .O(gate72inter0));
  nand2 gate288(.a(gate72inter0), .b(s_12), .O(gate72inter1));
  and2  gate289(.a(N341), .b(N273), .O(gate72inter2));
  inv1  gate290(.a(s_12), .O(gate72inter3));
  inv1  gate291(.a(s_13), .O(gate72inter4));
  nand2 gate292(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate293(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate294(.a(N273), .O(gate72inter7));
  inv1  gate295(.a(N341), .O(gate72inter8));
  nand2 gate296(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate297(.a(s_13), .b(gate72inter3), .O(gate72inter10));
  nor2  gate298(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate299(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate300(.a(gate72inter12), .b(gate72inter1), .O(N353));

  xor2  gate371(.a(N346), .b(N314), .O(gate73inter0));
  nand2 gate372(.a(gate73inter0), .b(s_24), .O(gate73inter1));
  and2  gate373(.a(N346), .b(N314), .O(gate73inter2));
  inv1  gate374(.a(s_24), .O(gate73inter3));
  inv1  gate375(.a(s_25), .O(gate73inter4));
  nand2 gate376(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate377(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate378(.a(N314), .O(gate73inter7));
  inv1  gate379(.a(N346), .O(gate73inter8));
  nand2 gate380(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate381(.a(s_25), .b(gate73inter3), .O(gate73inter10));
  nor2  gate382(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate383(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate384(.a(gate73inter12), .b(gate73inter1), .O(N354));
xor2 gate74( .a(N315), .b(N347), .O(N367) );

  xor2  gate385(.a(N348), .b(N316), .O(gate75inter0));
  nand2 gate386(.a(gate75inter0), .b(s_26), .O(gate75inter1));
  and2  gate387(.a(N348), .b(N316), .O(gate75inter2));
  inv1  gate388(.a(s_26), .O(gate75inter3));
  inv1  gate389(.a(s_27), .O(gate75inter4));
  nand2 gate390(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate391(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate392(.a(N316), .O(gate75inter7));
  inv1  gate393(.a(N348), .O(gate75inter8));
  nand2 gate394(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate395(.a(s_27), .b(gate75inter3), .O(gate75inter10));
  nor2  gate396(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate397(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate398(.a(gate75inter12), .b(gate75inter1), .O(N380));
xor2 gate76( .a(N317), .b(N349), .O(N393) );
xor2 gate77( .a(N318), .b(N350), .O(N406) );
xor2 gate78( .a(N319), .b(N351), .O(N419) );
xor2 gate79( .a(N320), .b(N352), .O(N432) );

  xor2  gate455(.a(N353), .b(N321), .O(gate80inter0));
  nand2 gate456(.a(gate80inter0), .b(s_36), .O(gate80inter1));
  and2  gate457(.a(N353), .b(N321), .O(gate80inter2));
  inv1  gate458(.a(s_36), .O(gate80inter3));
  inv1  gate459(.a(s_37), .O(gate80inter4));
  nand2 gate460(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate461(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate462(.a(N321), .O(gate80inter7));
  inv1  gate463(.a(N353), .O(gate80inter8));
  nand2 gate464(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate465(.a(s_37), .b(gate80inter3), .O(gate80inter10));
  nor2  gate466(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate467(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate468(.a(gate80inter12), .b(gate80inter1), .O(N445));
inv1 gate81( .a(N354), .O(N554) );
inv1 gate82( .a(N367), .O(N555) );
inv1 gate83( .a(N380), .O(N556) );
inv1 gate84( .a(N354), .O(N557) );
inv1 gate85( .a(N367), .O(N558) );
inv1 gate86( .a(N393), .O(N559) );
inv1 gate87( .a(N354), .O(N560) );
inv1 gate88( .a(N380), .O(N561) );
inv1 gate89( .a(N393), .O(N562) );
inv1 gate90( .a(N367), .O(N563) );
inv1 gate91( .a(N380), .O(N564) );
inv1 gate92( .a(N393), .O(N565) );
inv1 gate93( .a(N419), .O(N566) );
inv1 gate94( .a(N445), .O(N567) );
inv1 gate95( .a(N419), .O(N568) );
inv1 gate96( .a(N432), .O(N569) );
inv1 gate97( .a(N406), .O(N570) );
inv1 gate98( .a(N445), .O(N571) );
inv1 gate99( .a(N406), .O(N572) );
inv1 gate100( .a(N432), .O(N573) );
inv1 gate101( .a(N406), .O(N574) );
inv1 gate102( .a(N419), .O(N575) );
inv1 gate103( .a(N432), .O(N576) );
inv1 gate104( .a(N406), .O(N577) );
inv1 gate105( .a(N419), .O(N578) );
inv1 gate106( .a(N445), .O(N579) );
inv1 gate107( .a(N406), .O(N580) );
inv1 gate108( .a(N432), .O(N581) );
inv1 gate109( .a(N445), .O(N582) );
inv1 gate110( .a(N419), .O(N583) );
inv1 gate111( .a(N432), .O(N584) );
inv1 gate112( .a(N445), .O(N585) );
inv1 gate113( .a(N367), .O(N586) );
inv1 gate114( .a(N393), .O(N587) );
inv1 gate115( .a(N367), .O(N588) );
inv1 gate116( .a(N380), .O(N589) );
inv1 gate117( .a(N354), .O(N590) );
inv1 gate118( .a(N393), .O(N591) );
inv1 gate119( .a(N354), .O(N592) );
inv1 gate120( .a(N380), .O(N593) );
and4 gate121( .a(N554), .b(N555), .c(N556), .d(N393), .O(N594) );
and4 gate122( .a(N557), .b(N558), .c(N380), .d(N559), .O(N595) );
and4 gate123( .a(N560), .b(N367), .c(N561), .d(N562), .O(N596) );
and4 gate124( .a(N354), .b(N563), .c(N564), .d(N565), .O(N597) );
and4 gate125( .a(N574), .b(N575), .c(N576), .d(N445), .O(N598) );
and4 gate126( .a(N577), .b(N578), .c(N432), .d(N579), .O(N599) );
and4 gate127( .a(N580), .b(N419), .c(N581), .d(N582), .O(N600) );
and4 gate128( .a(N406), .b(N583), .c(N584), .d(N585), .O(N601) );
or4 gate129( .a(N594), .b(N595), .c(N596), .d(N597), .O(N602) );
or4 gate130( .a(N598), .b(N599), .c(N600), .d(N601), .O(N607) );
and5 gate131( .a(N406), .b(N566), .c(N432), .d(N567), .e(N602), .O(N620) );
and5 gate132( .a(N406), .b(N568), .c(N569), .d(N445), .e(N602), .O(N625) );
and5 gate133( .a(N570), .b(N419), .c(N432), .d(N571), .e(N602), .O(N630) );
and5 gate134( .a(N572), .b(N419), .c(N573), .d(N445), .e(N602), .O(N635) );
and5 gate135( .a(N354), .b(N586), .c(N380), .d(N587), .e(N607), .O(N640) );
and5 gate136( .a(N354), .b(N588), .c(N589), .d(N393), .e(N607), .O(N645) );
and5 gate137( .a(N590), .b(N367), .c(N380), .d(N591), .e(N607), .O(N650) );
and5 gate138( .a(N592), .b(N367), .c(N593), .d(N393), .e(N607), .O(N655) );
and2 gate139( .a(N354), .b(N620), .O(N692) );
and2 gate140( .a(N367), .b(N620), .O(N693) );
and2 gate141( .a(N380), .b(N620), .O(N694) );
and2 gate142( .a(N393), .b(N620), .O(N695) );
and2 gate143( .a(N354), .b(N625), .O(N696) );
and2 gate144( .a(N367), .b(N625), .O(N697) );
and2 gate145( .a(N380), .b(N625), .O(N698) );
and2 gate146( .a(N393), .b(N625), .O(N699) );
and2 gate147( .a(N354), .b(N630), .O(N700) );
and2 gate148( .a(N367), .b(N630), .O(N701) );
and2 gate149( .a(N380), .b(N630), .O(N702) );
and2 gate150( .a(N393), .b(N630), .O(N703) );
and2 gate151( .a(N354), .b(N635), .O(N704) );
and2 gate152( .a(N367), .b(N635), .O(N705) );
and2 gate153( .a(N380), .b(N635), .O(N706) );
and2 gate154( .a(N393), .b(N635), .O(N707) );
and2 gate155( .a(N406), .b(N640), .O(N708) );
and2 gate156( .a(N419), .b(N640), .O(N709) );
and2 gate157( .a(N432), .b(N640), .O(N710) );
and2 gate158( .a(N445), .b(N640), .O(N711) );
and2 gate159( .a(N406), .b(N645), .O(N712) );
and2 gate160( .a(N419), .b(N645), .O(N713) );
and2 gate161( .a(N432), .b(N645), .O(N714) );
and2 gate162( .a(N445), .b(N645), .O(N715) );
and2 gate163( .a(N406), .b(N650), .O(N716) );
and2 gate164( .a(N419), .b(N650), .O(N717) );
and2 gate165( .a(N432), .b(N650), .O(N718) );
and2 gate166( .a(N445), .b(N650), .O(N719) );
and2 gate167( .a(N406), .b(N655), .O(N720) );
and2 gate168( .a(N419), .b(N655), .O(N721) );
and2 gate169( .a(N432), .b(N655), .O(N722) );
and2 gate170( .a(N445), .b(N655), .O(N723) );
xor2 gate171( .a(N1), .b(N692), .O(N724) );
xor2 gate172( .a(N5), .b(N693), .O(N725) );
xor2 gate173( .a(N9), .b(N694), .O(N726) );
xor2 gate174( .a(N13), .b(N695), .O(N727) );
xor2 gate175( .a(N17), .b(N696), .O(N728) );
xor2 gate176( .a(N21), .b(N697), .O(N729) );
xor2 gate177( .a(N25), .b(N698), .O(N730) );

  xor2  gate623(.a(N699), .b(N29), .O(gate178inter0));
  nand2 gate624(.a(gate178inter0), .b(s_60), .O(gate178inter1));
  and2  gate625(.a(N699), .b(N29), .O(gate178inter2));
  inv1  gate626(.a(s_60), .O(gate178inter3));
  inv1  gate627(.a(s_61), .O(gate178inter4));
  nand2 gate628(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate629(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate630(.a(N29), .O(gate178inter7));
  inv1  gate631(.a(N699), .O(gate178inter8));
  nand2 gate632(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate633(.a(s_61), .b(gate178inter3), .O(gate178inter10));
  nor2  gate634(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate635(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate636(.a(gate178inter12), .b(gate178inter1), .O(N731));
xor2 gate179( .a(N33), .b(N700), .O(N732) );
xor2 gate180( .a(N37), .b(N701), .O(N733) );
xor2 gate181( .a(N41), .b(N702), .O(N734) );
xor2 gate182( .a(N45), .b(N703), .O(N735) );

  xor2  gate511(.a(N704), .b(N49), .O(gate183inter0));
  nand2 gate512(.a(gate183inter0), .b(s_44), .O(gate183inter1));
  and2  gate513(.a(N704), .b(N49), .O(gate183inter2));
  inv1  gate514(.a(s_44), .O(gate183inter3));
  inv1  gate515(.a(s_45), .O(gate183inter4));
  nand2 gate516(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate517(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate518(.a(N49), .O(gate183inter7));
  inv1  gate519(.a(N704), .O(gate183inter8));
  nand2 gate520(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate521(.a(s_45), .b(gate183inter3), .O(gate183inter10));
  nor2  gate522(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate523(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate524(.a(gate183inter12), .b(gate183inter1), .O(N736));
xor2 gate184( .a(N53), .b(N705), .O(N737) );

  xor2  gate441(.a(N706), .b(N57), .O(gate185inter0));
  nand2 gate442(.a(gate185inter0), .b(s_34), .O(gate185inter1));
  and2  gate443(.a(N706), .b(N57), .O(gate185inter2));
  inv1  gate444(.a(s_34), .O(gate185inter3));
  inv1  gate445(.a(s_35), .O(gate185inter4));
  nand2 gate446(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate447(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate448(.a(N57), .O(gate185inter7));
  inv1  gate449(.a(N706), .O(gate185inter8));
  nand2 gate450(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate451(.a(s_35), .b(gate185inter3), .O(gate185inter10));
  nor2  gate452(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate453(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate454(.a(gate185inter12), .b(gate185inter1), .O(N738));
xor2 gate186( .a(N61), .b(N707), .O(N739) );
xor2 gate187( .a(N65), .b(N708), .O(N740) );
xor2 gate188( .a(N69), .b(N709), .O(N741) );

  xor2  gate343(.a(N710), .b(N73), .O(gate189inter0));
  nand2 gate344(.a(gate189inter0), .b(s_20), .O(gate189inter1));
  and2  gate345(.a(N710), .b(N73), .O(gate189inter2));
  inv1  gate346(.a(s_20), .O(gate189inter3));
  inv1  gate347(.a(s_21), .O(gate189inter4));
  nand2 gate348(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate349(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate350(.a(N73), .O(gate189inter7));
  inv1  gate351(.a(N710), .O(gate189inter8));
  nand2 gate352(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate353(.a(s_21), .b(gate189inter3), .O(gate189inter10));
  nor2  gate354(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate355(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate356(.a(gate189inter12), .b(gate189inter1), .O(N742));
xor2 gate190( .a(N77), .b(N711), .O(N743) );

  xor2  gate497(.a(N712), .b(N81), .O(gate191inter0));
  nand2 gate498(.a(gate191inter0), .b(s_42), .O(gate191inter1));
  and2  gate499(.a(N712), .b(N81), .O(gate191inter2));
  inv1  gate500(.a(s_42), .O(gate191inter3));
  inv1  gate501(.a(s_43), .O(gate191inter4));
  nand2 gate502(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate503(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate504(.a(N81), .O(gate191inter7));
  inv1  gate505(.a(N712), .O(gate191inter8));
  nand2 gate506(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate507(.a(s_43), .b(gate191inter3), .O(gate191inter10));
  nor2  gate508(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate509(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate510(.a(gate191inter12), .b(gate191inter1), .O(N744));
xor2 gate192( .a(N85), .b(N713), .O(N745) );

  xor2  gate259(.a(N714), .b(N89), .O(gate193inter0));
  nand2 gate260(.a(gate193inter0), .b(s_8), .O(gate193inter1));
  and2  gate261(.a(N714), .b(N89), .O(gate193inter2));
  inv1  gate262(.a(s_8), .O(gate193inter3));
  inv1  gate263(.a(s_9), .O(gate193inter4));
  nand2 gate264(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate265(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate266(.a(N89), .O(gate193inter7));
  inv1  gate267(.a(N714), .O(gate193inter8));
  nand2 gate268(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate269(.a(s_9), .b(gate193inter3), .O(gate193inter10));
  nor2  gate270(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate271(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate272(.a(gate193inter12), .b(gate193inter1), .O(N746));

  xor2  gate357(.a(N715), .b(N93), .O(gate194inter0));
  nand2 gate358(.a(gate194inter0), .b(s_22), .O(gate194inter1));
  and2  gate359(.a(N715), .b(N93), .O(gate194inter2));
  inv1  gate360(.a(s_22), .O(gate194inter3));
  inv1  gate361(.a(s_23), .O(gate194inter4));
  nand2 gate362(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate363(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate364(.a(N93), .O(gate194inter7));
  inv1  gate365(.a(N715), .O(gate194inter8));
  nand2 gate366(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate367(.a(s_23), .b(gate194inter3), .O(gate194inter10));
  nor2  gate368(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate369(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate370(.a(gate194inter12), .b(gate194inter1), .O(N747));
xor2 gate195( .a(N97), .b(N716), .O(N748) );
xor2 gate196( .a(N101), .b(N717), .O(N749) );

  xor2  gate539(.a(N718), .b(N105), .O(gate197inter0));
  nand2 gate540(.a(gate197inter0), .b(s_48), .O(gate197inter1));
  and2  gate541(.a(N718), .b(N105), .O(gate197inter2));
  inv1  gate542(.a(s_48), .O(gate197inter3));
  inv1  gate543(.a(s_49), .O(gate197inter4));
  nand2 gate544(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate545(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate546(.a(N105), .O(gate197inter7));
  inv1  gate547(.a(N718), .O(gate197inter8));
  nand2 gate548(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate549(.a(s_49), .b(gate197inter3), .O(gate197inter10));
  nor2  gate550(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate551(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate552(.a(gate197inter12), .b(gate197inter1), .O(N750));
xor2 gate198( .a(N109), .b(N719), .O(N751) );
xor2 gate199( .a(N113), .b(N720), .O(N752) );
xor2 gate200( .a(N117), .b(N721), .O(N753) );
xor2 gate201( .a(N121), .b(N722), .O(N754) );
xor2 gate202( .a(N125), .b(N723), .O(N755) );

endmodule