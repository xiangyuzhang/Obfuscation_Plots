module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );

  xor2  gate813(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate814(.a(gate32inter0), .b(s_38), .O(gate32inter1));
  and2  gate815(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate816(.a(s_38), .O(gate32inter3));
  inv1  gate817(.a(s_39), .O(gate32inter4));
  nand2 gate818(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate819(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate820(.a(G12), .O(gate32inter7));
  inv1  gate821(.a(G16), .O(gate32inter8));
  nand2 gate822(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate823(.a(s_39), .b(gate32inter3), .O(gate32inter10));
  nor2  gate824(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate825(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate826(.a(gate32inter12), .b(gate32inter1), .O(G335));
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate1079(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1080(.a(gate36inter0), .b(s_76), .O(gate36inter1));
  and2  gate1081(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1082(.a(s_76), .O(gate36inter3));
  inv1  gate1083(.a(s_77), .O(gate36inter4));
  nand2 gate1084(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1085(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1086(.a(G26), .O(gate36inter7));
  inv1  gate1087(.a(G30), .O(gate36inter8));
  nand2 gate1088(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1089(.a(s_77), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1090(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1091(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1092(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate575(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate576(.a(gate41inter0), .b(s_4), .O(gate41inter1));
  and2  gate577(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate578(.a(s_4), .O(gate41inter3));
  inv1  gate579(.a(s_5), .O(gate41inter4));
  nand2 gate580(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate581(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate582(.a(G1), .O(gate41inter7));
  inv1  gate583(.a(G266), .O(gate41inter8));
  nand2 gate584(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate585(.a(s_5), .b(gate41inter3), .O(gate41inter10));
  nor2  gate586(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate587(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate588(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate1149(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate1150(.a(gate55inter0), .b(s_86), .O(gate55inter1));
  and2  gate1151(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate1152(.a(s_86), .O(gate55inter3));
  inv1  gate1153(.a(s_87), .O(gate55inter4));
  nand2 gate1154(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate1155(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate1156(.a(G15), .O(gate55inter7));
  inv1  gate1157(.a(G287), .O(gate55inter8));
  nand2 gate1158(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate1159(.a(s_87), .b(gate55inter3), .O(gate55inter10));
  nor2  gate1160(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate1161(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate1162(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate1121(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate1122(.a(gate63inter0), .b(s_82), .O(gate63inter1));
  and2  gate1123(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate1124(.a(s_82), .O(gate63inter3));
  inv1  gate1125(.a(s_83), .O(gate63inter4));
  nand2 gate1126(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate1127(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate1128(.a(G23), .O(gate63inter7));
  inv1  gate1129(.a(G299), .O(gate63inter8));
  nand2 gate1130(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate1131(.a(s_83), .b(gate63inter3), .O(gate63inter10));
  nor2  gate1132(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate1133(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate1134(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate561(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate562(.a(gate66inter0), .b(s_2), .O(gate66inter1));
  and2  gate563(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate564(.a(s_2), .O(gate66inter3));
  inv1  gate565(.a(s_3), .O(gate66inter4));
  nand2 gate566(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate567(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate568(.a(G26), .O(gate66inter7));
  inv1  gate569(.a(G302), .O(gate66inter8));
  nand2 gate570(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate571(.a(s_3), .b(gate66inter3), .O(gate66inter10));
  nor2  gate572(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate573(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate574(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate1219(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate1220(.a(gate70inter0), .b(s_96), .O(gate70inter1));
  and2  gate1221(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate1222(.a(s_96), .O(gate70inter3));
  inv1  gate1223(.a(s_97), .O(gate70inter4));
  nand2 gate1224(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate1225(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate1226(.a(G30), .O(gate70inter7));
  inv1  gate1227(.a(G308), .O(gate70inter8));
  nand2 gate1228(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate1229(.a(s_97), .b(gate70inter3), .O(gate70inter10));
  nor2  gate1230(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate1231(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate1232(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate1317(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate1318(.a(gate86inter0), .b(s_110), .O(gate86inter1));
  and2  gate1319(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate1320(.a(s_110), .O(gate86inter3));
  inv1  gate1321(.a(s_111), .O(gate86inter4));
  nand2 gate1322(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate1323(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate1324(.a(G8), .O(gate86inter7));
  inv1  gate1325(.a(G332), .O(gate86inter8));
  nand2 gate1326(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate1327(.a(s_111), .b(gate86inter3), .O(gate86inter10));
  nor2  gate1328(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate1329(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate1330(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate1261(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate1262(.a(gate90inter0), .b(s_102), .O(gate90inter1));
  and2  gate1263(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate1264(.a(s_102), .O(gate90inter3));
  inv1  gate1265(.a(s_103), .O(gate90inter4));
  nand2 gate1266(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate1267(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate1268(.a(G21), .O(gate90inter7));
  inv1  gate1269(.a(G338), .O(gate90inter8));
  nand2 gate1270(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate1271(.a(s_103), .b(gate90inter3), .O(gate90inter10));
  nor2  gate1272(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate1273(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate1274(.a(gate90inter12), .b(gate90inter1), .O(G411));
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );

  xor2  gate1205(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate1206(.a(gate111inter0), .b(s_94), .O(gate111inter1));
  and2  gate1207(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate1208(.a(s_94), .O(gate111inter3));
  inv1  gate1209(.a(s_95), .O(gate111inter4));
  nand2 gate1210(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate1211(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate1212(.a(G374), .O(gate111inter7));
  inv1  gate1213(.a(G375), .O(gate111inter8));
  nand2 gate1214(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate1215(.a(s_95), .b(gate111inter3), .O(gate111inter10));
  nor2  gate1216(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate1217(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate1218(.a(gate111inter12), .b(gate111inter1), .O(G444));
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate1023(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate1024(.a(gate116inter0), .b(s_68), .O(gate116inter1));
  and2  gate1025(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate1026(.a(s_68), .O(gate116inter3));
  inv1  gate1027(.a(s_69), .O(gate116inter4));
  nand2 gate1028(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate1029(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate1030(.a(G384), .O(gate116inter7));
  inv1  gate1031(.a(G385), .O(gate116inter8));
  nand2 gate1032(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate1033(.a(s_69), .b(gate116inter3), .O(gate116inter10));
  nor2  gate1034(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate1035(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate1036(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate589(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate590(.a(gate119inter0), .b(s_6), .O(gate119inter1));
  and2  gate591(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate592(.a(s_6), .O(gate119inter3));
  inv1  gate593(.a(s_7), .O(gate119inter4));
  nand2 gate594(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate595(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate596(.a(G390), .O(gate119inter7));
  inv1  gate597(.a(G391), .O(gate119inter8));
  nand2 gate598(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate599(.a(s_7), .b(gate119inter3), .O(gate119inter10));
  nor2  gate600(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate601(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate602(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate617(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate618(.a(gate126inter0), .b(s_10), .O(gate126inter1));
  and2  gate619(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate620(.a(s_10), .O(gate126inter3));
  inv1  gate621(.a(s_11), .O(gate126inter4));
  nand2 gate622(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate623(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate624(.a(G404), .O(gate126inter7));
  inv1  gate625(.a(G405), .O(gate126inter8));
  nand2 gate626(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate627(.a(s_11), .b(gate126inter3), .O(gate126inter10));
  nor2  gate628(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate629(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate630(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate981(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate982(.a(gate141inter0), .b(s_62), .O(gate141inter1));
  and2  gate983(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate984(.a(s_62), .O(gate141inter3));
  inv1  gate985(.a(s_63), .O(gate141inter4));
  nand2 gate986(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate987(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate988(.a(G450), .O(gate141inter7));
  inv1  gate989(.a(G453), .O(gate141inter8));
  nand2 gate990(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate991(.a(s_63), .b(gate141inter3), .O(gate141inter10));
  nor2  gate992(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate993(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate994(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );

  xor2  gate785(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate786(.a(gate152inter0), .b(s_34), .O(gate152inter1));
  and2  gate787(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate788(.a(s_34), .O(gate152inter3));
  inv1  gate789(.a(s_35), .O(gate152inter4));
  nand2 gate790(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate791(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate792(.a(G516), .O(gate152inter7));
  inv1  gate793(.a(G519), .O(gate152inter8));
  nand2 gate794(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate795(.a(s_35), .b(gate152inter3), .O(gate152inter10));
  nor2  gate796(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate797(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate798(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );

  xor2  gate659(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate660(.a(gate169inter0), .b(s_16), .O(gate169inter1));
  and2  gate661(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate662(.a(s_16), .O(gate169inter3));
  inv1  gate663(.a(s_17), .O(gate169inter4));
  nand2 gate664(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate665(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate666(.a(G474), .O(gate169inter7));
  inv1  gate667(.a(G546), .O(gate169inter8));
  nand2 gate668(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate669(.a(s_17), .b(gate169inter3), .O(gate169inter10));
  nor2  gate670(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate671(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate672(.a(gate169inter12), .b(gate169inter1), .O(G586));
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate869(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate870(.a(gate173inter0), .b(s_46), .O(gate173inter1));
  and2  gate871(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate872(.a(s_46), .O(gate173inter3));
  inv1  gate873(.a(s_47), .O(gate173inter4));
  nand2 gate874(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate875(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate876(.a(G486), .O(gate173inter7));
  inv1  gate877(.a(G552), .O(gate173inter8));
  nand2 gate878(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate879(.a(s_47), .b(gate173inter3), .O(gate173inter10));
  nor2  gate880(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate881(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate882(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate925(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate926(.a(gate175inter0), .b(s_54), .O(gate175inter1));
  and2  gate927(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate928(.a(s_54), .O(gate175inter3));
  inv1  gate929(.a(s_55), .O(gate175inter4));
  nand2 gate930(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate931(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate932(.a(G492), .O(gate175inter7));
  inv1  gate933(.a(G555), .O(gate175inter8));
  nand2 gate934(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate935(.a(s_55), .b(gate175inter3), .O(gate175inter10));
  nor2  gate936(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate937(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate938(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );

  xor2  gate547(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate548(.a(gate182inter0), .b(s_0), .O(gate182inter1));
  and2  gate549(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate550(.a(s_0), .O(gate182inter3));
  inv1  gate551(.a(s_1), .O(gate182inter4));
  nand2 gate552(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate553(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate554(.a(G513), .O(gate182inter7));
  inv1  gate555(.a(G564), .O(gate182inter8));
  nand2 gate556(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate557(.a(s_1), .b(gate182inter3), .O(gate182inter10));
  nor2  gate558(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate559(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate560(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );

  xor2  gate715(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate716(.a(gate202inter0), .b(s_24), .O(gate202inter1));
  and2  gate717(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate718(.a(s_24), .O(gate202inter3));
  inv1  gate719(.a(s_25), .O(gate202inter4));
  nand2 gate720(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate721(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate722(.a(G612), .O(gate202inter7));
  inv1  gate723(.a(G617), .O(gate202inter8));
  nand2 gate724(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate725(.a(s_25), .b(gate202inter3), .O(gate202inter10));
  nor2  gate726(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate727(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate728(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );

  xor2  gate673(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate674(.a(gate208inter0), .b(s_18), .O(gate208inter1));
  and2  gate675(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate676(.a(s_18), .O(gate208inter3));
  inv1  gate677(.a(s_19), .O(gate208inter4));
  nand2 gate678(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate679(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate680(.a(G627), .O(gate208inter7));
  inv1  gate681(.a(G637), .O(gate208inter8));
  nand2 gate682(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate683(.a(s_19), .b(gate208inter3), .O(gate208inter10));
  nor2  gate684(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate685(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate686(.a(gate208inter12), .b(gate208inter1), .O(G687));
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate953(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate954(.a(gate215inter0), .b(s_58), .O(gate215inter1));
  and2  gate955(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate956(.a(s_58), .O(gate215inter3));
  inv1  gate957(.a(s_59), .O(gate215inter4));
  nand2 gate958(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate959(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate960(.a(G607), .O(gate215inter7));
  inv1  gate961(.a(G675), .O(gate215inter8));
  nand2 gate962(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate963(.a(s_59), .b(gate215inter3), .O(gate215inter10));
  nor2  gate964(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate965(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate966(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate1135(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate1136(.a(gate218inter0), .b(s_84), .O(gate218inter1));
  and2  gate1137(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate1138(.a(s_84), .O(gate218inter3));
  inv1  gate1139(.a(s_85), .O(gate218inter4));
  nand2 gate1140(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate1141(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate1142(.a(G627), .O(gate218inter7));
  inv1  gate1143(.a(G678), .O(gate218inter8));
  nand2 gate1144(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate1145(.a(s_85), .b(gate218inter3), .O(gate218inter10));
  nor2  gate1146(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate1147(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate1148(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );

  xor2  gate757(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate758(.a(gate230inter0), .b(s_30), .O(gate230inter1));
  and2  gate759(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate760(.a(s_30), .O(gate230inter3));
  inv1  gate761(.a(s_31), .O(gate230inter4));
  nand2 gate762(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate763(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate764(.a(G700), .O(gate230inter7));
  inv1  gate765(.a(G701), .O(gate230inter8));
  nand2 gate766(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate767(.a(s_31), .b(gate230inter3), .O(gate230inter10));
  nor2  gate768(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate769(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate770(.a(gate230inter12), .b(gate230inter1), .O(G721));
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );

  xor2  gate645(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate646(.a(gate235inter0), .b(s_14), .O(gate235inter1));
  and2  gate647(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate648(.a(s_14), .O(gate235inter3));
  inv1  gate649(.a(s_15), .O(gate235inter4));
  nand2 gate650(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate651(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate652(.a(G248), .O(gate235inter7));
  inv1  gate653(.a(G724), .O(gate235inter8));
  nand2 gate654(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate655(.a(s_15), .b(gate235inter3), .O(gate235inter10));
  nor2  gate656(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate657(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate658(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate1093(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate1094(.a(gate241inter0), .b(s_78), .O(gate241inter1));
  and2  gate1095(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate1096(.a(s_78), .O(gate241inter3));
  inv1  gate1097(.a(s_79), .O(gate241inter4));
  nand2 gate1098(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate1099(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate1100(.a(G242), .O(gate241inter7));
  inv1  gate1101(.a(G730), .O(gate241inter8));
  nand2 gate1102(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate1103(.a(s_79), .b(gate241inter3), .O(gate241inter10));
  nor2  gate1104(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate1105(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate1106(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate1107(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1108(.a(gate243inter0), .b(s_80), .O(gate243inter1));
  and2  gate1109(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1110(.a(s_80), .O(gate243inter3));
  inv1  gate1111(.a(s_81), .O(gate243inter4));
  nand2 gate1112(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1113(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1114(.a(G245), .O(gate243inter7));
  inv1  gate1115(.a(G733), .O(gate243inter8));
  nand2 gate1116(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1117(.a(s_81), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1118(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1119(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1120(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );

  xor2  gate701(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate702(.a(gate246inter0), .b(s_22), .O(gate246inter1));
  and2  gate703(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate704(.a(s_22), .O(gate246inter3));
  inv1  gate705(.a(s_23), .O(gate246inter4));
  nand2 gate706(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate707(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate708(.a(G724), .O(gate246inter7));
  inv1  gate709(.a(G736), .O(gate246inter8));
  nand2 gate710(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate711(.a(s_23), .b(gate246inter3), .O(gate246inter10));
  nor2  gate712(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate713(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate714(.a(gate246inter12), .b(gate246inter1), .O(G759));
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate1163(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate1164(.a(gate252inter0), .b(s_88), .O(gate252inter1));
  and2  gate1165(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate1166(.a(s_88), .O(gate252inter3));
  inv1  gate1167(.a(s_89), .O(gate252inter4));
  nand2 gate1168(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate1169(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate1170(.a(G709), .O(gate252inter7));
  inv1  gate1171(.a(G745), .O(gate252inter8));
  nand2 gate1172(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate1173(.a(s_89), .b(gate252inter3), .O(gate252inter10));
  nor2  gate1174(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate1175(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate1176(.a(gate252inter12), .b(gate252inter1), .O(G765));

  xor2  gate799(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate800(.a(gate253inter0), .b(s_36), .O(gate253inter1));
  and2  gate801(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate802(.a(s_36), .O(gate253inter3));
  inv1  gate803(.a(s_37), .O(gate253inter4));
  nand2 gate804(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate805(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate806(.a(G260), .O(gate253inter7));
  inv1  gate807(.a(G748), .O(gate253inter8));
  nand2 gate808(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate809(.a(s_37), .b(gate253inter3), .O(gate253inter10));
  nor2  gate810(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate811(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate812(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );

  xor2  gate883(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate884(.a(gate259inter0), .b(s_48), .O(gate259inter1));
  and2  gate885(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate886(.a(s_48), .O(gate259inter3));
  inv1  gate887(.a(s_49), .O(gate259inter4));
  nand2 gate888(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate889(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate890(.a(G758), .O(gate259inter7));
  inv1  gate891(.a(G759), .O(gate259inter8));
  nand2 gate892(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate893(.a(s_49), .b(gate259inter3), .O(gate259inter10));
  nor2  gate894(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate895(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate896(.a(gate259inter12), .b(gate259inter1), .O(G776));
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate827(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate828(.a(gate267inter0), .b(s_40), .O(gate267inter1));
  and2  gate829(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate830(.a(s_40), .O(gate267inter3));
  inv1  gate831(.a(s_41), .O(gate267inter4));
  nand2 gate832(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate833(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate834(.a(G648), .O(gate267inter7));
  inv1  gate835(.a(G776), .O(gate267inter8));
  nand2 gate836(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate837(.a(s_41), .b(gate267inter3), .O(gate267inter10));
  nor2  gate838(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate839(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate840(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate1009(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate1010(.a(gate269inter0), .b(s_66), .O(gate269inter1));
  and2  gate1011(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate1012(.a(s_66), .O(gate269inter3));
  inv1  gate1013(.a(s_67), .O(gate269inter4));
  nand2 gate1014(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate1015(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate1016(.a(G654), .O(gate269inter7));
  inv1  gate1017(.a(G782), .O(gate269inter8));
  nand2 gate1018(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate1019(.a(s_67), .b(gate269inter3), .O(gate269inter10));
  nor2  gate1020(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate1021(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate1022(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );

  xor2  gate911(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate912(.a(gate277inter0), .b(s_52), .O(gate277inter1));
  and2  gate913(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate914(.a(s_52), .O(gate277inter3));
  inv1  gate915(.a(s_53), .O(gate277inter4));
  nand2 gate916(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate917(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate918(.a(G648), .O(gate277inter7));
  inv1  gate919(.a(G800), .O(gate277inter8));
  nand2 gate920(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate921(.a(s_53), .b(gate277inter3), .O(gate277inter10));
  nor2  gate922(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate923(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate924(.a(gate277inter12), .b(gate277inter1), .O(G822));

  xor2  gate1233(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate1234(.a(gate278inter0), .b(s_98), .O(gate278inter1));
  and2  gate1235(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate1236(.a(s_98), .O(gate278inter3));
  inv1  gate1237(.a(s_99), .O(gate278inter4));
  nand2 gate1238(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate1239(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate1240(.a(G776), .O(gate278inter7));
  inv1  gate1241(.a(G800), .O(gate278inter8));
  nand2 gate1242(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate1243(.a(s_99), .b(gate278inter3), .O(gate278inter10));
  nor2  gate1244(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate1245(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate1246(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate771(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate772(.a(gate292inter0), .b(s_32), .O(gate292inter1));
  and2  gate773(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate774(.a(s_32), .O(gate292inter3));
  inv1  gate775(.a(s_33), .O(gate292inter4));
  nand2 gate776(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate777(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate778(.a(G824), .O(gate292inter7));
  inv1  gate779(.a(G825), .O(gate292inter8));
  nand2 gate780(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate781(.a(s_33), .b(gate292inter3), .O(gate292inter10));
  nor2  gate782(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate783(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate784(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate855(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate856(.a(gate294inter0), .b(s_44), .O(gate294inter1));
  and2  gate857(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate858(.a(s_44), .O(gate294inter3));
  inv1  gate859(.a(s_45), .O(gate294inter4));
  nand2 gate860(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate861(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate862(.a(G832), .O(gate294inter7));
  inv1  gate863(.a(G833), .O(gate294inter8));
  nand2 gate864(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate865(.a(s_45), .b(gate294inter3), .O(gate294inter10));
  nor2  gate866(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate867(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate868(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate743(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate744(.a(gate388inter0), .b(s_28), .O(gate388inter1));
  and2  gate745(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate746(.a(s_28), .O(gate388inter3));
  inv1  gate747(.a(s_29), .O(gate388inter4));
  nand2 gate748(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate749(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate750(.a(G2), .O(gate388inter7));
  inv1  gate751(.a(G1039), .O(gate388inter8));
  nand2 gate752(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate753(.a(s_29), .b(gate388inter3), .O(gate388inter10));
  nor2  gate754(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate755(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate756(.a(gate388inter12), .b(gate388inter1), .O(G1135));
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate1177(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate1178(.a(gate393inter0), .b(s_90), .O(gate393inter1));
  and2  gate1179(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate1180(.a(s_90), .O(gate393inter3));
  inv1  gate1181(.a(s_91), .O(gate393inter4));
  nand2 gate1182(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate1183(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate1184(.a(G7), .O(gate393inter7));
  inv1  gate1185(.a(G1054), .O(gate393inter8));
  nand2 gate1186(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate1187(.a(s_91), .b(gate393inter3), .O(gate393inter10));
  nor2  gate1188(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate1189(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate1190(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );

  xor2  gate897(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate898(.a(gate404inter0), .b(s_50), .O(gate404inter1));
  and2  gate899(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate900(.a(s_50), .O(gate404inter3));
  inv1  gate901(.a(s_51), .O(gate404inter4));
  nand2 gate902(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate903(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate904(.a(G18), .O(gate404inter7));
  inv1  gate905(.a(G1087), .O(gate404inter8));
  nand2 gate906(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate907(.a(s_51), .b(gate404inter3), .O(gate404inter10));
  nor2  gate908(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate909(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate910(.a(gate404inter12), .b(gate404inter1), .O(G1183));
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate939(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate940(.a(gate409inter0), .b(s_56), .O(gate409inter1));
  and2  gate941(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate942(.a(s_56), .O(gate409inter3));
  inv1  gate943(.a(s_57), .O(gate409inter4));
  nand2 gate944(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate945(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate946(.a(G23), .O(gate409inter7));
  inv1  gate947(.a(G1102), .O(gate409inter8));
  nand2 gate948(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate949(.a(s_57), .b(gate409inter3), .O(gate409inter10));
  nor2  gate950(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate951(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate952(.a(gate409inter12), .b(gate409inter1), .O(G1198));
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );

  xor2  gate687(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate688(.a(gate412inter0), .b(s_20), .O(gate412inter1));
  and2  gate689(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate690(.a(s_20), .O(gate412inter3));
  inv1  gate691(.a(s_21), .O(gate412inter4));
  nand2 gate692(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate693(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate694(.a(G26), .O(gate412inter7));
  inv1  gate695(.a(G1111), .O(gate412inter8));
  nand2 gate696(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate697(.a(s_21), .b(gate412inter3), .O(gate412inter10));
  nor2  gate698(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate699(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate700(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate1065(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate1066(.a(gate428inter0), .b(s_74), .O(gate428inter1));
  and2  gate1067(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate1068(.a(s_74), .O(gate428inter3));
  inv1  gate1069(.a(s_75), .O(gate428inter4));
  nand2 gate1070(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate1071(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate1072(.a(G1048), .O(gate428inter7));
  inv1  gate1073(.a(G1144), .O(gate428inter8));
  nand2 gate1074(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate1075(.a(s_75), .b(gate428inter3), .O(gate428inter10));
  nor2  gate1076(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate1077(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate1078(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate1037(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate1038(.a(gate434inter0), .b(s_70), .O(gate434inter1));
  and2  gate1039(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate1040(.a(s_70), .O(gate434inter3));
  inv1  gate1041(.a(s_71), .O(gate434inter4));
  nand2 gate1042(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate1043(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate1044(.a(G1057), .O(gate434inter7));
  inv1  gate1045(.a(G1153), .O(gate434inter8));
  nand2 gate1046(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate1047(.a(s_71), .b(gate434inter3), .O(gate434inter10));
  nor2  gate1048(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate1049(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate1050(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );

  xor2  gate1289(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate1290(.a(gate447inter0), .b(s_106), .O(gate447inter1));
  and2  gate1291(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate1292(.a(s_106), .O(gate447inter3));
  inv1  gate1293(.a(s_107), .O(gate447inter4));
  nand2 gate1294(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate1295(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate1296(.a(G15), .O(gate447inter7));
  inv1  gate1297(.a(G1174), .O(gate447inter8));
  nand2 gate1298(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate1299(.a(s_107), .b(gate447inter3), .O(gate447inter10));
  nor2  gate1300(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate1301(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate1302(.a(gate447inter12), .b(gate447inter1), .O(G1256));
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );

  xor2  gate1191(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate1192(.a(gate449inter0), .b(s_92), .O(gate449inter1));
  and2  gate1193(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate1194(.a(s_92), .O(gate449inter3));
  inv1  gate1195(.a(s_93), .O(gate449inter4));
  nand2 gate1196(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate1197(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate1198(.a(G16), .O(gate449inter7));
  inv1  gate1199(.a(G1177), .O(gate449inter8));
  nand2 gate1200(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate1201(.a(s_93), .b(gate449inter3), .O(gate449inter10));
  nor2  gate1202(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate1203(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate1204(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate1275(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate1276(.a(gate456inter0), .b(s_104), .O(gate456inter1));
  and2  gate1277(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate1278(.a(s_104), .O(gate456inter3));
  inv1  gate1279(.a(s_105), .O(gate456inter4));
  nand2 gate1280(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate1281(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate1282(.a(G1090), .O(gate456inter7));
  inv1  gate1283(.a(G1186), .O(gate456inter8));
  nand2 gate1284(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate1285(.a(s_105), .b(gate456inter3), .O(gate456inter10));
  nor2  gate1286(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate1287(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate1288(.a(gate456inter12), .b(gate456inter1), .O(G1265));

  xor2  gate1051(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate1052(.a(gate457inter0), .b(s_72), .O(gate457inter1));
  and2  gate1053(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate1054(.a(s_72), .O(gate457inter3));
  inv1  gate1055(.a(s_73), .O(gate457inter4));
  nand2 gate1056(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate1057(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate1058(.a(G20), .O(gate457inter7));
  inv1  gate1059(.a(G1189), .O(gate457inter8));
  nand2 gate1060(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate1061(.a(s_73), .b(gate457inter3), .O(gate457inter10));
  nor2  gate1062(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate1063(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate1064(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate841(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate842(.a(gate461inter0), .b(s_42), .O(gate461inter1));
  and2  gate843(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate844(.a(s_42), .O(gate461inter3));
  inv1  gate845(.a(s_43), .O(gate461inter4));
  nand2 gate846(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate847(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate848(.a(G22), .O(gate461inter7));
  inv1  gate849(.a(G1195), .O(gate461inter8));
  nand2 gate850(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate851(.a(s_43), .b(gate461inter3), .O(gate461inter10));
  nor2  gate852(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate853(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate854(.a(gate461inter12), .b(gate461inter1), .O(G1270));
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate995(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate996(.a(gate474inter0), .b(s_64), .O(gate474inter1));
  and2  gate997(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate998(.a(s_64), .O(gate474inter3));
  inv1  gate999(.a(s_65), .O(gate474inter4));
  nand2 gate1000(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate1001(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate1002(.a(G1117), .O(gate474inter7));
  inv1  gate1003(.a(G1213), .O(gate474inter8));
  nand2 gate1004(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate1005(.a(s_65), .b(gate474inter3), .O(gate474inter10));
  nor2  gate1006(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate1007(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate1008(.a(gate474inter12), .b(gate474inter1), .O(G1283));
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate1303(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate1304(.a(gate476inter0), .b(s_108), .O(gate476inter1));
  and2  gate1305(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate1306(.a(s_108), .O(gate476inter3));
  inv1  gate1307(.a(s_109), .O(gate476inter4));
  nand2 gate1308(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate1309(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate1310(.a(G1120), .O(gate476inter7));
  inv1  gate1311(.a(G1216), .O(gate476inter8));
  nand2 gate1312(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate1313(.a(s_109), .b(gate476inter3), .O(gate476inter10));
  nor2  gate1314(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate1315(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate1316(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );

  xor2  gate729(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate730(.a(gate483inter0), .b(s_26), .O(gate483inter1));
  and2  gate731(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate732(.a(s_26), .O(gate483inter3));
  inv1  gate733(.a(s_27), .O(gate483inter4));
  nand2 gate734(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate735(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate736(.a(G1228), .O(gate483inter7));
  inv1  gate737(.a(G1229), .O(gate483inter8));
  nand2 gate738(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate739(.a(s_27), .b(gate483inter3), .O(gate483inter10));
  nor2  gate740(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate741(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate742(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate603(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate604(.a(gate488inter0), .b(s_8), .O(gate488inter1));
  and2  gate605(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate606(.a(s_8), .O(gate488inter3));
  inv1  gate607(.a(s_9), .O(gate488inter4));
  nand2 gate608(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate609(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate610(.a(G1238), .O(gate488inter7));
  inv1  gate611(.a(G1239), .O(gate488inter8));
  nand2 gate612(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate613(.a(s_9), .b(gate488inter3), .O(gate488inter10));
  nor2  gate614(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate615(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate616(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate631(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate632(.a(gate501inter0), .b(s_12), .O(gate501inter1));
  and2  gate633(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate634(.a(s_12), .O(gate501inter3));
  inv1  gate635(.a(s_13), .O(gate501inter4));
  nand2 gate636(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate637(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate638(.a(G1264), .O(gate501inter7));
  inv1  gate639(.a(G1265), .O(gate501inter8));
  nand2 gate640(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate641(.a(s_13), .b(gate501inter3), .O(gate501inter10));
  nor2  gate642(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate643(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate644(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );

  xor2  gate967(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate968(.a(gate505inter0), .b(s_60), .O(gate505inter1));
  and2  gate969(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate970(.a(s_60), .O(gate505inter3));
  inv1  gate971(.a(s_61), .O(gate505inter4));
  nand2 gate972(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate973(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate974(.a(G1272), .O(gate505inter7));
  inv1  gate975(.a(G1273), .O(gate505inter8));
  nand2 gate976(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate977(.a(s_61), .b(gate505inter3), .O(gate505inter10));
  nor2  gate978(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate979(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate980(.a(gate505inter12), .b(gate505inter1), .O(G1314));
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );

  xor2  gate1247(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate1248(.a(gate512inter0), .b(s_100), .O(gate512inter1));
  and2  gate1249(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate1250(.a(s_100), .O(gate512inter3));
  inv1  gate1251(.a(s_101), .O(gate512inter4));
  nand2 gate1252(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate1253(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate1254(.a(G1286), .O(gate512inter7));
  inv1  gate1255(.a(G1287), .O(gate512inter8));
  nand2 gate1256(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate1257(.a(s_101), .b(gate512inter3), .O(gate512inter10));
  nor2  gate1258(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate1259(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate1260(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule