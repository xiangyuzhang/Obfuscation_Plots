module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281, s_282, s_283, s_284, s_285, s_286, s_287, s_288, s_289, s_290, s_291, s_292, s_293, s_294, s_295, s_296, s_297, s_298, s_299, s_300, s_301, s_302, s_303, s_304, s_305, s_306, s_307, s_308, s_309, s_310, s_311, s_312, s_313, s_314, s_315, s_316, s_317, s_318, s_319, s_320, s_321, s_322, s_323, s_324, s_325, s_326, s_327, s_328, s_329, s_330, s_331, s_332, s_333, s_334, s_335, s_336, s_337, s_338, s_339, s_340, s_341, s_342, s_343, s_344, s_345, s_346, s_347, s_348, s_349, s_350, s_351, s_352, s_353, s_354, s_355, s_356, s_357, s_358, s_359, s_360, s_361, s_362, s_363, s_364, s_365, s_366, s_367, s_368, s_369, s_370, s_371, s_372, s_373, s_374, s_375, s_376, s_377, s_378, s_379, s_380, s_381;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );

  xor2  gate757(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate758(.a(gate10inter0), .b(s_30), .O(gate10inter1));
  and2  gate759(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate760(.a(s_30), .O(gate10inter3));
  inv1  gate761(.a(s_31), .O(gate10inter4));
  nand2 gate762(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate763(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate764(.a(G3), .O(gate10inter7));
  inv1  gate765(.a(G4), .O(gate10inter8));
  nand2 gate766(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate767(.a(s_31), .b(gate10inter3), .O(gate10inter10));
  nor2  gate768(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate769(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate770(.a(gate10inter12), .b(gate10inter1), .O(G269));

  xor2  gate575(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate576(.a(gate11inter0), .b(s_4), .O(gate11inter1));
  and2  gate577(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate578(.a(s_4), .O(gate11inter3));
  inv1  gate579(.a(s_5), .O(gate11inter4));
  nand2 gate580(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate581(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate582(.a(G5), .O(gate11inter7));
  inv1  gate583(.a(G6), .O(gate11inter8));
  nand2 gate584(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate585(.a(s_5), .b(gate11inter3), .O(gate11inter10));
  nor2  gate586(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate587(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate588(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate2325(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate2326(.a(gate13inter0), .b(s_254), .O(gate13inter1));
  and2  gate2327(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate2328(.a(s_254), .O(gate13inter3));
  inv1  gate2329(.a(s_255), .O(gate13inter4));
  nand2 gate2330(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate2331(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate2332(.a(G9), .O(gate13inter7));
  inv1  gate2333(.a(G10), .O(gate13inter8));
  nand2 gate2334(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate2335(.a(s_255), .b(gate13inter3), .O(gate13inter10));
  nor2  gate2336(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate2337(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate2338(.a(gate13inter12), .b(gate13inter1), .O(G278));

  xor2  gate1373(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate1374(.a(gate14inter0), .b(s_118), .O(gate14inter1));
  and2  gate1375(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate1376(.a(s_118), .O(gate14inter3));
  inv1  gate1377(.a(s_119), .O(gate14inter4));
  nand2 gate1378(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate1379(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate1380(.a(G11), .O(gate14inter7));
  inv1  gate1381(.a(G12), .O(gate14inter8));
  nand2 gate1382(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate1383(.a(s_119), .b(gate14inter3), .O(gate14inter10));
  nor2  gate1384(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate1385(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate1386(.a(gate14inter12), .b(gate14inter1), .O(G281));

  xor2  gate2101(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate2102(.a(gate15inter0), .b(s_222), .O(gate15inter1));
  and2  gate2103(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate2104(.a(s_222), .O(gate15inter3));
  inv1  gate2105(.a(s_223), .O(gate15inter4));
  nand2 gate2106(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate2107(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate2108(.a(G13), .O(gate15inter7));
  inv1  gate2109(.a(G14), .O(gate15inter8));
  nand2 gate2110(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate2111(.a(s_223), .b(gate15inter3), .O(gate15inter10));
  nor2  gate2112(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate2113(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate2114(.a(gate15inter12), .b(gate15inter1), .O(G284));

  xor2  gate2339(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate2340(.a(gate16inter0), .b(s_256), .O(gate16inter1));
  and2  gate2341(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate2342(.a(s_256), .O(gate16inter3));
  inv1  gate2343(.a(s_257), .O(gate16inter4));
  nand2 gate2344(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate2345(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate2346(.a(G15), .O(gate16inter7));
  inv1  gate2347(.a(G16), .O(gate16inter8));
  nand2 gate2348(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate2349(.a(s_257), .b(gate16inter3), .O(gate16inter10));
  nor2  gate2350(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate2351(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate2352(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate1751(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate1752(.a(gate19inter0), .b(s_172), .O(gate19inter1));
  and2  gate1753(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate1754(.a(s_172), .O(gate19inter3));
  inv1  gate1755(.a(s_173), .O(gate19inter4));
  nand2 gate1756(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate1757(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate1758(.a(G21), .O(gate19inter7));
  inv1  gate1759(.a(G22), .O(gate19inter8));
  nand2 gate1760(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate1761(.a(s_173), .b(gate19inter3), .O(gate19inter10));
  nor2  gate1762(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate1763(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate1764(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate1835(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate1836(.a(gate23inter0), .b(s_184), .O(gate23inter1));
  and2  gate1837(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate1838(.a(s_184), .O(gate23inter3));
  inv1  gate1839(.a(s_185), .O(gate23inter4));
  nand2 gate1840(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate1841(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate1842(.a(G29), .O(gate23inter7));
  inv1  gate1843(.a(G30), .O(gate23inter8));
  nand2 gate1844(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate1845(.a(s_185), .b(gate23inter3), .O(gate23inter10));
  nor2  gate1846(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate1847(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate1848(.a(gate23inter12), .b(gate23inter1), .O(G308));

  xor2  gate2815(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate2816(.a(gate24inter0), .b(s_324), .O(gate24inter1));
  and2  gate2817(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate2818(.a(s_324), .O(gate24inter3));
  inv1  gate2819(.a(s_325), .O(gate24inter4));
  nand2 gate2820(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate2821(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate2822(.a(G31), .O(gate24inter7));
  inv1  gate2823(.a(G32), .O(gate24inter8));
  nand2 gate2824(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate2825(.a(s_325), .b(gate24inter3), .O(gate24inter10));
  nor2  gate2826(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate2827(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate2828(.a(gate24inter12), .b(gate24inter1), .O(G311));

  xor2  gate1611(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate1612(.a(gate25inter0), .b(s_152), .O(gate25inter1));
  and2  gate1613(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate1614(.a(s_152), .O(gate25inter3));
  inv1  gate1615(.a(s_153), .O(gate25inter4));
  nand2 gate1616(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate1617(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate1618(.a(G1), .O(gate25inter7));
  inv1  gate1619(.a(G5), .O(gate25inter8));
  nand2 gate1620(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate1621(.a(s_153), .b(gate25inter3), .O(gate25inter10));
  nor2  gate1622(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate1623(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate1624(.a(gate25inter12), .b(gate25inter1), .O(G314));

  xor2  gate2521(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate2522(.a(gate26inter0), .b(s_282), .O(gate26inter1));
  and2  gate2523(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate2524(.a(s_282), .O(gate26inter3));
  inv1  gate2525(.a(s_283), .O(gate26inter4));
  nand2 gate2526(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate2527(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate2528(.a(G9), .O(gate26inter7));
  inv1  gate2529(.a(G13), .O(gate26inter8));
  nand2 gate2530(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate2531(.a(s_283), .b(gate26inter3), .O(gate26inter10));
  nor2  gate2532(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate2533(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate2534(.a(gate26inter12), .b(gate26inter1), .O(G317));

  xor2  gate1149(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate1150(.a(gate27inter0), .b(s_86), .O(gate27inter1));
  and2  gate1151(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate1152(.a(s_86), .O(gate27inter3));
  inv1  gate1153(.a(s_87), .O(gate27inter4));
  nand2 gate1154(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate1155(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate1156(.a(G2), .O(gate27inter7));
  inv1  gate1157(.a(G6), .O(gate27inter8));
  nand2 gate1158(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate1159(.a(s_87), .b(gate27inter3), .O(gate27inter10));
  nor2  gate1160(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate1161(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate1162(.a(gate27inter12), .b(gate27inter1), .O(G320));

  xor2  gate1569(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate1570(.a(gate28inter0), .b(s_146), .O(gate28inter1));
  and2  gate1571(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate1572(.a(s_146), .O(gate28inter3));
  inv1  gate1573(.a(s_147), .O(gate28inter4));
  nand2 gate1574(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate1575(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate1576(.a(G10), .O(gate28inter7));
  inv1  gate1577(.a(G14), .O(gate28inter8));
  nand2 gate1578(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate1579(.a(s_147), .b(gate28inter3), .O(gate28inter10));
  nor2  gate1580(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate1581(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate1582(.a(gate28inter12), .b(gate28inter1), .O(G323));
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate855(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate856(.a(gate31inter0), .b(s_44), .O(gate31inter1));
  and2  gate857(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate858(.a(s_44), .O(gate31inter3));
  inv1  gate859(.a(s_45), .O(gate31inter4));
  nand2 gate860(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate861(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate862(.a(G4), .O(gate31inter7));
  inv1  gate863(.a(G8), .O(gate31inter8));
  nand2 gate864(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate865(.a(s_45), .b(gate31inter3), .O(gate31inter10));
  nor2  gate866(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate867(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate868(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate603(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate604(.a(gate37inter0), .b(s_8), .O(gate37inter1));
  and2  gate605(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate606(.a(s_8), .O(gate37inter3));
  inv1  gate607(.a(s_9), .O(gate37inter4));
  nand2 gate608(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate609(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate610(.a(G19), .O(gate37inter7));
  inv1  gate611(.a(G23), .O(gate37inter8));
  nand2 gate612(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate613(.a(s_9), .b(gate37inter3), .O(gate37inter10));
  nor2  gate614(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate615(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate616(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate2689(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate2690(.a(gate39inter0), .b(s_306), .O(gate39inter1));
  and2  gate2691(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate2692(.a(s_306), .O(gate39inter3));
  inv1  gate2693(.a(s_307), .O(gate39inter4));
  nand2 gate2694(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate2695(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate2696(.a(G20), .O(gate39inter7));
  inv1  gate2697(.a(G24), .O(gate39inter8));
  nand2 gate2698(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate2699(.a(s_307), .b(gate39inter3), .O(gate39inter10));
  nor2  gate2700(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate2701(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate2702(.a(gate39inter12), .b(gate39inter1), .O(G356));

  xor2  gate813(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate814(.a(gate40inter0), .b(s_38), .O(gate40inter1));
  and2  gate815(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate816(.a(s_38), .O(gate40inter3));
  inv1  gate817(.a(s_39), .O(gate40inter4));
  nand2 gate818(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate819(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate820(.a(G28), .O(gate40inter7));
  inv1  gate821(.a(G32), .O(gate40inter8));
  nand2 gate822(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate823(.a(s_39), .b(gate40inter3), .O(gate40inter10));
  nor2  gate824(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate825(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate826(.a(gate40inter12), .b(gate40inter1), .O(G359));
nand2 gate41( .a(G1), .b(G266), .O(G362) );

  xor2  gate785(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate786(.a(gate42inter0), .b(s_34), .O(gate42inter1));
  and2  gate787(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate788(.a(s_34), .O(gate42inter3));
  inv1  gate789(.a(s_35), .O(gate42inter4));
  nand2 gate790(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate791(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate792(.a(G2), .O(gate42inter7));
  inv1  gate793(.a(G266), .O(gate42inter8));
  nand2 gate794(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate795(.a(s_35), .b(gate42inter3), .O(gate42inter10));
  nor2  gate796(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate797(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate798(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate3025(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate3026(.a(gate44inter0), .b(s_354), .O(gate44inter1));
  and2  gate3027(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate3028(.a(s_354), .O(gate44inter3));
  inv1  gate3029(.a(s_355), .O(gate44inter4));
  nand2 gate3030(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate3031(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate3032(.a(G4), .O(gate44inter7));
  inv1  gate3033(.a(G269), .O(gate44inter8));
  nand2 gate3034(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate3035(.a(s_355), .b(gate44inter3), .O(gate44inter10));
  nor2  gate3036(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate3037(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate3038(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );

  xor2  gate1513(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate1514(.a(gate47inter0), .b(s_138), .O(gate47inter1));
  and2  gate1515(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate1516(.a(s_138), .O(gate47inter3));
  inv1  gate1517(.a(s_139), .O(gate47inter4));
  nand2 gate1518(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate1519(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate1520(.a(G7), .O(gate47inter7));
  inv1  gate1521(.a(G275), .O(gate47inter8));
  nand2 gate1522(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate1523(.a(s_139), .b(gate47inter3), .O(gate47inter10));
  nor2  gate1524(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate1525(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate1526(.a(gate47inter12), .b(gate47inter1), .O(G368));
nand2 gate48( .a(G8), .b(G275), .O(G369) );

  xor2  gate1695(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate1696(.a(gate49inter0), .b(s_164), .O(gate49inter1));
  and2  gate1697(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate1698(.a(s_164), .O(gate49inter3));
  inv1  gate1699(.a(s_165), .O(gate49inter4));
  nand2 gate1700(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate1701(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate1702(.a(G9), .O(gate49inter7));
  inv1  gate1703(.a(G278), .O(gate49inter8));
  nand2 gate1704(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate1705(.a(s_165), .b(gate49inter3), .O(gate49inter10));
  nor2  gate1706(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate1707(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate1708(.a(gate49inter12), .b(gate49inter1), .O(G370));

  xor2  gate617(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate618(.a(gate50inter0), .b(s_10), .O(gate50inter1));
  and2  gate619(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate620(.a(s_10), .O(gate50inter3));
  inv1  gate621(.a(s_11), .O(gate50inter4));
  nand2 gate622(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate623(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate624(.a(G10), .O(gate50inter7));
  inv1  gate625(.a(G278), .O(gate50inter8));
  nand2 gate626(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate627(.a(s_11), .b(gate50inter3), .O(gate50inter10));
  nor2  gate628(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate629(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate630(.a(gate50inter12), .b(gate50inter1), .O(G371));
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate1219(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate1220(.a(gate52inter0), .b(s_96), .O(gate52inter1));
  and2  gate1221(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate1222(.a(s_96), .O(gate52inter3));
  inv1  gate1223(.a(s_97), .O(gate52inter4));
  nand2 gate1224(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate1225(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate1226(.a(G12), .O(gate52inter7));
  inv1  gate1227(.a(G281), .O(gate52inter8));
  nand2 gate1228(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate1229(.a(s_97), .b(gate52inter3), .O(gate52inter10));
  nor2  gate1230(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate1231(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate1232(.a(gate52inter12), .b(gate52inter1), .O(G373));

  xor2  gate1275(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate1276(.a(gate53inter0), .b(s_104), .O(gate53inter1));
  and2  gate1277(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate1278(.a(s_104), .O(gate53inter3));
  inv1  gate1279(.a(s_105), .O(gate53inter4));
  nand2 gate1280(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate1281(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate1282(.a(G13), .O(gate53inter7));
  inv1  gate1283(.a(G284), .O(gate53inter8));
  nand2 gate1284(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate1285(.a(s_105), .b(gate53inter3), .O(gate53inter10));
  nor2  gate1286(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate1287(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate1288(.a(gate53inter12), .b(gate53inter1), .O(G374));
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate1597(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate1598(.a(gate55inter0), .b(s_150), .O(gate55inter1));
  and2  gate1599(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate1600(.a(s_150), .O(gate55inter3));
  inv1  gate1601(.a(s_151), .O(gate55inter4));
  nand2 gate1602(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate1603(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate1604(.a(G15), .O(gate55inter7));
  inv1  gate1605(.a(G287), .O(gate55inter8));
  nand2 gate1606(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate1607(.a(s_151), .b(gate55inter3), .O(gate55inter10));
  nor2  gate1608(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate1609(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate1610(.a(gate55inter12), .b(gate55inter1), .O(G376));

  xor2  gate645(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate646(.a(gate56inter0), .b(s_14), .O(gate56inter1));
  and2  gate647(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate648(.a(s_14), .O(gate56inter3));
  inv1  gate649(.a(s_15), .O(gate56inter4));
  nand2 gate650(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate651(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate652(.a(G16), .O(gate56inter7));
  inv1  gate653(.a(G287), .O(gate56inter8));
  nand2 gate654(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate655(.a(s_15), .b(gate56inter3), .O(gate56inter10));
  nor2  gate656(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate657(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate658(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );

  xor2  gate1709(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate1710(.a(gate61inter0), .b(s_166), .O(gate61inter1));
  and2  gate1711(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate1712(.a(s_166), .O(gate61inter3));
  inv1  gate1713(.a(s_167), .O(gate61inter4));
  nand2 gate1714(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate1715(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate1716(.a(G21), .O(gate61inter7));
  inv1  gate1717(.a(G296), .O(gate61inter8));
  nand2 gate1718(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate1719(.a(s_167), .b(gate61inter3), .O(gate61inter10));
  nor2  gate1720(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate1721(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate1722(.a(gate61inter12), .b(gate61inter1), .O(G382));
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate897(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate898(.a(gate63inter0), .b(s_50), .O(gate63inter1));
  and2  gate899(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate900(.a(s_50), .O(gate63inter3));
  inv1  gate901(.a(s_51), .O(gate63inter4));
  nand2 gate902(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate903(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate904(.a(G23), .O(gate63inter7));
  inv1  gate905(.a(G299), .O(gate63inter8));
  nand2 gate906(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate907(.a(s_51), .b(gate63inter3), .O(gate63inter10));
  nor2  gate908(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate909(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate910(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate2283(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate2284(.a(gate69inter0), .b(s_248), .O(gate69inter1));
  and2  gate2285(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate2286(.a(s_248), .O(gate69inter3));
  inv1  gate2287(.a(s_249), .O(gate69inter4));
  nand2 gate2288(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate2289(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate2290(.a(G29), .O(gate69inter7));
  inv1  gate2291(.a(G308), .O(gate69inter8));
  nand2 gate2292(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate2293(.a(s_249), .b(gate69inter3), .O(gate69inter10));
  nor2  gate2294(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate2295(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate2296(.a(gate69inter12), .b(gate69inter1), .O(G390));
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate799(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate800(.a(gate74inter0), .b(s_36), .O(gate74inter1));
  and2  gate801(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate802(.a(s_36), .O(gate74inter3));
  inv1  gate803(.a(s_37), .O(gate74inter4));
  nand2 gate804(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate805(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate806(.a(G5), .O(gate74inter7));
  inv1  gate807(.a(G314), .O(gate74inter8));
  nand2 gate808(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate809(.a(s_37), .b(gate74inter3), .O(gate74inter10));
  nor2  gate810(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate811(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate812(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate2759(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate2760(.a(gate77inter0), .b(s_316), .O(gate77inter1));
  and2  gate2761(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate2762(.a(s_316), .O(gate77inter3));
  inv1  gate2763(.a(s_317), .O(gate77inter4));
  nand2 gate2764(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate2765(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate2766(.a(G2), .O(gate77inter7));
  inv1  gate2767(.a(G320), .O(gate77inter8));
  nand2 gate2768(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate2769(.a(s_317), .b(gate77inter3), .O(gate77inter10));
  nor2  gate2770(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate2771(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate2772(.a(gate77inter12), .b(gate77inter1), .O(G398));

  xor2  gate2745(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate2746(.a(gate78inter0), .b(s_314), .O(gate78inter1));
  and2  gate2747(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate2748(.a(s_314), .O(gate78inter3));
  inv1  gate2749(.a(s_315), .O(gate78inter4));
  nand2 gate2750(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate2751(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate2752(.a(G6), .O(gate78inter7));
  inv1  gate2753(.a(G320), .O(gate78inter8));
  nand2 gate2754(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate2755(.a(s_315), .b(gate78inter3), .O(gate78inter10));
  nor2  gate2756(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate2757(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate2758(.a(gate78inter12), .b(gate78inter1), .O(G399));

  xor2  gate2997(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate2998(.a(gate79inter0), .b(s_350), .O(gate79inter1));
  and2  gate2999(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate3000(.a(s_350), .O(gate79inter3));
  inv1  gate3001(.a(s_351), .O(gate79inter4));
  nand2 gate3002(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate3003(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate3004(.a(G10), .O(gate79inter7));
  inv1  gate3005(.a(G323), .O(gate79inter8));
  nand2 gate3006(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate3007(.a(s_351), .b(gate79inter3), .O(gate79inter10));
  nor2  gate3008(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate3009(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate3010(.a(gate79inter12), .b(gate79inter1), .O(G400));
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );

  xor2  gate3207(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate3208(.a(gate83inter0), .b(s_380), .O(gate83inter1));
  and2  gate3209(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate3210(.a(s_380), .O(gate83inter3));
  inv1  gate3211(.a(s_381), .O(gate83inter4));
  nand2 gate3212(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate3213(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate3214(.a(G11), .O(gate83inter7));
  inv1  gate3215(.a(G329), .O(gate83inter8));
  nand2 gate3216(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate3217(.a(s_381), .b(gate83inter3), .O(gate83inter10));
  nor2  gate3218(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate3219(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate3220(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate1947(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate1948(.a(gate86inter0), .b(s_200), .O(gate86inter1));
  and2  gate1949(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate1950(.a(s_200), .O(gate86inter3));
  inv1  gate1951(.a(s_201), .O(gate86inter4));
  nand2 gate1952(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate1953(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate1954(.a(G8), .O(gate86inter7));
  inv1  gate1955(.a(G332), .O(gate86inter8));
  nand2 gate1956(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate1957(.a(s_201), .b(gate86inter3), .O(gate86inter10));
  nor2  gate1958(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate1959(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate1960(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate2227(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate2228(.a(gate88inter0), .b(s_240), .O(gate88inter1));
  and2  gate2229(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate2230(.a(s_240), .O(gate88inter3));
  inv1  gate2231(.a(s_241), .O(gate88inter4));
  nand2 gate2232(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate2233(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate2234(.a(G16), .O(gate88inter7));
  inv1  gate2235(.a(G335), .O(gate88inter8));
  nand2 gate2236(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate2237(.a(s_241), .b(gate88inter3), .O(gate88inter10));
  nor2  gate2238(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate2239(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate2240(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );

  xor2  gate673(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate674(.a(gate92inter0), .b(s_18), .O(gate92inter1));
  and2  gate675(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate676(.a(s_18), .O(gate92inter3));
  inv1  gate677(.a(s_19), .O(gate92inter4));
  nand2 gate678(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate679(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate680(.a(G29), .O(gate92inter7));
  inv1  gate681(.a(G341), .O(gate92inter8));
  nand2 gate682(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate683(.a(s_19), .b(gate92inter3), .O(gate92inter10));
  nor2  gate684(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate685(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate686(.a(gate92inter12), .b(gate92inter1), .O(G413));

  xor2  gate771(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate772(.a(gate93inter0), .b(s_32), .O(gate93inter1));
  and2  gate773(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate774(.a(s_32), .O(gate93inter3));
  inv1  gate775(.a(s_33), .O(gate93inter4));
  nand2 gate776(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate777(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate778(.a(G18), .O(gate93inter7));
  inv1  gate779(.a(G344), .O(gate93inter8));
  nand2 gate780(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate781(.a(s_33), .b(gate93inter3), .O(gate93inter10));
  nor2  gate782(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate783(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate784(.a(gate93inter12), .b(gate93inter1), .O(G414));
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate3151(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate3152(.a(gate95inter0), .b(s_372), .O(gate95inter1));
  and2  gate3153(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate3154(.a(s_372), .O(gate95inter3));
  inv1  gate3155(.a(s_373), .O(gate95inter4));
  nand2 gate3156(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate3157(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate3158(.a(G26), .O(gate95inter7));
  inv1  gate3159(.a(G347), .O(gate95inter8));
  nand2 gate3160(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate3161(.a(s_373), .b(gate95inter3), .O(gate95inter10));
  nor2  gate3162(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate3163(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate3164(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );

  xor2  gate561(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate562(.a(gate97inter0), .b(s_2), .O(gate97inter1));
  and2  gate563(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate564(.a(s_2), .O(gate97inter3));
  inv1  gate565(.a(s_3), .O(gate97inter4));
  nand2 gate566(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate567(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate568(.a(G19), .O(gate97inter7));
  inv1  gate569(.a(G350), .O(gate97inter8));
  nand2 gate570(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate571(.a(s_3), .b(gate97inter3), .O(gate97inter10));
  nor2  gate572(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate573(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate574(.a(gate97inter12), .b(gate97inter1), .O(G418));

  xor2  gate1933(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate1934(.a(gate98inter0), .b(s_198), .O(gate98inter1));
  and2  gate1935(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate1936(.a(s_198), .O(gate98inter3));
  inv1  gate1937(.a(s_199), .O(gate98inter4));
  nand2 gate1938(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1939(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1940(.a(G23), .O(gate98inter7));
  inv1  gate1941(.a(G350), .O(gate98inter8));
  nand2 gate1942(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1943(.a(s_199), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1944(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1945(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1946(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );

  xor2  gate981(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate982(.a(gate103inter0), .b(s_62), .O(gate103inter1));
  and2  gate983(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate984(.a(s_62), .O(gate103inter3));
  inv1  gate985(.a(s_63), .O(gate103inter4));
  nand2 gate986(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate987(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate988(.a(G28), .O(gate103inter7));
  inv1  gate989(.a(G359), .O(gate103inter8));
  nand2 gate990(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate991(.a(s_63), .b(gate103inter3), .O(gate103inter10));
  nor2  gate992(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate993(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate994(.a(gate103inter12), .b(gate103inter1), .O(G424));
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate2017(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate2018(.a(gate106inter0), .b(s_210), .O(gate106inter1));
  and2  gate2019(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate2020(.a(s_210), .O(gate106inter3));
  inv1  gate2021(.a(s_211), .O(gate106inter4));
  nand2 gate2022(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate2023(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate2024(.a(G364), .O(gate106inter7));
  inv1  gate2025(.a(G365), .O(gate106inter8));
  nand2 gate2026(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate2027(.a(s_211), .b(gate106inter3), .O(gate106inter10));
  nor2  gate2028(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate2029(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate2030(.a(gate106inter12), .b(gate106inter1), .O(G429));

  xor2  gate2605(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate2606(.a(gate107inter0), .b(s_294), .O(gate107inter1));
  and2  gate2607(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate2608(.a(s_294), .O(gate107inter3));
  inv1  gate2609(.a(s_295), .O(gate107inter4));
  nand2 gate2610(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate2611(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate2612(.a(G366), .O(gate107inter7));
  inv1  gate2613(.a(G367), .O(gate107inter8));
  nand2 gate2614(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate2615(.a(s_295), .b(gate107inter3), .O(gate107inter10));
  nor2  gate2616(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate2617(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate2618(.a(gate107inter12), .b(gate107inter1), .O(G432));

  xor2  gate1961(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate1962(.a(gate108inter0), .b(s_202), .O(gate108inter1));
  and2  gate1963(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate1964(.a(s_202), .O(gate108inter3));
  inv1  gate1965(.a(s_203), .O(gate108inter4));
  nand2 gate1966(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate1967(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate1968(.a(G368), .O(gate108inter7));
  inv1  gate1969(.a(G369), .O(gate108inter8));
  nand2 gate1970(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate1971(.a(s_203), .b(gate108inter3), .O(gate108inter10));
  nor2  gate1972(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate1973(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate1974(.a(gate108inter12), .b(gate108inter1), .O(G435));

  xor2  gate3067(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate3068(.a(gate109inter0), .b(s_360), .O(gate109inter1));
  and2  gate3069(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate3070(.a(s_360), .O(gate109inter3));
  inv1  gate3071(.a(s_361), .O(gate109inter4));
  nand2 gate3072(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate3073(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate3074(.a(G370), .O(gate109inter7));
  inv1  gate3075(.a(G371), .O(gate109inter8));
  nand2 gate3076(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate3077(.a(s_361), .b(gate109inter3), .O(gate109inter10));
  nor2  gate3078(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate3079(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate3080(.a(gate109inter12), .b(gate109inter1), .O(G438));

  xor2  gate3053(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate3054(.a(gate110inter0), .b(s_358), .O(gate110inter1));
  and2  gate3055(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate3056(.a(s_358), .O(gate110inter3));
  inv1  gate3057(.a(s_359), .O(gate110inter4));
  nand2 gate3058(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate3059(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate3060(.a(G372), .O(gate110inter7));
  inv1  gate3061(.a(G373), .O(gate110inter8));
  nand2 gate3062(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate3063(.a(s_359), .b(gate110inter3), .O(gate110inter10));
  nor2  gate3064(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate3065(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate3066(.a(gate110inter12), .b(gate110inter1), .O(G441));

  xor2  gate1499(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate1500(.a(gate111inter0), .b(s_136), .O(gate111inter1));
  and2  gate1501(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate1502(.a(s_136), .O(gate111inter3));
  inv1  gate1503(.a(s_137), .O(gate111inter4));
  nand2 gate1504(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate1505(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate1506(.a(G374), .O(gate111inter7));
  inv1  gate1507(.a(G375), .O(gate111inter8));
  nand2 gate1508(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate1509(.a(s_137), .b(gate111inter3), .O(gate111inter10));
  nor2  gate1510(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate1511(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate1512(.a(gate111inter12), .b(gate111inter1), .O(G444));

  xor2  gate1765(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate1766(.a(gate112inter0), .b(s_174), .O(gate112inter1));
  and2  gate1767(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate1768(.a(s_174), .O(gate112inter3));
  inv1  gate1769(.a(s_175), .O(gate112inter4));
  nand2 gate1770(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate1771(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate1772(.a(G376), .O(gate112inter7));
  inv1  gate1773(.a(G377), .O(gate112inter8));
  nand2 gate1774(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate1775(.a(s_175), .b(gate112inter3), .O(gate112inter10));
  nor2  gate1776(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate1777(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate1778(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );

  xor2  gate1009(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate1010(.a(gate114inter0), .b(s_66), .O(gate114inter1));
  and2  gate1011(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate1012(.a(s_66), .O(gate114inter3));
  inv1  gate1013(.a(s_67), .O(gate114inter4));
  nand2 gate1014(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate1015(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate1016(.a(G380), .O(gate114inter7));
  inv1  gate1017(.a(G381), .O(gate114inter8));
  nand2 gate1018(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate1019(.a(s_67), .b(gate114inter3), .O(gate114inter10));
  nor2  gate1020(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate1021(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate1022(.a(gate114inter12), .b(gate114inter1), .O(G453));

  xor2  gate1737(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate1738(.a(gate115inter0), .b(s_170), .O(gate115inter1));
  and2  gate1739(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate1740(.a(s_170), .O(gate115inter3));
  inv1  gate1741(.a(s_171), .O(gate115inter4));
  nand2 gate1742(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate1743(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate1744(.a(G382), .O(gate115inter7));
  inv1  gate1745(.a(G383), .O(gate115inter8));
  nand2 gate1746(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate1747(.a(s_171), .b(gate115inter3), .O(gate115inter10));
  nor2  gate1748(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate1749(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate1750(.a(gate115inter12), .b(gate115inter1), .O(G456));

  xor2  gate2941(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate2942(.a(gate116inter0), .b(s_342), .O(gate116inter1));
  and2  gate2943(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate2944(.a(s_342), .O(gate116inter3));
  inv1  gate2945(.a(s_343), .O(gate116inter4));
  nand2 gate2946(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate2947(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate2948(.a(G384), .O(gate116inter7));
  inv1  gate2949(.a(G385), .O(gate116inter8));
  nand2 gate2950(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate2951(.a(s_343), .b(gate116inter3), .O(gate116inter10));
  nor2  gate2952(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate2953(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate2954(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate869(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate870(.a(gate118inter0), .b(s_46), .O(gate118inter1));
  and2  gate871(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate872(.a(s_46), .O(gate118inter3));
  inv1  gate873(.a(s_47), .O(gate118inter4));
  nand2 gate874(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate875(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate876(.a(G388), .O(gate118inter7));
  inv1  gate877(.a(G389), .O(gate118inter8));
  nand2 gate878(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate879(.a(s_47), .b(gate118inter3), .O(gate118inter10));
  nor2  gate880(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate881(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate882(.a(gate118inter12), .b(gate118inter1), .O(G465));
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate2255(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate2256(.a(gate121inter0), .b(s_244), .O(gate121inter1));
  and2  gate2257(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate2258(.a(s_244), .O(gate121inter3));
  inv1  gate2259(.a(s_245), .O(gate121inter4));
  nand2 gate2260(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate2261(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate2262(.a(G394), .O(gate121inter7));
  inv1  gate2263(.a(G395), .O(gate121inter8));
  nand2 gate2264(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate2265(.a(s_245), .b(gate121inter3), .O(gate121inter10));
  nor2  gate2266(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate2267(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate2268(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );

  xor2  gate3165(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate3166(.a(gate127inter0), .b(s_374), .O(gate127inter1));
  and2  gate3167(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate3168(.a(s_374), .O(gate127inter3));
  inv1  gate3169(.a(s_375), .O(gate127inter4));
  nand2 gate3170(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate3171(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate3172(.a(G406), .O(gate127inter7));
  inv1  gate3173(.a(G407), .O(gate127inter8));
  nand2 gate3174(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate3175(.a(s_375), .b(gate127inter3), .O(gate127inter10));
  nor2  gate3176(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate3177(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate3178(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );

  xor2  gate1079(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate1080(.a(gate129inter0), .b(s_76), .O(gate129inter1));
  and2  gate1081(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate1082(.a(s_76), .O(gate129inter3));
  inv1  gate1083(.a(s_77), .O(gate129inter4));
  nand2 gate1084(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate1085(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate1086(.a(G410), .O(gate129inter7));
  inv1  gate1087(.a(G411), .O(gate129inter8));
  nand2 gate1088(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate1089(.a(s_77), .b(gate129inter3), .O(gate129inter10));
  nor2  gate1090(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate1091(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate1092(.a(gate129inter12), .b(gate129inter1), .O(G498));
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate1443(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate1444(.a(gate138inter0), .b(s_128), .O(gate138inter1));
  and2  gate1445(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate1446(.a(s_128), .O(gate138inter3));
  inv1  gate1447(.a(s_129), .O(gate138inter4));
  nand2 gate1448(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate1449(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate1450(.a(G432), .O(gate138inter7));
  inv1  gate1451(.a(G435), .O(gate138inter8));
  nand2 gate1452(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate1453(.a(s_129), .b(gate138inter3), .O(gate138inter10));
  nor2  gate1454(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate1455(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate1456(.a(gate138inter12), .b(gate138inter1), .O(G525));

  xor2  gate1485(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate1486(.a(gate139inter0), .b(s_134), .O(gate139inter1));
  and2  gate1487(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate1488(.a(s_134), .O(gate139inter3));
  inv1  gate1489(.a(s_135), .O(gate139inter4));
  nand2 gate1490(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate1491(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate1492(.a(G438), .O(gate139inter7));
  inv1  gate1493(.a(G441), .O(gate139inter8));
  nand2 gate1494(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate1495(.a(s_135), .b(gate139inter3), .O(gate139inter10));
  nor2  gate1496(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate1497(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate1498(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate2731(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate2732(.a(gate142inter0), .b(s_312), .O(gate142inter1));
  and2  gate2733(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate2734(.a(s_312), .O(gate142inter3));
  inv1  gate2735(.a(s_313), .O(gate142inter4));
  nand2 gate2736(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate2737(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate2738(.a(G456), .O(gate142inter7));
  inv1  gate2739(.a(G459), .O(gate142inter8));
  nand2 gate2740(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate2741(.a(s_313), .b(gate142inter3), .O(gate142inter10));
  nor2  gate2742(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate2743(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate2744(.a(gate142inter12), .b(gate142inter1), .O(G537));
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate2843(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate2844(.a(gate147inter0), .b(s_328), .O(gate147inter1));
  and2  gate2845(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate2846(.a(s_328), .O(gate147inter3));
  inv1  gate2847(.a(s_329), .O(gate147inter4));
  nand2 gate2848(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate2849(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate2850(.a(G486), .O(gate147inter7));
  inv1  gate2851(.a(G489), .O(gate147inter8));
  nand2 gate2852(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate2853(.a(s_329), .b(gate147inter3), .O(gate147inter10));
  nor2  gate2854(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate2855(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate2856(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate1135(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate1136(.a(gate150inter0), .b(s_84), .O(gate150inter1));
  and2  gate1137(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate1138(.a(s_84), .O(gate150inter3));
  inv1  gate1139(.a(s_85), .O(gate150inter4));
  nand2 gate1140(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate1141(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate1142(.a(G504), .O(gate150inter7));
  inv1  gate1143(.a(G507), .O(gate150inter8));
  nand2 gate1144(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate1145(.a(s_85), .b(gate150inter3), .O(gate150inter10));
  nor2  gate1146(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate1147(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate1148(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate1191(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate1192(.a(gate153inter0), .b(s_92), .O(gate153inter1));
  and2  gate1193(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate1194(.a(s_92), .O(gate153inter3));
  inv1  gate1195(.a(s_93), .O(gate153inter4));
  nand2 gate1196(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate1197(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate1198(.a(G426), .O(gate153inter7));
  inv1  gate1199(.a(G522), .O(gate153inter8));
  nand2 gate1200(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate1201(.a(s_93), .b(gate153inter3), .O(gate153inter10));
  nor2  gate1202(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate1203(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate1204(.a(gate153inter12), .b(gate153inter1), .O(G570));
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate1849(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate1850(.a(gate155inter0), .b(s_186), .O(gate155inter1));
  and2  gate1851(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate1852(.a(s_186), .O(gate155inter3));
  inv1  gate1853(.a(s_187), .O(gate155inter4));
  nand2 gate1854(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1855(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1856(.a(G432), .O(gate155inter7));
  inv1  gate1857(.a(G525), .O(gate155inter8));
  nand2 gate1858(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1859(.a(s_187), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1860(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1861(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1862(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate1625(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate1626(.a(gate158inter0), .b(s_154), .O(gate158inter1));
  and2  gate1627(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate1628(.a(s_154), .O(gate158inter3));
  inv1  gate1629(.a(s_155), .O(gate158inter4));
  nand2 gate1630(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate1631(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate1632(.a(G441), .O(gate158inter7));
  inv1  gate1633(.a(G528), .O(gate158inter8));
  nand2 gate1634(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate1635(.a(s_155), .b(gate158inter3), .O(gate158inter10));
  nor2  gate1636(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate1637(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate1638(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate1051(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate1052(.a(gate161inter0), .b(s_72), .O(gate161inter1));
  and2  gate1053(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate1054(.a(s_72), .O(gate161inter3));
  inv1  gate1055(.a(s_73), .O(gate161inter4));
  nand2 gate1056(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate1057(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate1058(.a(G450), .O(gate161inter7));
  inv1  gate1059(.a(G534), .O(gate161inter8));
  nand2 gate1060(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate1061(.a(s_73), .b(gate161inter3), .O(gate161inter10));
  nor2  gate1062(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate1063(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate1064(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate2661(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate2662(.a(gate165inter0), .b(s_302), .O(gate165inter1));
  and2  gate2663(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate2664(.a(s_302), .O(gate165inter3));
  inv1  gate2665(.a(s_303), .O(gate165inter4));
  nand2 gate2666(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate2667(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate2668(.a(G462), .O(gate165inter7));
  inv1  gate2669(.a(G540), .O(gate165inter8));
  nand2 gate2670(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate2671(.a(s_303), .b(gate165inter3), .O(gate165inter10));
  nor2  gate2672(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate2673(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate2674(.a(gate165inter12), .b(gate165inter1), .O(G582));

  xor2  gate2003(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate2004(.a(gate166inter0), .b(s_208), .O(gate166inter1));
  and2  gate2005(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate2006(.a(s_208), .O(gate166inter3));
  inv1  gate2007(.a(s_209), .O(gate166inter4));
  nand2 gate2008(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate2009(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate2010(.a(G465), .O(gate166inter7));
  inv1  gate2011(.a(G540), .O(gate166inter8));
  nand2 gate2012(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate2013(.a(s_209), .b(gate166inter3), .O(gate166inter10));
  nor2  gate2014(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate2015(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate2016(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );

  xor2  gate1527(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate1528(.a(gate168inter0), .b(s_140), .O(gate168inter1));
  and2  gate1529(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate1530(.a(s_140), .O(gate168inter3));
  inv1  gate1531(.a(s_141), .O(gate168inter4));
  nand2 gate1532(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate1533(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate1534(.a(G471), .O(gate168inter7));
  inv1  gate1535(.a(G543), .O(gate168inter8));
  nand2 gate1536(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate1537(.a(s_141), .b(gate168inter3), .O(gate168inter10));
  nor2  gate1538(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate1539(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate1540(.a(gate168inter12), .b(gate168inter1), .O(G585));

  xor2  gate2423(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate2424(.a(gate169inter0), .b(s_268), .O(gate169inter1));
  and2  gate2425(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate2426(.a(s_268), .O(gate169inter3));
  inv1  gate2427(.a(s_269), .O(gate169inter4));
  nand2 gate2428(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate2429(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate2430(.a(G474), .O(gate169inter7));
  inv1  gate2431(.a(G546), .O(gate169inter8));
  nand2 gate2432(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate2433(.a(s_269), .b(gate169inter3), .O(gate169inter10));
  nor2  gate2434(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate2435(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate2436(.a(gate169inter12), .b(gate169inter1), .O(G586));

  xor2  gate2885(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate2886(.a(gate170inter0), .b(s_334), .O(gate170inter1));
  and2  gate2887(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate2888(.a(s_334), .O(gate170inter3));
  inv1  gate2889(.a(s_335), .O(gate170inter4));
  nand2 gate2890(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate2891(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate2892(.a(G477), .O(gate170inter7));
  inv1  gate2893(.a(G546), .O(gate170inter8));
  nand2 gate2894(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate2895(.a(s_335), .b(gate170inter3), .O(gate170inter10));
  nor2  gate2896(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate2897(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate2898(.a(gate170inter12), .b(gate170inter1), .O(G587));

  xor2  gate1555(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate1556(.a(gate171inter0), .b(s_144), .O(gate171inter1));
  and2  gate1557(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate1558(.a(s_144), .O(gate171inter3));
  inv1  gate1559(.a(s_145), .O(gate171inter4));
  nand2 gate1560(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate1561(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate1562(.a(G480), .O(gate171inter7));
  inv1  gate1563(.a(G549), .O(gate171inter8));
  nand2 gate1564(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate1565(.a(s_145), .b(gate171inter3), .O(gate171inter10));
  nor2  gate1566(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate1567(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate1568(.a(gate171inter12), .b(gate171inter1), .O(G588));

  xor2  gate1471(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate1472(.a(gate172inter0), .b(s_132), .O(gate172inter1));
  and2  gate1473(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate1474(.a(s_132), .O(gate172inter3));
  inv1  gate1475(.a(s_133), .O(gate172inter4));
  nand2 gate1476(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate1477(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate1478(.a(G483), .O(gate172inter7));
  inv1  gate1479(.a(G549), .O(gate172inter8));
  nand2 gate1480(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate1481(.a(s_133), .b(gate172inter3), .O(gate172inter10));
  nor2  gate1482(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate1483(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate1484(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );

  xor2  gate2507(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate2508(.a(gate176inter0), .b(s_280), .O(gate176inter1));
  and2  gate2509(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate2510(.a(s_280), .O(gate176inter3));
  inv1  gate2511(.a(s_281), .O(gate176inter4));
  nand2 gate2512(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate2513(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate2514(.a(G495), .O(gate176inter7));
  inv1  gate2515(.a(G555), .O(gate176inter8));
  nand2 gate2516(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate2517(.a(s_281), .b(gate176inter3), .O(gate176inter10));
  nor2  gate2518(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate2519(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate2520(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );

  xor2  gate1359(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate1360(.a(gate179inter0), .b(s_116), .O(gate179inter1));
  and2  gate1361(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate1362(.a(s_116), .O(gate179inter3));
  inv1  gate1363(.a(s_117), .O(gate179inter4));
  nand2 gate1364(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate1365(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate1366(.a(G504), .O(gate179inter7));
  inv1  gate1367(.a(G561), .O(gate179inter8));
  nand2 gate1368(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate1369(.a(s_117), .b(gate179inter3), .O(gate179inter10));
  nor2  gate1370(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate1371(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate1372(.a(gate179inter12), .b(gate179inter1), .O(G596));

  xor2  gate2409(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate2410(.a(gate180inter0), .b(s_266), .O(gate180inter1));
  and2  gate2411(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate2412(.a(s_266), .O(gate180inter3));
  inv1  gate2413(.a(s_267), .O(gate180inter4));
  nand2 gate2414(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate2415(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate2416(.a(G507), .O(gate180inter7));
  inv1  gate2417(.a(G561), .O(gate180inter8));
  nand2 gate2418(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate2419(.a(s_267), .b(gate180inter3), .O(gate180inter10));
  nor2  gate2420(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate2421(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate2422(.a(gate180inter12), .b(gate180inter1), .O(G597));
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate547(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate548(.a(gate183inter0), .b(s_0), .O(gate183inter1));
  and2  gate549(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate550(.a(s_0), .O(gate183inter3));
  inv1  gate551(.a(s_1), .O(gate183inter4));
  nand2 gate552(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate553(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate554(.a(G516), .O(gate183inter7));
  inv1  gate555(.a(G567), .O(gate183inter8));
  nand2 gate556(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate557(.a(s_1), .b(gate183inter3), .O(gate183inter10));
  nor2  gate558(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate559(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate560(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate2269(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate2270(.a(gate187inter0), .b(s_246), .O(gate187inter1));
  and2  gate2271(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate2272(.a(s_246), .O(gate187inter3));
  inv1  gate2273(.a(s_247), .O(gate187inter4));
  nand2 gate2274(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate2275(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate2276(.a(G574), .O(gate187inter7));
  inv1  gate2277(.a(G575), .O(gate187inter8));
  nand2 gate2278(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate2279(.a(s_247), .b(gate187inter3), .O(gate187inter10));
  nor2  gate2280(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate2281(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate2282(.a(gate187inter12), .b(gate187inter1), .O(G612));
nand2 gate188( .a(G576), .b(G577), .O(G617) );

  xor2  gate1317(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate1318(.a(gate189inter0), .b(s_110), .O(gate189inter1));
  and2  gate1319(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate1320(.a(s_110), .O(gate189inter3));
  inv1  gate1321(.a(s_111), .O(gate189inter4));
  nand2 gate1322(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate1323(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate1324(.a(G578), .O(gate189inter7));
  inv1  gate1325(.a(G579), .O(gate189inter8));
  nand2 gate1326(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate1327(.a(s_111), .b(gate189inter3), .O(gate189inter10));
  nor2  gate1328(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate1329(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate1330(.a(gate189inter12), .b(gate189inter1), .O(G622));
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate1863(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate1864(.a(gate193inter0), .b(s_188), .O(gate193inter1));
  and2  gate1865(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate1866(.a(s_188), .O(gate193inter3));
  inv1  gate1867(.a(s_189), .O(gate193inter4));
  nand2 gate1868(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate1869(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate1870(.a(G586), .O(gate193inter7));
  inv1  gate1871(.a(G587), .O(gate193inter8));
  nand2 gate1872(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate1873(.a(s_189), .b(gate193inter3), .O(gate193inter10));
  nor2  gate1874(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate1875(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate1876(.a(gate193inter12), .b(gate193inter1), .O(G642));

  xor2  gate2913(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate2914(.a(gate194inter0), .b(s_338), .O(gate194inter1));
  and2  gate2915(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate2916(.a(s_338), .O(gate194inter3));
  inv1  gate2917(.a(s_339), .O(gate194inter4));
  nand2 gate2918(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate2919(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate2920(.a(G588), .O(gate194inter7));
  inv1  gate2921(.a(G589), .O(gate194inter8));
  nand2 gate2922(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate2923(.a(s_339), .b(gate194inter3), .O(gate194inter10));
  nor2  gate2924(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate2925(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate2926(.a(gate194inter12), .b(gate194inter1), .O(G645));

  xor2  gate1261(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate1262(.a(gate195inter0), .b(s_102), .O(gate195inter1));
  and2  gate1263(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate1264(.a(s_102), .O(gate195inter3));
  inv1  gate1265(.a(s_103), .O(gate195inter4));
  nand2 gate1266(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate1267(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate1268(.a(G590), .O(gate195inter7));
  inv1  gate1269(.a(G591), .O(gate195inter8));
  nand2 gate1270(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate1271(.a(s_103), .b(gate195inter3), .O(gate195inter10));
  nor2  gate1272(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate1273(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate1274(.a(gate195inter12), .b(gate195inter1), .O(G648));

  xor2  gate3179(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate3180(.a(gate196inter0), .b(s_376), .O(gate196inter1));
  and2  gate3181(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate3182(.a(s_376), .O(gate196inter3));
  inv1  gate3183(.a(s_377), .O(gate196inter4));
  nand2 gate3184(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate3185(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate3186(.a(G592), .O(gate196inter7));
  inv1  gate3187(.a(G593), .O(gate196inter8));
  nand2 gate3188(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate3189(.a(s_377), .b(gate196inter3), .O(gate196inter10));
  nor2  gate3190(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate3191(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate3192(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );

  xor2  gate2969(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate2970(.a(gate199inter0), .b(s_346), .O(gate199inter1));
  and2  gate2971(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate2972(.a(s_346), .O(gate199inter3));
  inv1  gate2973(.a(s_347), .O(gate199inter4));
  nand2 gate2974(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate2975(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate2976(.a(G598), .O(gate199inter7));
  inv1  gate2977(.a(G599), .O(gate199inter8));
  nand2 gate2978(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate2979(.a(s_347), .b(gate199inter3), .O(gate199inter10));
  nor2  gate2980(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate2981(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate2982(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate967(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate968(.a(gate201inter0), .b(s_60), .O(gate201inter1));
  and2  gate969(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate970(.a(s_60), .O(gate201inter3));
  inv1  gate971(.a(s_61), .O(gate201inter4));
  nand2 gate972(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate973(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate974(.a(G602), .O(gate201inter7));
  inv1  gate975(.a(G607), .O(gate201inter8));
  nand2 gate976(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate977(.a(s_61), .b(gate201inter3), .O(gate201inter10));
  nor2  gate978(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate979(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate980(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );

  xor2  gate1681(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate1682(.a(gate204inter0), .b(s_162), .O(gate204inter1));
  and2  gate1683(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate1684(.a(s_162), .O(gate204inter3));
  inv1  gate1685(.a(s_163), .O(gate204inter4));
  nand2 gate1686(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate1687(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate1688(.a(G607), .O(gate204inter7));
  inv1  gate1689(.a(G617), .O(gate204inter8));
  nand2 gate1690(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate1691(.a(s_163), .b(gate204inter3), .O(gate204inter10));
  nor2  gate1692(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate1693(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate1694(.a(gate204inter12), .b(gate204inter1), .O(G675));
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate1793(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate1794(.a(gate206inter0), .b(s_178), .O(gate206inter1));
  and2  gate1795(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate1796(.a(s_178), .O(gate206inter3));
  inv1  gate1797(.a(s_179), .O(gate206inter4));
  nand2 gate1798(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate1799(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate1800(.a(G632), .O(gate206inter7));
  inv1  gate1801(.a(G637), .O(gate206inter8));
  nand2 gate1802(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate1803(.a(s_179), .b(gate206inter3), .O(gate206inter10));
  nor2  gate1804(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate1805(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate1806(.a(gate206inter12), .b(gate206inter1), .O(G681));

  xor2  gate2577(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate2578(.a(gate207inter0), .b(s_290), .O(gate207inter1));
  and2  gate2579(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate2580(.a(s_290), .O(gate207inter3));
  inv1  gate2581(.a(s_291), .O(gate207inter4));
  nand2 gate2582(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate2583(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate2584(.a(G622), .O(gate207inter7));
  inv1  gate2585(.a(G632), .O(gate207inter8));
  nand2 gate2586(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate2587(.a(s_291), .b(gate207inter3), .O(gate207inter10));
  nor2  gate2588(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate2589(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate2590(.a(gate207inter12), .b(gate207inter1), .O(G684));

  xor2  gate925(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate926(.a(gate208inter0), .b(s_54), .O(gate208inter1));
  and2  gate927(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate928(.a(s_54), .O(gate208inter3));
  inv1  gate929(.a(s_55), .O(gate208inter4));
  nand2 gate930(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate931(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate932(.a(G627), .O(gate208inter7));
  inv1  gate933(.a(G637), .O(gate208inter8));
  nand2 gate934(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate935(.a(s_55), .b(gate208inter3), .O(gate208inter10));
  nor2  gate936(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate937(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate938(.a(gate208inter12), .b(gate208inter1), .O(G687));
nand2 gate209( .a(G602), .b(G666), .O(G690) );

  xor2  gate1289(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate1290(.a(gate210inter0), .b(s_106), .O(gate210inter1));
  and2  gate1291(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate1292(.a(s_106), .O(gate210inter3));
  inv1  gate1293(.a(s_107), .O(gate210inter4));
  nand2 gate1294(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate1295(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate1296(.a(G607), .O(gate210inter7));
  inv1  gate1297(.a(G666), .O(gate210inter8));
  nand2 gate1298(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate1299(.a(s_107), .b(gate210inter3), .O(gate210inter10));
  nor2  gate1300(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate1301(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate1302(.a(gate210inter12), .b(gate210inter1), .O(G691));

  xor2  gate2633(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate2634(.a(gate211inter0), .b(s_298), .O(gate211inter1));
  and2  gate2635(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate2636(.a(s_298), .O(gate211inter3));
  inv1  gate2637(.a(s_299), .O(gate211inter4));
  nand2 gate2638(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate2639(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate2640(.a(G612), .O(gate211inter7));
  inv1  gate2641(.a(G669), .O(gate211inter8));
  nand2 gate2642(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate2643(.a(s_299), .b(gate211inter3), .O(gate211inter10));
  nor2  gate2644(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate2645(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate2646(.a(gate211inter12), .b(gate211inter1), .O(G692));

  xor2  gate1093(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate1094(.a(gate212inter0), .b(s_78), .O(gate212inter1));
  and2  gate1095(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate1096(.a(s_78), .O(gate212inter3));
  inv1  gate1097(.a(s_79), .O(gate212inter4));
  nand2 gate1098(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate1099(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate1100(.a(G617), .O(gate212inter7));
  inv1  gate1101(.a(G669), .O(gate212inter8));
  nand2 gate1102(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate1103(.a(s_79), .b(gate212inter3), .O(gate212inter10));
  nor2  gate1104(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate1105(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate1106(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate953(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate954(.a(gate214inter0), .b(s_58), .O(gate214inter1));
  and2  gate955(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate956(.a(s_58), .O(gate214inter3));
  inv1  gate957(.a(s_59), .O(gate214inter4));
  nand2 gate958(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate959(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate960(.a(G612), .O(gate214inter7));
  inv1  gate961(.a(G672), .O(gate214inter8));
  nand2 gate962(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate963(.a(s_59), .b(gate214inter3), .O(gate214inter10));
  nor2  gate964(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate965(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate966(.a(gate214inter12), .b(gate214inter1), .O(G695));

  xor2  gate2563(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate2564(.a(gate215inter0), .b(s_288), .O(gate215inter1));
  and2  gate2565(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate2566(.a(s_288), .O(gate215inter3));
  inv1  gate2567(.a(s_289), .O(gate215inter4));
  nand2 gate2568(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate2569(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate2570(.a(G607), .O(gate215inter7));
  inv1  gate2571(.a(G675), .O(gate215inter8));
  nand2 gate2572(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate2573(.a(s_289), .b(gate215inter3), .O(gate215inter10));
  nor2  gate2574(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate2575(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate2576(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );

  xor2  gate1303(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate1304(.a(gate217inter0), .b(s_108), .O(gate217inter1));
  and2  gate1305(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate1306(.a(s_108), .O(gate217inter3));
  inv1  gate1307(.a(s_109), .O(gate217inter4));
  nand2 gate1308(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate1309(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate1310(.a(G622), .O(gate217inter7));
  inv1  gate1311(.a(G678), .O(gate217inter8));
  nand2 gate1312(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate1313(.a(s_109), .b(gate217inter3), .O(gate217inter10));
  nor2  gate1314(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate1315(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate1316(.a(gate217inter12), .b(gate217inter1), .O(G698));
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate1163(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate1164(.a(gate220inter0), .b(s_88), .O(gate220inter1));
  and2  gate1165(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate1166(.a(s_88), .O(gate220inter3));
  inv1  gate1167(.a(s_89), .O(gate220inter4));
  nand2 gate1168(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate1169(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate1170(.a(G637), .O(gate220inter7));
  inv1  gate1171(.a(G681), .O(gate220inter8));
  nand2 gate1172(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate1173(.a(s_89), .b(gate220inter3), .O(gate220inter10));
  nor2  gate1174(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate1175(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate1176(.a(gate220inter12), .b(gate220inter1), .O(G701));
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate2171(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate2172(.a(gate224inter0), .b(s_232), .O(gate224inter1));
  and2  gate2173(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate2174(.a(s_232), .O(gate224inter3));
  inv1  gate2175(.a(s_233), .O(gate224inter4));
  nand2 gate2176(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate2177(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate2178(.a(G637), .O(gate224inter7));
  inv1  gate2179(.a(G687), .O(gate224inter8));
  nand2 gate2180(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate2181(.a(s_233), .b(gate224inter3), .O(gate224inter10));
  nor2  gate2182(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate2183(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate2184(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate1429(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate1430(.a(gate227inter0), .b(s_126), .O(gate227inter1));
  and2  gate1431(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate1432(.a(s_126), .O(gate227inter3));
  inv1  gate1433(.a(s_127), .O(gate227inter4));
  nand2 gate1434(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate1435(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate1436(.a(G694), .O(gate227inter7));
  inv1  gate1437(.a(G695), .O(gate227inter8));
  nand2 gate1438(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate1439(.a(s_127), .b(gate227inter3), .O(gate227inter10));
  nor2  gate1440(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate1441(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate1442(.a(gate227inter12), .b(gate227inter1), .O(G712));
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );

  xor2  gate1247(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate1248(.a(gate230inter0), .b(s_100), .O(gate230inter1));
  and2  gate1249(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate1250(.a(s_100), .O(gate230inter3));
  inv1  gate1251(.a(s_101), .O(gate230inter4));
  nand2 gate1252(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate1253(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate1254(.a(G700), .O(gate230inter7));
  inv1  gate1255(.a(G701), .O(gate230inter8));
  nand2 gate1256(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate1257(.a(s_101), .b(gate230inter3), .O(gate230inter10));
  nor2  gate1258(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate1259(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate1260(.a(gate230inter12), .b(gate230inter1), .O(G721));

  xor2  gate1457(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate1458(.a(gate231inter0), .b(s_130), .O(gate231inter1));
  and2  gate1459(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate1460(.a(s_130), .O(gate231inter3));
  inv1  gate1461(.a(s_131), .O(gate231inter4));
  nand2 gate1462(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate1463(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate1464(.a(G702), .O(gate231inter7));
  inv1  gate1465(.a(G703), .O(gate231inter8));
  nand2 gate1466(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate1467(.a(s_131), .b(gate231inter3), .O(gate231inter10));
  nor2  gate1468(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate1469(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate1470(.a(gate231inter12), .b(gate231inter1), .O(G724));

  xor2  gate1107(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate1108(.a(gate232inter0), .b(s_80), .O(gate232inter1));
  and2  gate1109(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate1110(.a(s_80), .O(gate232inter3));
  inv1  gate1111(.a(s_81), .O(gate232inter4));
  nand2 gate1112(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate1113(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate1114(.a(G704), .O(gate232inter7));
  inv1  gate1115(.a(G705), .O(gate232inter8));
  nand2 gate1116(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate1117(.a(s_81), .b(gate232inter3), .O(gate232inter10));
  nor2  gate1118(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate1119(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate1120(.a(gate232inter12), .b(gate232inter1), .O(G727));

  xor2  gate2395(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate2396(.a(gate233inter0), .b(s_264), .O(gate233inter1));
  and2  gate2397(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate2398(.a(s_264), .O(gate233inter3));
  inv1  gate2399(.a(s_265), .O(gate233inter4));
  nand2 gate2400(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate2401(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate2402(.a(G242), .O(gate233inter7));
  inv1  gate2403(.a(G718), .O(gate233inter8));
  nand2 gate2404(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate2405(.a(s_265), .b(gate233inter3), .O(gate233inter10));
  nor2  gate2406(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate2407(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate2408(.a(gate233inter12), .b(gate233inter1), .O(G730));

  xor2  gate2451(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate2452(.a(gate234inter0), .b(s_272), .O(gate234inter1));
  and2  gate2453(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate2454(.a(s_272), .O(gate234inter3));
  inv1  gate2455(.a(s_273), .O(gate234inter4));
  nand2 gate2456(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate2457(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate2458(.a(G245), .O(gate234inter7));
  inv1  gate2459(.a(G721), .O(gate234inter8));
  nand2 gate2460(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate2461(.a(s_273), .b(gate234inter3), .O(gate234inter10));
  nor2  gate2462(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate2463(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate2464(.a(gate234inter12), .b(gate234inter1), .O(G733));

  xor2  gate2927(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate2928(.a(gate235inter0), .b(s_340), .O(gate235inter1));
  and2  gate2929(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate2930(.a(s_340), .O(gate235inter3));
  inv1  gate2931(.a(s_341), .O(gate235inter4));
  nand2 gate2932(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate2933(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate2934(.a(G248), .O(gate235inter7));
  inv1  gate2935(.a(G724), .O(gate235inter8));
  nand2 gate2936(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate2937(.a(s_341), .b(gate235inter3), .O(gate235inter10));
  nor2  gate2938(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate2939(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate2940(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate631(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate632(.a(gate237inter0), .b(s_12), .O(gate237inter1));
  and2  gate633(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate634(.a(s_12), .O(gate237inter3));
  inv1  gate635(.a(s_13), .O(gate237inter4));
  nand2 gate636(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate637(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate638(.a(G254), .O(gate237inter7));
  inv1  gate639(.a(G706), .O(gate237inter8));
  nand2 gate640(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate641(.a(s_13), .b(gate237inter3), .O(gate237inter10));
  nor2  gate642(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate643(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate644(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate1037(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate1038(.a(gate241inter0), .b(s_70), .O(gate241inter1));
  and2  gate1039(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate1040(.a(s_70), .O(gate241inter3));
  inv1  gate1041(.a(s_71), .O(gate241inter4));
  nand2 gate1042(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate1043(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate1044(.a(G242), .O(gate241inter7));
  inv1  gate1045(.a(G730), .O(gate241inter8));
  nand2 gate1046(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate1047(.a(s_71), .b(gate241inter3), .O(gate241inter10));
  nor2  gate1048(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate1049(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate1050(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate659(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate660(.a(gate245inter0), .b(s_16), .O(gate245inter1));
  and2  gate661(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate662(.a(s_16), .O(gate245inter3));
  inv1  gate663(.a(s_17), .O(gate245inter4));
  nand2 gate664(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate665(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate666(.a(G248), .O(gate245inter7));
  inv1  gate667(.a(G736), .O(gate245inter8));
  nand2 gate668(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate669(.a(s_17), .b(gate245inter3), .O(gate245inter10));
  nor2  gate670(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate671(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate672(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate1401(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate1402(.a(gate248inter0), .b(s_122), .O(gate248inter1));
  and2  gate1403(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate1404(.a(s_122), .O(gate248inter3));
  inv1  gate1405(.a(s_123), .O(gate248inter4));
  nand2 gate1406(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate1407(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate1408(.a(G727), .O(gate248inter7));
  inv1  gate1409(.a(G739), .O(gate248inter8));
  nand2 gate1410(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate1411(.a(s_123), .b(gate248inter3), .O(gate248inter10));
  nor2  gate1412(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate1413(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate1414(.a(gate248inter12), .b(gate248inter1), .O(G761));

  xor2  gate589(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate590(.a(gate249inter0), .b(s_6), .O(gate249inter1));
  and2  gate591(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate592(.a(s_6), .O(gate249inter3));
  inv1  gate593(.a(s_7), .O(gate249inter4));
  nand2 gate594(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate595(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate596(.a(G254), .O(gate249inter7));
  inv1  gate597(.a(G742), .O(gate249inter8));
  nand2 gate598(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate599(.a(s_7), .b(gate249inter3), .O(gate249inter10));
  nor2  gate600(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate601(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate602(.a(gate249inter12), .b(gate249inter1), .O(G762));

  xor2  gate2157(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate2158(.a(gate250inter0), .b(s_230), .O(gate250inter1));
  and2  gate2159(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate2160(.a(s_230), .O(gate250inter3));
  inv1  gate2161(.a(s_231), .O(gate250inter4));
  nand2 gate2162(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate2163(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate2164(.a(G706), .O(gate250inter7));
  inv1  gate2165(.a(G742), .O(gate250inter8));
  nand2 gate2166(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate2167(.a(s_231), .b(gate250inter3), .O(gate250inter10));
  nor2  gate2168(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate2169(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate2170(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate1667(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate1668(.a(gate253inter0), .b(s_160), .O(gate253inter1));
  and2  gate1669(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate1670(.a(s_160), .O(gate253inter3));
  inv1  gate1671(.a(s_161), .O(gate253inter4));
  nand2 gate1672(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate1673(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate1674(.a(G260), .O(gate253inter7));
  inv1  gate1675(.a(G748), .O(gate253inter8));
  nand2 gate1676(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate1677(.a(s_161), .b(gate253inter3), .O(gate253inter10));
  nor2  gate1678(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate1679(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate1680(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate1177(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate1178(.a(gate257inter0), .b(s_90), .O(gate257inter1));
  and2  gate1179(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate1180(.a(s_90), .O(gate257inter3));
  inv1  gate1181(.a(s_91), .O(gate257inter4));
  nand2 gate1182(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate1183(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate1184(.a(G754), .O(gate257inter7));
  inv1  gate1185(.a(G755), .O(gate257inter8));
  nand2 gate1186(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate1187(.a(s_91), .b(gate257inter3), .O(gate257inter10));
  nor2  gate1188(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate1189(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate1190(.a(gate257inter12), .b(gate257inter1), .O(G770));

  xor2  gate1891(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate1892(.a(gate258inter0), .b(s_192), .O(gate258inter1));
  and2  gate1893(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate1894(.a(s_192), .O(gate258inter3));
  inv1  gate1895(.a(s_193), .O(gate258inter4));
  nand2 gate1896(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate1897(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate1898(.a(G756), .O(gate258inter7));
  inv1  gate1899(.a(G757), .O(gate258inter8));
  nand2 gate1900(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate1901(.a(s_193), .b(gate258inter3), .O(gate258inter10));
  nor2  gate1902(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate1903(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate1904(.a(gate258inter12), .b(gate258inter1), .O(G773));

  xor2  gate2143(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate2144(.a(gate259inter0), .b(s_228), .O(gate259inter1));
  and2  gate2145(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate2146(.a(s_228), .O(gate259inter3));
  inv1  gate2147(.a(s_229), .O(gate259inter4));
  nand2 gate2148(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate2149(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate2150(.a(G758), .O(gate259inter7));
  inv1  gate2151(.a(G759), .O(gate259inter8));
  nand2 gate2152(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate2153(.a(s_229), .b(gate259inter3), .O(gate259inter10));
  nor2  gate2154(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate2155(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate2156(.a(gate259inter12), .b(gate259inter1), .O(G776));
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate911(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate912(.a(gate263inter0), .b(s_52), .O(gate263inter1));
  and2  gate913(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate914(.a(s_52), .O(gate263inter3));
  inv1  gate915(.a(s_53), .O(gate263inter4));
  nand2 gate916(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate917(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate918(.a(G766), .O(gate263inter7));
  inv1  gate919(.a(G767), .O(gate263inter8));
  nand2 gate920(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate921(.a(s_53), .b(gate263inter3), .O(gate263inter10));
  nor2  gate922(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate923(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate924(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate1541(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate1542(.a(gate265inter0), .b(s_142), .O(gate265inter1));
  and2  gate1543(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate1544(.a(s_142), .O(gate265inter3));
  inv1  gate1545(.a(s_143), .O(gate265inter4));
  nand2 gate1546(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate1547(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate1548(.a(G642), .O(gate265inter7));
  inv1  gate1549(.a(G770), .O(gate265inter8));
  nand2 gate1550(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate1551(.a(s_143), .b(gate265inter3), .O(gate265inter10));
  nor2  gate1552(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate1553(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate1554(.a(gate265inter12), .b(gate265inter1), .O(G794));
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate1233(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate1234(.a(gate267inter0), .b(s_98), .O(gate267inter1));
  and2  gate1235(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate1236(.a(s_98), .O(gate267inter3));
  inv1  gate1237(.a(s_99), .O(gate267inter4));
  nand2 gate1238(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate1239(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate1240(.a(G648), .O(gate267inter7));
  inv1  gate1241(.a(G776), .O(gate267inter8));
  nand2 gate1242(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate1243(.a(s_99), .b(gate267inter3), .O(gate267inter10));
  nor2  gate1244(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate1245(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate1246(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate2787(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate2788(.a(gate269inter0), .b(s_320), .O(gate269inter1));
  and2  gate2789(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate2790(.a(s_320), .O(gate269inter3));
  inv1  gate2791(.a(s_321), .O(gate269inter4));
  nand2 gate2792(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate2793(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate2794(.a(G654), .O(gate269inter7));
  inv1  gate2795(.a(G782), .O(gate269inter8));
  nand2 gate2796(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate2797(.a(s_321), .b(gate269inter3), .O(gate269inter10));
  nor2  gate2798(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate2799(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate2800(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate2773(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate2774(.a(gate274inter0), .b(s_318), .O(gate274inter1));
  and2  gate2775(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate2776(.a(s_318), .O(gate274inter3));
  inv1  gate2777(.a(s_319), .O(gate274inter4));
  nand2 gate2778(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate2779(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate2780(.a(G770), .O(gate274inter7));
  inv1  gate2781(.a(G794), .O(gate274inter8));
  nand2 gate2782(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate2783(.a(s_319), .b(gate274inter3), .O(gate274inter10));
  nor2  gate2784(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate2785(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate2786(.a(gate274inter12), .b(gate274inter1), .O(G819));

  xor2  gate2437(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate2438(.a(gate275inter0), .b(s_270), .O(gate275inter1));
  and2  gate2439(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate2440(.a(s_270), .O(gate275inter3));
  inv1  gate2441(.a(s_271), .O(gate275inter4));
  nand2 gate2442(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate2443(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate2444(.a(G645), .O(gate275inter7));
  inv1  gate2445(.a(G797), .O(gate275inter8));
  nand2 gate2446(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate2447(.a(s_271), .b(gate275inter3), .O(gate275inter10));
  nor2  gate2448(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate2449(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate2450(.a(gate275inter12), .b(gate275inter1), .O(G820));

  xor2  gate715(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate716(.a(gate276inter0), .b(s_24), .O(gate276inter1));
  and2  gate717(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate718(.a(s_24), .O(gate276inter3));
  inv1  gate719(.a(s_25), .O(gate276inter4));
  nand2 gate720(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate721(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate722(.a(G773), .O(gate276inter7));
  inv1  gate723(.a(G797), .O(gate276inter8));
  nand2 gate724(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate725(.a(s_25), .b(gate276inter3), .O(gate276inter10));
  nor2  gate726(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate727(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate728(.a(gate276inter12), .b(gate276inter1), .O(G821));

  xor2  gate1821(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate1822(.a(gate277inter0), .b(s_182), .O(gate277inter1));
  and2  gate1823(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate1824(.a(s_182), .O(gate277inter3));
  inv1  gate1825(.a(s_183), .O(gate277inter4));
  nand2 gate1826(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate1827(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate1828(.a(G648), .O(gate277inter7));
  inv1  gate1829(.a(G800), .O(gate277inter8));
  nand2 gate1830(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate1831(.a(s_183), .b(gate277inter3), .O(gate277inter10));
  nor2  gate1832(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate1833(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate1834(.a(gate277inter12), .b(gate277inter1), .O(G822));

  xor2  gate1345(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate1346(.a(gate278inter0), .b(s_114), .O(gate278inter1));
  and2  gate1347(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate1348(.a(s_114), .O(gate278inter3));
  inv1  gate1349(.a(s_115), .O(gate278inter4));
  nand2 gate1350(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate1351(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate1352(.a(G776), .O(gate278inter7));
  inv1  gate1353(.a(G800), .O(gate278inter8));
  nand2 gate1354(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate1355(.a(s_115), .b(gate278inter3), .O(gate278inter10));
  nor2  gate1356(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate1357(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate1358(.a(gate278inter12), .b(gate278inter1), .O(G823));

  xor2  gate743(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate744(.a(gate279inter0), .b(s_28), .O(gate279inter1));
  and2  gate745(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate746(.a(s_28), .O(gate279inter3));
  inv1  gate747(.a(s_29), .O(gate279inter4));
  nand2 gate748(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate749(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate750(.a(G651), .O(gate279inter7));
  inv1  gate751(.a(G803), .O(gate279inter8));
  nand2 gate752(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate753(.a(s_29), .b(gate279inter3), .O(gate279inter10));
  nor2  gate754(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate755(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate756(.a(gate279inter12), .b(gate279inter1), .O(G824));

  xor2  gate2087(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate2088(.a(gate280inter0), .b(s_220), .O(gate280inter1));
  and2  gate2089(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate2090(.a(s_220), .O(gate280inter3));
  inv1  gate2091(.a(s_221), .O(gate280inter4));
  nand2 gate2092(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate2093(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate2094(.a(G779), .O(gate280inter7));
  inv1  gate2095(.a(G803), .O(gate280inter8));
  nand2 gate2096(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate2097(.a(s_221), .b(gate280inter3), .O(gate280inter10));
  nor2  gate2098(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate2099(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate2100(.a(gate280inter12), .b(gate280inter1), .O(G825));
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate2829(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate2830(.a(gate283inter0), .b(s_326), .O(gate283inter1));
  and2  gate2831(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate2832(.a(s_326), .O(gate283inter3));
  inv1  gate2833(.a(s_327), .O(gate283inter4));
  nand2 gate2834(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate2835(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate2836(.a(G657), .O(gate283inter7));
  inv1  gate2837(.a(G809), .O(gate283inter8));
  nand2 gate2838(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate2839(.a(s_327), .b(gate283inter3), .O(gate283inter10));
  nor2  gate2840(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate2841(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate2842(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate2059(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate2060(.a(gate285inter0), .b(s_216), .O(gate285inter1));
  and2  gate2061(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate2062(.a(s_216), .O(gate285inter3));
  inv1  gate2063(.a(s_217), .O(gate285inter4));
  nand2 gate2064(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate2065(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate2066(.a(G660), .O(gate285inter7));
  inv1  gate2067(.a(G812), .O(gate285inter8));
  nand2 gate2068(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate2069(.a(s_217), .b(gate285inter3), .O(gate285inter10));
  nor2  gate2070(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate2071(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate2072(.a(gate285inter12), .b(gate285inter1), .O(G830));

  xor2  gate939(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate940(.a(gate286inter0), .b(s_56), .O(gate286inter1));
  and2  gate941(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate942(.a(s_56), .O(gate286inter3));
  inv1  gate943(.a(s_57), .O(gate286inter4));
  nand2 gate944(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate945(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate946(.a(G788), .O(gate286inter7));
  inv1  gate947(.a(G812), .O(gate286inter8));
  nand2 gate948(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate949(.a(s_57), .b(gate286inter3), .O(gate286inter10));
  nor2  gate950(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate951(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate952(.a(gate286inter12), .b(gate286inter1), .O(G831));

  xor2  gate3039(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate3040(.a(gate287inter0), .b(s_356), .O(gate287inter1));
  and2  gate3041(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate3042(.a(s_356), .O(gate287inter3));
  inv1  gate3043(.a(s_357), .O(gate287inter4));
  nand2 gate3044(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate3045(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate3046(.a(G663), .O(gate287inter7));
  inv1  gate3047(.a(G815), .O(gate287inter8));
  nand2 gate3048(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate3049(.a(s_357), .b(gate287inter3), .O(gate287inter10));
  nor2  gate3050(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate3051(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate3052(.a(gate287inter12), .b(gate287inter1), .O(G832));

  xor2  gate1023(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate1024(.a(gate288inter0), .b(s_68), .O(gate288inter1));
  and2  gate1025(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate1026(.a(s_68), .O(gate288inter3));
  inv1  gate1027(.a(s_69), .O(gate288inter4));
  nand2 gate1028(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate1029(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate1030(.a(G791), .O(gate288inter7));
  inv1  gate1031(.a(G815), .O(gate288inter8));
  nand2 gate1032(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate1033(.a(s_69), .b(gate288inter3), .O(gate288inter10));
  nor2  gate1034(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate1035(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate1036(.a(gate288inter12), .b(gate288inter1), .O(G833));

  xor2  gate1415(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate1416(.a(gate289inter0), .b(s_124), .O(gate289inter1));
  and2  gate1417(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate1418(.a(s_124), .O(gate289inter3));
  inv1  gate1419(.a(s_125), .O(gate289inter4));
  nand2 gate1420(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate1421(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate1422(.a(G818), .O(gate289inter7));
  inv1  gate1423(.a(G819), .O(gate289inter8));
  nand2 gate1424(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate1425(.a(s_125), .b(gate289inter3), .O(gate289inter10));
  nor2  gate1426(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate1427(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate1428(.a(gate289inter12), .b(gate289inter1), .O(G834));

  xor2  gate2297(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate2298(.a(gate290inter0), .b(s_250), .O(gate290inter1));
  and2  gate2299(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate2300(.a(s_250), .O(gate290inter3));
  inv1  gate2301(.a(s_251), .O(gate290inter4));
  nand2 gate2302(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate2303(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate2304(.a(G820), .O(gate290inter7));
  inv1  gate2305(.a(G821), .O(gate290inter8));
  nand2 gate2306(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate2307(.a(s_251), .b(gate290inter3), .O(gate290inter10));
  nor2  gate2308(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate2309(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate2310(.a(gate290inter12), .b(gate290inter1), .O(G847));

  xor2  gate2549(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate2550(.a(gate291inter0), .b(s_286), .O(gate291inter1));
  and2  gate2551(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate2552(.a(s_286), .O(gate291inter3));
  inv1  gate2553(.a(s_287), .O(gate291inter4));
  nand2 gate2554(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate2555(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate2556(.a(G822), .O(gate291inter7));
  inv1  gate2557(.a(G823), .O(gate291inter8));
  nand2 gate2558(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate2559(.a(s_287), .b(gate291inter3), .O(gate291inter10));
  nor2  gate2560(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate2561(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate2562(.a(gate291inter12), .b(gate291inter1), .O(G860));

  xor2  gate2465(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate2466(.a(gate292inter0), .b(s_274), .O(gate292inter1));
  and2  gate2467(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate2468(.a(s_274), .O(gate292inter3));
  inv1  gate2469(.a(s_275), .O(gate292inter4));
  nand2 gate2470(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate2471(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate2472(.a(G824), .O(gate292inter7));
  inv1  gate2473(.a(G825), .O(gate292inter8));
  nand2 gate2474(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate2475(.a(s_275), .b(gate292inter3), .O(gate292inter10));
  nor2  gate2476(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate2477(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate2478(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate2479(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate2480(.a(gate294inter0), .b(s_276), .O(gate294inter1));
  and2  gate2481(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate2482(.a(s_276), .O(gate294inter3));
  inv1  gate2483(.a(s_277), .O(gate294inter4));
  nand2 gate2484(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate2485(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate2486(.a(G832), .O(gate294inter7));
  inv1  gate2487(.a(G833), .O(gate294inter8));
  nand2 gate2488(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate2489(.a(s_277), .b(gate294inter3), .O(gate294inter10));
  nor2  gate2490(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate2491(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate2492(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate2675(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate2676(.a(gate296inter0), .b(s_304), .O(gate296inter1));
  and2  gate2677(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate2678(.a(s_304), .O(gate296inter3));
  inv1  gate2679(.a(s_305), .O(gate296inter4));
  nand2 gate2680(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate2681(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate2682(.a(G826), .O(gate296inter7));
  inv1  gate2683(.a(G827), .O(gate296inter8));
  nand2 gate2684(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate2685(.a(s_305), .b(gate296inter3), .O(gate296inter10));
  nor2  gate2686(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate2687(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate2688(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate1779(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate1780(.a(gate391inter0), .b(s_176), .O(gate391inter1));
  and2  gate1781(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate1782(.a(s_176), .O(gate391inter3));
  inv1  gate1783(.a(s_177), .O(gate391inter4));
  nand2 gate1784(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate1785(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate1786(.a(G5), .O(gate391inter7));
  inv1  gate1787(.a(G1048), .O(gate391inter8));
  nand2 gate1788(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate1789(.a(s_177), .b(gate391inter3), .O(gate391inter10));
  nor2  gate1790(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate1791(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate1792(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate1331(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate1332(.a(gate393inter0), .b(s_112), .O(gate393inter1));
  and2  gate1333(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate1334(.a(s_112), .O(gate393inter3));
  inv1  gate1335(.a(s_113), .O(gate393inter4));
  nand2 gate1336(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate1337(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate1338(.a(G7), .O(gate393inter7));
  inv1  gate1339(.a(G1054), .O(gate393inter8));
  nand2 gate1340(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate1341(.a(s_113), .b(gate393inter3), .O(gate393inter10));
  nor2  gate1342(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate1343(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate1344(.a(gate393inter12), .b(gate393inter1), .O(G1150));

  xor2  gate3081(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate3082(.a(gate394inter0), .b(s_362), .O(gate394inter1));
  and2  gate3083(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate3084(.a(s_362), .O(gate394inter3));
  inv1  gate3085(.a(s_363), .O(gate394inter4));
  nand2 gate3086(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate3087(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate3088(.a(G8), .O(gate394inter7));
  inv1  gate3089(.a(G1057), .O(gate394inter8));
  nand2 gate3090(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate3091(.a(s_363), .b(gate394inter3), .O(gate394inter10));
  nor2  gate3092(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate3093(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate3094(.a(gate394inter12), .b(gate394inter1), .O(G1153));

  xor2  gate3109(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate3110(.a(gate395inter0), .b(s_366), .O(gate395inter1));
  and2  gate3111(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate3112(.a(s_366), .O(gate395inter3));
  inv1  gate3113(.a(s_367), .O(gate395inter4));
  nand2 gate3114(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate3115(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate3116(.a(G9), .O(gate395inter7));
  inv1  gate3117(.a(G1060), .O(gate395inter8));
  nand2 gate3118(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate3119(.a(s_367), .b(gate395inter3), .O(gate395inter10));
  nor2  gate3120(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate3121(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate3122(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate2899(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate2900(.a(gate397inter0), .b(s_336), .O(gate397inter1));
  and2  gate2901(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate2902(.a(s_336), .O(gate397inter3));
  inv1  gate2903(.a(s_337), .O(gate397inter4));
  nand2 gate2904(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate2905(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate2906(.a(G11), .O(gate397inter7));
  inv1  gate2907(.a(G1066), .O(gate397inter8));
  nand2 gate2908(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate2909(.a(s_337), .b(gate397inter3), .O(gate397inter10));
  nor2  gate2910(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate2911(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate2912(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate1919(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate1920(.a(gate402inter0), .b(s_196), .O(gate402inter1));
  and2  gate1921(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate1922(.a(s_196), .O(gate402inter3));
  inv1  gate1923(.a(s_197), .O(gate402inter4));
  nand2 gate1924(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate1925(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate1926(.a(G16), .O(gate402inter7));
  inv1  gate1927(.a(G1081), .O(gate402inter8));
  nand2 gate1928(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate1929(.a(s_197), .b(gate402inter3), .O(gate402inter10));
  nor2  gate1930(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate1931(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate1932(.a(gate402inter12), .b(gate402inter1), .O(G1177));
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate1065(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate1066(.a(gate407inter0), .b(s_74), .O(gate407inter1));
  and2  gate1067(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate1068(.a(s_74), .O(gate407inter3));
  inv1  gate1069(.a(s_75), .O(gate407inter4));
  nand2 gate1070(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate1071(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate1072(.a(G21), .O(gate407inter7));
  inv1  gate1073(.a(G1096), .O(gate407inter8));
  nand2 gate1074(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate1075(.a(s_75), .b(gate407inter3), .O(gate407inter10));
  nor2  gate1076(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate1077(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate1078(.a(gate407inter12), .b(gate407inter1), .O(G1192));

  xor2  gate3123(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate3124(.a(gate408inter0), .b(s_368), .O(gate408inter1));
  and2  gate3125(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate3126(.a(s_368), .O(gate408inter3));
  inv1  gate3127(.a(s_369), .O(gate408inter4));
  nand2 gate3128(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate3129(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate3130(.a(G22), .O(gate408inter7));
  inv1  gate3131(.a(G1099), .O(gate408inter8));
  nand2 gate3132(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate3133(.a(s_369), .b(gate408inter3), .O(gate408inter10));
  nor2  gate3134(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate3135(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate3136(.a(gate408inter12), .b(gate408inter1), .O(G1195));
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate2801(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate2802(.a(gate410inter0), .b(s_322), .O(gate410inter1));
  and2  gate2803(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate2804(.a(s_322), .O(gate410inter3));
  inv1  gate2805(.a(s_323), .O(gate410inter4));
  nand2 gate2806(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate2807(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate2808(.a(G24), .O(gate410inter7));
  inv1  gate2809(.a(G1105), .O(gate410inter8));
  nand2 gate2810(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate2811(.a(s_323), .b(gate410inter3), .O(gate410inter10));
  nor2  gate2812(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate2813(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate2814(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate729(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate730(.a(gate417inter0), .b(s_26), .O(gate417inter1));
  and2  gate731(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate732(.a(s_26), .O(gate417inter3));
  inv1  gate733(.a(s_27), .O(gate417inter4));
  nand2 gate734(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate735(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate736(.a(G31), .O(gate417inter7));
  inv1  gate737(.a(G1126), .O(gate417inter8));
  nand2 gate738(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate739(.a(s_27), .b(gate417inter3), .O(gate417inter10));
  nor2  gate740(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate741(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate742(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate1387(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate1388(.a(gate421inter0), .b(s_120), .O(gate421inter1));
  and2  gate1389(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate1390(.a(s_120), .O(gate421inter3));
  inv1  gate1391(.a(s_121), .O(gate421inter4));
  nand2 gate1392(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate1393(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate1394(.a(G2), .O(gate421inter7));
  inv1  gate1395(.a(G1135), .O(gate421inter8));
  nand2 gate1396(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate1397(.a(s_121), .b(gate421inter3), .O(gate421inter10));
  nor2  gate1398(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate1399(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate1400(.a(gate421inter12), .b(gate421inter1), .O(G1230));

  xor2  gate2199(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate2200(.a(gate422inter0), .b(s_236), .O(gate422inter1));
  and2  gate2201(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate2202(.a(s_236), .O(gate422inter3));
  inv1  gate2203(.a(s_237), .O(gate422inter4));
  nand2 gate2204(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate2205(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate2206(.a(G1039), .O(gate422inter7));
  inv1  gate2207(.a(G1135), .O(gate422inter8));
  nand2 gate2208(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate2209(.a(s_237), .b(gate422inter3), .O(gate422inter10));
  nor2  gate2210(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate2211(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate2212(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );

  xor2  gate1121(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate1122(.a(gate426inter0), .b(s_82), .O(gate426inter1));
  and2  gate1123(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate1124(.a(s_82), .O(gate426inter3));
  inv1  gate1125(.a(s_83), .O(gate426inter4));
  nand2 gate1126(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate1127(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate1128(.a(G1045), .O(gate426inter7));
  inv1  gate1129(.a(G1141), .O(gate426inter8));
  nand2 gate1130(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate1131(.a(s_83), .b(gate426inter3), .O(gate426inter10));
  nor2  gate1132(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate1133(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate1134(.a(gate426inter12), .b(gate426inter1), .O(G1235));

  xor2  gate2493(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate2494(.a(gate427inter0), .b(s_278), .O(gate427inter1));
  and2  gate2495(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate2496(.a(s_278), .O(gate427inter3));
  inv1  gate2497(.a(s_279), .O(gate427inter4));
  nand2 gate2498(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate2499(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate2500(.a(G5), .O(gate427inter7));
  inv1  gate2501(.a(G1144), .O(gate427inter8));
  nand2 gate2502(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate2503(.a(s_279), .b(gate427inter3), .O(gate427inter10));
  nor2  gate2504(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate2505(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate2506(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate2535(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate2536(.a(gate430inter0), .b(s_284), .O(gate430inter1));
  and2  gate2537(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate2538(.a(s_284), .O(gate430inter3));
  inv1  gate2539(.a(s_285), .O(gate430inter4));
  nand2 gate2540(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate2541(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate2542(.a(G1051), .O(gate430inter7));
  inv1  gate2543(.a(G1147), .O(gate430inter8));
  nand2 gate2544(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate2545(.a(s_285), .b(gate430inter3), .O(gate430inter10));
  nor2  gate2546(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate2547(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate2548(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate1583(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate1584(.a(gate432inter0), .b(s_148), .O(gate432inter1));
  and2  gate1585(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate1586(.a(s_148), .O(gate432inter3));
  inv1  gate1587(.a(s_149), .O(gate432inter4));
  nand2 gate1588(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate1589(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate1590(.a(G1054), .O(gate432inter7));
  inv1  gate1591(.a(G1150), .O(gate432inter8));
  nand2 gate1592(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate1593(.a(s_149), .b(gate432inter3), .O(gate432inter10));
  nor2  gate1594(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate1595(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate1596(.a(gate432inter12), .b(gate432inter1), .O(G1241));

  xor2  gate1723(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate1724(.a(gate433inter0), .b(s_168), .O(gate433inter1));
  and2  gate1725(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate1726(.a(s_168), .O(gate433inter3));
  inv1  gate1727(.a(s_169), .O(gate433inter4));
  nand2 gate1728(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate1729(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate1730(.a(G8), .O(gate433inter7));
  inv1  gate1731(.a(G1153), .O(gate433inter8));
  nand2 gate1732(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate1733(.a(s_169), .b(gate433inter3), .O(gate433inter10));
  nor2  gate1734(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate1735(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate1736(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate883(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate884(.a(gate438inter0), .b(s_48), .O(gate438inter1));
  and2  gate885(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate886(.a(s_48), .O(gate438inter3));
  inv1  gate887(.a(s_49), .O(gate438inter4));
  nand2 gate888(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate889(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate890(.a(G1063), .O(gate438inter7));
  inv1  gate891(.a(G1159), .O(gate438inter8));
  nand2 gate892(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate893(.a(s_49), .b(gate438inter3), .O(gate438inter10));
  nor2  gate894(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate895(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate896(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate2983(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate2984(.a(gate441inter0), .b(s_348), .O(gate441inter1));
  and2  gate2985(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate2986(.a(s_348), .O(gate441inter3));
  inv1  gate2987(.a(s_349), .O(gate441inter4));
  nand2 gate2988(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate2989(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate2990(.a(G12), .O(gate441inter7));
  inv1  gate2991(.a(G1165), .O(gate441inter8));
  nand2 gate2992(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate2993(.a(s_349), .b(gate441inter3), .O(gate441inter10));
  nor2  gate2994(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate2995(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate2996(.a(gate441inter12), .b(gate441inter1), .O(G1250));

  xor2  gate2353(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate2354(.a(gate442inter0), .b(s_258), .O(gate442inter1));
  and2  gate2355(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate2356(.a(s_258), .O(gate442inter3));
  inv1  gate2357(.a(s_259), .O(gate442inter4));
  nand2 gate2358(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate2359(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate2360(.a(G1069), .O(gate442inter7));
  inv1  gate2361(.a(G1165), .O(gate442inter8));
  nand2 gate2362(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate2363(.a(s_259), .b(gate442inter3), .O(gate442inter10));
  nor2  gate2364(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate2365(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate2366(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate2115(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate2116(.a(gate445inter0), .b(s_224), .O(gate445inter1));
  and2  gate2117(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate2118(.a(s_224), .O(gate445inter3));
  inv1  gate2119(.a(s_225), .O(gate445inter4));
  nand2 gate2120(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate2121(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate2122(.a(G14), .O(gate445inter7));
  inv1  gate2123(.a(G1171), .O(gate445inter8));
  nand2 gate2124(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate2125(.a(s_225), .b(gate445inter3), .O(gate445inter10));
  nor2  gate2126(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate2127(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate2128(.a(gate445inter12), .b(gate445inter1), .O(G1254));

  xor2  gate2647(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate2648(.a(gate446inter0), .b(s_300), .O(gate446inter1));
  and2  gate2649(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate2650(.a(s_300), .O(gate446inter3));
  inv1  gate2651(.a(s_301), .O(gate446inter4));
  nand2 gate2652(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate2653(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate2654(.a(G1075), .O(gate446inter7));
  inv1  gate2655(.a(G1171), .O(gate446inter8));
  nand2 gate2656(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate2657(.a(s_301), .b(gate446inter3), .O(gate446inter10));
  nor2  gate2658(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate2659(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate2660(.a(gate446inter12), .b(gate446inter1), .O(G1255));

  xor2  gate2213(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate2214(.a(gate447inter0), .b(s_238), .O(gate447inter1));
  and2  gate2215(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate2216(.a(s_238), .O(gate447inter3));
  inv1  gate2217(.a(s_239), .O(gate447inter4));
  nand2 gate2218(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate2219(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate2220(.a(G15), .O(gate447inter7));
  inv1  gate2221(.a(G1174), .O(gate447inter8));
  nand2 gate2222(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate2223(.a(s_239), .b(gate447inter3), .O(gate447inter10));
  nor2  gate2224(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate2225(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate2226(.a(gate447inter12), .b(gate447inter1), .O(G1256));

  xor2  gate701(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate702(.a(gate448inter0), .b(s_22), .O(gate448inter1));
  and2  gate703(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate704(.a(s_22), .O(gate448inter3));
  inv1  gate705(.a(s_23), .O(gate448inter4));
  nand2 gate706(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate707(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate708(.a(G1078), .O(gate448inter7));
  inv1  gate709(.a(G1174), .O(gate448inter8));
  nand2 gate710(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate711(.a(s_23), .b(gate448inter3), .O(gate448inter10));
  nor2  gate712(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate713(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate714(.a(gate448inter12), .b(gate448inter1), .O(G1257));

  xor2  gate1653(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate1654(.a(gate449inter0), .b(s_158), .O(gate449inter1));
  and2  gate1655(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate1656(.a(s_158), .O(gate449inter3));
  inv1  gate1657(.a(s_159), .O(gate449inter4));
  nand2 gate1658(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate1659(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate1660(.a(G16), .O(gate449inter7));
  inv1  gate1661(.a(G1177), .O(gate449inter8));
  nand2 gate1662(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate1663(.a(s_159), .b(gate449inter3), .O(gate449inter10));
  nor2  gate1664(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate1665(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate1666(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );

  xor2  gate2073(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate2074(.a(gate451inter0), .b(s_218), .O(gate451inter1));
  and2  gate2075(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate2076(.a(s_218), .O(gate451inter3));
  inv1  gate2077(.a(s_219), .O(gate451inter4));
  nand2 gate2078(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate2079(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate2080(.a(G17), .O(gate451inter7));
  inv1  gate2081(.a(G1180), .O(gate451inter8));
  nand2 gate2082(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate2083(.a(s_219), .b(gate451inter3), .O(gate451inter10));
  nor2  gate2084(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate2085(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate2086(.a(gate451inter12), .b(gate451inter1), .O(G1260));

  xor2  gate687(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate688(.a(gate452inter0), .b(s_20), .O(gate452inter1));
  and2  gate689(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate690(.a(s_20), .O(gate452inter3));
  inv1  gate691(.a(s_21), .O(gate452inter4));
  nand2 gate692(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate693(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate694(.a(G1084), .O(gate452inter7));
  inv1  gate695(.a(G1180), .O(gate452inter8));
  nand2 gate696(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate697(.a(s_21), .b(gate452inter3), .O(gate452inter10));
  nor2  gate698(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate699(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate700(.a(gate452inter12), .b(gate452inter1), .O(G1261));

  xor2  gate3193(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate3194(.a(gate453inter0), .b(s_378), .O(gate453inter1));
  and2  gate3195(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate3196(.a(s_378), .O(gate453inter3));
  inv1  gate3197(.a(s_379), .O(gate453inter4));
  nand2 gate3198(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate3199(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate3200(.a(G18), .O(gate453inter7));
  inv1  gate3201(.a(G1183), .O(gate453inter8));
  nand2 gate3202(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate3203(.a(s_379), .b(gate453inter3), .O(gate453inter10));
  nor2  gate3204(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate3205(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate3206(.a(gate453inter12), .b(gate453inter1), .O(G1262));

  xor2  gate1639(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate1640(.a(gate454inter0), .b(s_156), .O(gate454inter1));
  and2  gate1641(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate1642(.a(s_156), .O(gate454inter3));
  inv1  gate1643(.a(s_157), .O(gate454inter4));
  nand2 gate1644(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate1645(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate1646(.a(G1087), .O(gate454inter7));
  inv1  gate1647(.a(G1183), .O(gate454inter8));
  nand2 gate1648(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate1649(.a(s_157), .b(gate454inter3), .O(gate454inter10));
  nor2  gate1650(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate1651(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate1652(.a(gate454inter12), .b(gate454inter1), .O(G1263));
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate3137(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate3138(.a(gate457inter0), .b(s_370), .O(gate457inter1));
  and2  gate3139(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate3140(.a(s_370), .O(gate457inter3));
  inv1  gate3141(.a(s_371), .O(gate457inter4));
  nand2 gate3142(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate3143(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate3144(.a(G20), .O(gate457inter7));
  inv1  gate3145(.a(G1189), .O(gate457inter8));
  nand2 gate3146(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate3147(.a(s_371), .b(gate457inter3), .O(gate457inter10));
  nor2  gate3148(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate3149(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate3150(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate2619(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate2620(.a(gate460inter0), .b(s_296), .O(gate460inter1));
  and2  gate2621(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate2622(.a(s_296), .O(gate460inter3));
  inv1  gate2623(.a(s_297), .O(gate460inter4));
  nand2 gate2624(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate2625(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate2626(.a(G1096), .O(gate460inter7));
  inv1  gate2627(.a(G1192), .O(gate460inter8));
  nand2 gate2628(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate2629(.a(s_297), .b(gate460inter3), .O(gate460inter10));
  nor2  gate2630(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate2631(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate2632(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );

  xor2  gate1989(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate1990(.a(gate462inter0), .b(s_206), .O(gate462inter1));
  and2  gate1991(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate1992(.a(s_206), .O(gate462inter3));
  inv1  gate1993(.a(s_207), .O(gate462inter4));
  nand2 gate1994(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate1995(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate1996(.a(G1099), .O(gate462inter7));
  inv1  gate1997(.a(G1195), .O(gate462inter8));
  nand2 gate1998(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate1999(.a(s_207), .b(gate462inter3), .O(gate462inter10));
  nor2  gate2000(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate2001(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate2002(.a(gate462inter12), .b(gate462inter1), .O(G1271));

  xor2  gate2031(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate2032(.a(gate463inter0), .b(s_212), .O(gate463inter1));
  and2  gate2033(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate2034(.a(s_212), .O(gate463inter3));
  inv1  gate2035(.a(s_213), .O(gate463inter4));
  nand2 gate2036(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate2037(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate2038(.a(G23), .O(gate463inter7));
  inv1  gate2039(.a(G1198), .O(gate463inter8));
  nand2 gate2040(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate2041(.a(s_213), .b(gate463inter3), .O(gate463inter10));
  nor2  gate2042(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate2043(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate2044(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate827(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate828(.a(gate465inter0), .b(s_40), .O(gate465inter1));
  and2  gate829(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate830(.a(s_40), .O(gate465inter3));
  inv1  gate831(.a(s_41), .O(gate465inter4));
  nand2 gate832(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate833(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate834(.a(G24), .O(gate465inter7));
  inv1  gate835(.a(G1201), .O(gate465inter8));
  nand2 gate836(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate837(.a(s_41), .b(gate465inter3), .O(gate465inter10));
  nor2  gate838(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate839(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate840(.a(gate465inter12), .b(gate465inter1), .O(G1274));

  xor2  gate1807(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate1808(.a(gate466inter0), .b(s_180), .O(gate466inter1));
  and2  gate1809(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate1810(.a(s_180), .O(gate466inter3));
  inv1  gate1811(.a(s_181), .O(gate466inter4));
  nand2 gate1812(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate1813(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate1814(.a(G1105), .O(gate466inter7));
  inv1  gate1815(.a(G1201), .O(gate466inter8));
  nand2 gate1816(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate1817(.a(s_181), .b(gate466inter3), .O(gate466inter10));
  nor2  gate1818(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate1819(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate1820(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );

  xor2  gate2241(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate2242(.a(gate470inter0), .b(s_242), .O(gate470inter1));
  and2  gate2243(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate2244(.a(s_242), .O(gate470inter3));
  inv1  gate2245(.a(s_243), .O(gate470inter4));
  nand2 gate2246(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate2247(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate2248(.a(G1111), .O(gate470inter7));
  inv1  gate2249(.a(G1207), .O(gate470inter8));
  nand2 gate2250(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate2251(.a(s_243), .b(gate470inter3), .O(gate470inter10));
  nor2  gate2252(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate2253(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate2254(.a(gate470inter12), .b(gate470inter1), .O(G1279));

  xor2  gate2955(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate2956(.a(gate471inter0), .b(s_344), .O(gate471inter1));
  and2  gate2957(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate2958(.a(s_344), .O(gate471inter3));
  inv1  gate2959(.a(s_345), .O(gate471inter4));
  nand2 gate2960(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate2961(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate2962(.a(G27), .O(gate471inter7));
  inv1  gate2963(.a(G1210), .O(gate471inter8));
  nand2 gate2964(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate2965(.a(s_345), .b(gate471inter3), .O(gate471inter10));
  nor2  gate2966(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate2967(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate2968(.a(gate471inter12), .b(gate471inter1), .O(G1280));

  xor2  gate995(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate996(.a(gate472inter0), .b(s_64), .O(gate472inter1));
  and2  gate997(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate998(.a(s_64), .O(gate472inter3));
  inv1  gate999(.a(s_65), .O(gate472inter4));
  nand2 gate1000(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate1001(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate1002(.a(G1114), .O(gate472inter7));
  inv1  gate1003(.a(G1210), .O(gate472inter8));
  nand2 gate1004(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate1005(.a(s_65), .b(gate472inter3), .O(gate472inter10));
  nor2  gate1006(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate1007(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate1008(.a(gate472inter12), .b(gate472inter1), .O(G1281));

  xor2  gate841(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate842(.a(gate473inter0), .b(s_42), .O(gate473inter1));
  and2  gate843(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate844(.a(s_42), .O(gate473inter3));
  inv1  gate845(.a(s_43), .O(gate473inter4));
  nand2 gate846(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate847(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate848(.a(G28), .O(gate473inter7));
  inv1  gate849(.a(G1213), .O(gate473inter8));
  nand2 gate850(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate851(.a(s_43), .b(gate473inter3), .O(gate473inter10));
  nor2  gate852(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate853(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate854(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate2185(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate2186(.a(gate475inter0), .b(s_234), .O(gate475inter1));
  and2  gate2187(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate2188(.a(s_234), .O(gate475inter3));
  inv1  gate2189(.a(s_235), .O(gate475inter4));
  nand2 gate2190(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate2191(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate2192(.a(G29), .O(gate475inter7));
  inv1  gate2193(.a(G1216), .O(gate475inter8));
  nand2 gate2194(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate2195(.a(s_235), .b(gate475inter3), .O(gate475inter10));
  nor2  gate2196(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate2197(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate2198(.a(gate475inter12), .b(gate475inter1), .O(G1284));
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate2591(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate2592(.a(gate477inter0), .b(s_292), .O(gate477inter1));
  and2  gate2593(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate2594(.a(s_292), .O(gate477inter3));
  inv1  gate2595(.a(s_293), .O(gate477inter4));
  nand2 gate2596(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate2597(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate2598(.a(G30), .O(gate477inter7));
  inv1  gate2599(.a(G1219), .O(gate477inter8));
  nand2 gate2600(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate2601(.a(s_293), .b(gate477inter3), .O(gate477inter10));
  nor2  gate2602(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate2603(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate2604(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate2703(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate2704(.a(gate481inter0), .b(s_308), .O(gate481inter1));
  and2  gate2705(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate2706(.a(s_308), .O(gate481inter3));
  inv1  gate2707(.a(s_309), .O(gate481inter4));
  nand2 gate2708(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate2709(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate2710(.a(G32), .O(gate481inter7));
  inv1  gate2711(.a(G1225), .O(gate481inter8));
  nand2 gate2712(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate2713(.a(s_309), .b(gate481inter3), .O(gate481inter10));
  nor2  gate2714(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate2715(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate2716(.a(gate481inter12), .b(gate481inter1), .O(G1290));
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate1975(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate1976(.a(gate486inter0), .b(s_204), .O(gate486inter1));
  and2  gate1977(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate1978(.a(s_204), .O(gate486inter3));
  inv1  gate1979(.a(s_205), .O(gate486inter4));
  nand2 gate1980(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate1981(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate1982(.a(G1234), .O(gate486inter7));
  inv1  gate1983(.a(G1235), .O(gate486inter8));
  nand2 gate1984(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate1985(.a(s_205), .b(gate486inter3), .O(gate486inter10));
  nor2  gate1986(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate1987(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate1988(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate2045(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate2046(.a(gate490inter0), .b(s_214), .O(gate490inter1));
  and2  gate2047(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate2048(.a(s_214), .O(gate490inter3));
  inv1  gate2049(.a(s_215), .O(gate490inter4));
  nand2 gate2050(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate2051(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate2052(.a(G1242), .O(gate490inter7));
  inv1  gate2053(.a(G1243), .O(gate490inter8));
  nand2 gate2054(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate2055(.a(s_215), .b(gate490inter3), .O(gate490inter10));
  nor2  gate2056(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate2057(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate2058(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate1877(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate1878(.a(gate492inter0), .b(s_190), .O(gate492inter1));
  and2  gate1879(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate1880(.a(s_190), .O(gate492inter3));
  inv1  gate1881(.a(s_191), .O(gate492inter4));
  nand2 gate1882(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate1883(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate1884(.a(G1246), .O(gate492inter7));
  inv1  gate1885(.a(G1247), .O(gate492inter8));
  nand2 gate1886(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate1887(.a(s_191), .b(gate492inter3), .O(gate492inter10));
  nor2  gate1888(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate1889(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate1890(.a(gate492inter12), .b(gate492inter1), .O(G1301));

  xor2  gate3011(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate3012(.a(gate493inter0), .b(s_352), .O(gate493inter1));
  and2  gate3013(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate3014(.a(s_352), .O(gate493inter3));
  inv1  gate3015(.a(s_353), .O(gate493inter4));
  nand2 gate3016(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate3017(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate3018(.a(G1248), .O(gate493inter7));
  inv1  gate3019(.a(G1249), .O(gate493inter8));
  nand2 gate3020(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate3021(.a(s_353), .b(gate493inter3), .O(gate493inter10));
  nor2  gate3022(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate3023(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate3024(.a(gate493inter12), .b(gate493inter1), .O(G1302));

  xor2  gate1905(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1906(.a(gate494inter0), .b(s_194), .O(gate494inter1));
  and2  gate1907(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1908(.a(s_194), .O(gate494inter3));
  inv1  gate1909(.a(s_195), .O(gate494inter4));
  nand2 gate1910(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1911(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1912(.a(G1250), .O(gate494inter7));
  inv1  gate1913(.a(G1251), .O(gate494inter8));
  nand2 gate1914(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1915(.a(s_195), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1916(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1917(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1918(.a(gate494inter12), .b(gate494inter1), .O(G1303));

  xor2  gate2367(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate2368(.a(gate495inter0), .b(s_260), .O(gate495inter1));
  and2  gate2369(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate2370(.a(s_260), .O(gate495inter3));
  inv1  gate2371(.a(s_261), .O(gate495inter4));
  nand2 gate2372(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate2373(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate2374(.a(G1252), .O(gate495inter7));
  inv1  gate2375(.a(G1253), .O(gate495inter8));
  nand2 gate2376(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate2377(.a(s_261), .b(gate495inter3), .O(gate495inter10));
  nor2  gate2378(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate2379(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate2380(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate2717(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate2718(.a(gate499inter0), .b(s_310), .O(gate499inter1));
  and2  gate2719(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate2720(.a(s_310), .O(gate499inter3));
  inv1  gate2721(.a(s_311), .O(gate499inter4));
  nand2 gate2722(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate2723(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate2724(.a(G1260), .O(gate499inter7));
  inv1  gate2725(.a(G1261), .O(gate499inter8));
  nand2 gate2726(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate2727(.a(s_311), .b(gate499inter3), .O(gate499inter10));
  nor2  gate2728(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate2729(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate2730(.a(gate499inter12), .b(gate499inter1), .O(G1308));

  xor2  gate2381(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate2382(.a(gate500inter0), .b(s_262), .O(gate500inter1));
  and2  gate2383(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate2384(.a(s_262), .O(gate500inter3));
  inv1  gate2385(.a(s_263), .O(gate500inter4));
  nand2 gate2386(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate2387(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate2388(.a(G1262), .O(gate500inter7));
  inv1  gate2389(.a(G1263), .O(gate500inter8));
  nand2 gate2390(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate2391(.a(s_263), .b(gate500inter3), .O(gate500inter10));
  nor2  gate2392(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate2393(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate2394(.a(gate500inter12), .b(gate500inter1), .O(G1309));

  xor2  gate2129(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate2130(.a(gate501inter0), .b(s_226), .O(gate501inter1));
  and2  gate2131(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate2132(.a(s_226), .O(gate501inter3));
  inv1  gate2133(.a(s_227), .O(gate501inter4));
  nand2 gate2134(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate2135(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate2136(.a(G1264), .O(gate501inter7));
  inv1  gate2137(.a(G1265), .O(gate501inter8));
  nand2 gate2138(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate2139(.a(s_227), .b(gate501inter3), .O(gate501inter10));
  nor2  gate2140(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate2141(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate2142(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate3095(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate3096(.a(gate504inter0), .b(s_364), .O(gate504inter1));
  and2  gate3097(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate3098(.a(s_364), .O(gate504inter3));
  inv1  gate3099(.a(s_365), .O(gate504inter4));
  nand2 gate3100(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate3101(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate3102(.a(G1270), .O(gate504inter7));
  inv1  gate3103(.a(G1271), .O(gate504inter8));
  nand2 gate3104(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate3105(.a(s_365), .b(gate504inter3), .O(gate504inter10));
  nor2  gate3106(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate3107(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate3108(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );

  xor2  gate2871(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate2872(.a(gate507inter0), .b(s_332), .O(gate507inter1));
  and2  gate2873(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate2874(.a(s_332), .O(gate507inter3));
  inv1  gate2875(.a(s_333), .O(gate507inter4));
  nand2 gate2876(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate2877(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate2878(.a(G1276), .O(gate507inter7));
  inv1  gate2879(.a(G1277), .O(gate507inter8));
  nand2 gate2880(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate2881(.a(s_333), .b(gate507inter3), .O(gate507inter10));
  nor2  gate2882(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate2883(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate2884(.a(gate507inter12), .b(gate507inter1), .O(G1316));

  xor2  gate1205(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate1206(.a(gate508inter0), .b(s_94), .O(gate508inter1));
  and2  gate1207(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate1208(.a(s_94), .O(gate508inter3));
  inv1  gate1209(.a(s_95), .O(gate508inter4));
  nand2 gate1210(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate1211(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate1212(.a(G1278), .O(gate508inter7));
  inv1  gate1213(.a(G1279), .O(gate508inter8));
  nand2 gate1214(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate1215(.a(s_95), .b(gate508inter3), .O(gate508inter10));
  nor2  gate1216(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate1217(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate1218(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate2857(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate2858(.a(gate511inter0), .b(s_330), .O(gate511inter1));
  and2  gate2859(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate2860(.a(s_330), .O(gate511inter3));
  inv1  gate2861(.a(s_331), .O(gate511inter4));
  nand2 gate2862(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate2863(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate2864(.a(G1284), .O(gate511inter7));
  inv1  gate2865(.a(G1285), .O(gate511inter8));
  nand2 gate2866(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate2867(.a(s_331), .b(gate511inter3), .O(gate511inter10));
  nor2  gate2868(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate2869(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate2870(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );

  xor2  gate2311(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate2312(.a(gate513inter0), .b(s_252), .O(gate513inter1));
  and2  gate2313(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate2314(.a(s_252), .O(gate513inter3));
  inv1  gate2315(.a(s_253), .O(gate513inter4));
  nand2 gate2316(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate2317(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate2318(.a(G1288), .O(gate513inter7));
  inv1  gate2319(.a(G1289), .O(gate513inter8));
  nand2 gate2320(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate2321(.a(s_253), .b(gate513inter3), .O(gate513inter10));
  nor2  gate2322(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate2323(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate2324(.a(gate513inter12), .b(gate513inter1), .O(G1322));
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule