module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate1625(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate1626(.a(gate11inter0), .b(s_154), .O(gate11inter1));
  and2  gate1627(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate1628(.a(s_154), .O(gate11inter3));
  inv1  gate1629(.a(s_155), .O(gate11inter4));
  nand2 gate1630(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate1631(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate1632(.a(G5), .O(gate11inter7));
  inv1  gate1633(.a(G6), .O(gate11inter8));
  nand2 gate1634(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate1635(.a(s_155), .b(gate11inter3), .O(gate11inter10));
  nor2  gate1636(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate1637(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate1638(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate1023(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate1024(.a(gate16inter0), .b(s_68), .O(gate16inter1));
  and2  gate1025(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate1026(.a(s_68), .O(gate16inter3));
  inv1  gate1027(.a(s_69), .O(gate16inter4));
  nand2 gate1028(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate1029(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate1030(.a(G15), .O(gate16inter7));
  inv1  gate1031(.a(G16), .O(gate16inter8));
  nand2 gate1032(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate1033(.a(s_69), .b(gate16inter3), .O(gate16inter10));
  nor2  gate1034(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate1035(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate1036(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate827(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate828(.a(gate19inter0), .b(s_40), .O(gate19inter1));
  and2  gate829(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate830(.a(s_40), .O(gate19inter3));
  inv1  gate831(.a(s_41), .O(gate19inter4));
  nand2 gate832(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate833(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate834(.a(G21), .O(gate19inter7));
  inv1  gate835(.a(G22), .O(gate19inter8));
  nand2 gate836(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate837(.a(s_41), .b(gate19inter3), .O(gate19inter10));
  nor2  gate838(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate839(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate840(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate1261(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate1262(.a(gate21inter0), .b(s_102), .O(gate21inter1));
  and2  gate1263(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate1264(.a(s_102), .O(gate21inter3));
  inv1  gate1265(.a(s_103), .O(gate21inter4));
  nand2 gate1266(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate1267(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate1268(.a(G25), .O(gate21inter7));
  inv1  gate1269(.a(G26), .O(gate21inter8));
  nand2 gate1270(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate1271(.a(s_103), .b(gate21inter3), .O(gate21inter10));
  nor2  gate1272(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate1273(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate1274(.a(gate21inter12), .b(gate21inter1), .O(G302));

  xor2  gate1709(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate1710(.a(gate22inter0), .b(s_166), .O(gate22inter1));
  and2  gate1711(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate1712(.a(s_166), .O(gate22inter3));
  inv1  gate1713(.a(s_167), .O(gate22inter4));
  nand2 gate1714(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate1715(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate1716(.a(G27), .O(gate22inter7));
  inv1  gate1717(.a(G28), .O(gate22inter8));
  nand2 gate1718(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate1719(.a(s_167), .b(gate22inter3), .O(gate22inter10));
  nor2  gate1720(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate1721(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate1722(.a(gate22inter12), .b(gate22inter1), .O(G305));
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );

  xor2  gate1093(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate1094(.a(gate35inter0), .b(s_78), .O(gate35inter1));
  and2  gate1095(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate1096(.a(s_78), .O(gate35inter3));
  inv1  gate1097(.a(s_79), .O(gate35inter4));
  nand2 gate1098(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate1099(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate1100(.a(G18), .O(gate35inter7));
  inv1  gate1101(.a(G22), .O(gate35inter8));
  nand2 gate1102(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate1103(.a(s_79), .b(gate35inter3), .O(gate35inter10));
  nor2  gate1104(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate1105(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate1106(.a(gate35inter12), .b(gate35inter1), .O(G344));
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate1639(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate1640(.a(gate39inter0), .b(s_156), .O(gate39inter1));
  and2  gate1641(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate1642(.a(s_156), .O(gate39inter3));
  inv1  gate1643(.a(s_157), .O(gate39inter4));
  nand2 gate1644(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate1645(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate1646(.a(G20), .O(gate39inter7));
  inv1  gate1647(.a(G24), .O(gate39inter8));
  nand2 gate1648(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate1649(.a(s_157), .b(gate39inter3), .O(gate39inter10));
  nor2  gate1650(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate1651(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate1652(.a(gate39inter12), .b(gate39inter1), .O(G356));

  xor2  gate1065(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate1066(.a(gate40inter0), .b(s_74), .O(gate40inter1));
  and2  gate1067(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate1068(.a(s_74), .O(gate40inter3));
  inv1  gate1069(.a(s_75), .O(gate40inter4));
  nand2 gate1070(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate1071(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate1072(.a(G28), .O(gate40inter7));
  inv1  gate1073(.a(G32), .O(gate40inter8));
  nand2 gate1074(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate1075(.a(s_75), .b(gate40inter3), .O(gate40inter10));
  nor2  gate1076(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate1077(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate1078(.a(gate40inter12), .b(gate40inter1), .O(G359));
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate1303(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate1304(.a(gate43inter0), .b(s_108), .O(gate43inter1));
  and2  gate1305(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate1306(.a(s_108), .O(gate43inter3));
  inv1  gate1307(.a(s_109), .O(gate43inter4));
  nand2 gate1308(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate1309(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate1310(.a(G3), .O(gate43inter7));
  inv1  gate1311(.a(G269), .O(gate43inter8));
  nand2 gate1312(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate1313(.a(s_109), .b(gate43inter3), .O(gate43inter10));
  nor2  gate1314(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate1315(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate1316(.a(gate43inter12), .b(gate43inter1), .O(G364));
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate1149(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate1150(.a(gate51inter0), .b(s_86), .O(gate51inter1));
  and2  gate1151(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate1152(.a(s_86), .O(gate51inter3));
  inv1  gate1153(.a(s_87), .O(gate51inter4));
  nand2 gate1154(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate1155(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate1156(.a(G11), .O(gate51inter7));
  inv1  gate1157(.a(G281), .O(gate51inter8));
  nand2 gate1158(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate1159(.a(s_87), .b(gate51inter3), .O(gate51inter10));
  nor2  gate1160(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate1161(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate1162(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );

  xor2  gate1289(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate1290(.a(gate56inter0), .b(s_106), .O(gate56inter1));
  and2  gate1291(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate1292(.a(s_106), .O(gate56inter3));
  inv1  gate1293(.a(s_107), .O(gate56inter4));
  nand2 gate1294(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate1295(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate1296(.a(G16), .O(gate56inter7));
  inv1  gate1297(.a(G287), .O(gate56inter8));
  nand2 gate1298(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate1299(.a(s_107), .b(gate56inter3), .O(gate56inter10));
  nor2  gate1300(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate1301(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate1302(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate1191(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate1192(.a(gate59inter0), .b(s_92), .O(gate59inter1));
  and2  gate1193(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate1194(.a(s_92), .O(gate59inter3));
  inv1  gate1195(.a(s_93), .O(gate59inter4));
  nand2 gate1196(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate1197(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate1198(.a(G19), .O(gate59inter7));
  inv1  gate1199(.a(G293), .O(gate59inter8));
  nand2 gate1200(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate1201(.a(s_93), .b(gate59inter3), .O(gate59inter10));
  nor2  gate1202(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate1203(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate1204(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );

  xor2  gate1205(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate1206(.a(gate64inter0), .b(s_94), .O(gate64inter1));
  and2  gate1207(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate1208(.a(s_94), .O(gate64inter3));
  inv1  gate1209(.a(s_95), .O(gate64inter4));
  nand2 gate1210(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate1211(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate1212(.a(G24), .O(gate64inter7));
  inv1  gate1213(.a(G299), .O(gate64inter8));
  nand2 gate1214(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate1215(.a(s_95), .b(gate64inter3), .O(gate64inter10));
  nor2  gate1216(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate1217(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate1218(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate1681(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate1682(.a(gate74inter0), .b(s_162), .O(gate74inter1));
  and2  gate1683(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate1684(.a(s_162), .O(gate74inter3));
  inv1  gate1685(.a(s_163), .O(gate74inter4));
  nand2 gate1686(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate1687(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate1688(.a(G5), .O(gate74inter7));
  inv1  gate1689(.a(G314), .O(gate74inter8));
  nand2 gate1690(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate1691(.a(s_163), .b(gate74inter3), .O(gate74inter10));
  nor2  gate1692(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate1693(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate1694(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate1331(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate1332(.a(gate86inter0), .b(s_112), .O(gate86inter1));
  and2  gate1333(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate1334(.a(s_112), .O(gate86inter3));
  inv1  gate1335(.a(s_113), .O(gate86inter4));
  nand2 gate1336(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate1337(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate1338(.a(G8), .O(gate86inter7));
  inv1  gate1339(.a(G332), .O(gate86inter8));
  nand2 gate1340(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate1341(.a(s_113), .b(gate86inter3), .O(gate86inter10));
  nor2  gate1342(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate1343(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate1344(.a(gate86inter12), .b(gate86inter1), .O(G407));

  xor2  gate617(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate618(.a(gate87inter0), .b(s_10), .O(gate87inter1));
  and2  gate619(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate620(.a(s_10), .O(gate87inter3));
  inv1  gate621(.a(s_11), .O(gate87inter4));
  nand2 gate622(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate623(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate624(.a(G12), .O(gate87inter7));
  inv1  gate625(.a(G335), .O(gate87inter8));
  nand2 gate626(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate627(.a(s_11), .b(gate87inter3), .O(gate87inter10));
  nor2  gate628(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate629(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate630(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate589(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate590(.a(gate100inter0), .b(s_6), .O(gate100inter1));
  and2  gate591(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate592(.a(s_6), .O(gate100inter3));
  inv1  gate593(.a(s_7), .O(gate100inter4));
  nand2 gate594(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate595(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate596(.a(G31), .O(gate100inter7));
  inv1  gate597(.a(G353), .O(gate100inter8));
  nand2 gate598(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate599(.a(s_7), .b(gate100inter3), .O(gate100inter10));
  nor2  gate600(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate601(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate602(.a(gate100inter12), .b(gate100inter1), .O(G421));

  xor2  gate911(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate912(.a(gate101inter0), .b(s_52), .O(gate101inter1));
  and2  gate913(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate914(.a(s_52), .O(gate101inter3));
  inv1  gate915(.a(s_53), .O(gate101inter4));
  nand2 gate916(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate917(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate918(.a(G20), .O(gate101inter7));
  inv1  gate919(.a(G356), .O(gate101inter8));
  nand2 gate920(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate921(.a(s_53), .b(gate101inter3), .O(gate101inter10));
  nor2  gate922(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate923(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate924(.a(gate101inter12), .b(gate101inter1), .O(G422));

  xor2  gate1079(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate1080(.a(gate102inter0), .b(s_76), .O(gate102inter1));
  and2  gate1081(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate1082(.a(s_76), .O(gate102inter3));
  inv1  gate1083(.a(s_77), .O(gate102inter4));
  nand2 gate1084(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate1085(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate1086(.a(G24), .O(gate102inter7));
  inv1  gate1087(.a(G356), .O(gate102inter8));
  nand2 gate1088(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate1089(.a(s_77), .b(gate102inter3), .O(gate102inter10));
  nor2  gate1090(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate1091(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate1092(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate1611(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate1612(.a(gate104inter0), .b(s_152), .O(gate104inter1));
  and2  gate1613(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate1614(.a(s_152), .O(gate104inter3));
  inv1  gate1615(.a(s_153), .O(gate104inter4));
  nand2 gate1616(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate1617(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate1618(.a(G32), .O(gate104inter7));
  inv1  gate1619(.a(G359), .O(gate104inter8));
  nand2 gate1620(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate1621(.a(s_153), .b(gate104inter3), .O(gate104inter10));
  nor2  gate1622(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate1623(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate1624(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate1443(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate1444(.a(gate106inter0), .b(s_128), .O(gate106inter1));
  and2  gate1445(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate1446(.a(s_128), .O(gate106inter3));
  inv1  gate1447(.a(s_129), .O(gate106inter4));
  nand2 gate1448(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate1449(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate1450(.a(G364), .O(gate106inter7));
  inv1  gate1451(.a(G365), .O(gate106inter8));
  nand2 gate1452(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate1453(.a(s_129), .b(gate106inter3), .O(gate106inter10));
  nor2  gate1454(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate1455(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate1456(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate1597(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate1598(.a(gate112inter0), .b(s_150), .O(gate112inter1));
  and2  gate1599(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate1600(.a(s_150), .O(gate112inter3));
  inv1  gate1601(.a(s_151), .O(gate112inter4));
  nand2 gate1602(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate1603(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate1604(.a(G376), .O(gate112inter7));
  inv1  gate1605(.a(G377), .O(gate112inter8));
  nand2 gate1606(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate1607(.a(s_151), .b(gate112inter3), .O(gate112inter10));
  nor2  gate1608(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate1609(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate1610(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );

  xor2  gate1219(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate1220(.a(gate114inter0), .b(s_96), .O(gate114inter1));
  and2  gate1221(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate1222(.a(s_96), .O(gate114inter3));
  inv1  gate1223(.a(s_97), .O(gate114inter4));
  nand2 gate1224(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate1225(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate1226(.a(G380), .O(gate114inter7));
  inv1  gate1227(.a(G381), .O(gate114inter8));
  nand2 gate1228(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate1229(.a(s_97), .b(gate114inter3), .O(gate114inter10));
  nor2  gate1230(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate1231(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate1232(.a(gate114inter12), .b(gate114inter1), .O(G453));
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );

  xor2  gate785(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate786(.a(gate122inter0), .b(s_34), .O(gate122inter1));
  and2  gate787(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate788(.a(s_34), .O(gate122inter3));
  inv1  gate789(.a(s_35), .O(gate122inter4));
  nand2 gate790(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate791(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate792(.a(G396), .O(gate122inter7));
  inv1  gate793(.a(G397), .O(gate122inter8));
  nand2 gate794(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate795(.a(s_35), .b(gate122inter3), .O(gate122inter10));
  nor2  gate796(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate797(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate798(.a(gate122inter12), .b(gate122inter1), .O(G477));
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate1555(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate1556(.a(gate126inter0), .b(s_144), .O(gate126inter1));
  and2  gate1557(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate1558(.a(s_144), .O(gate126inter3));
  inv1  gate1559(.a(s_145), .O(gate126inter4));
  nand2 gate1560(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate1561(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate1562(.a(G404), .O(gate126inter7));
  inv1  gate1563(.a(G405), .O(gate126inter8));
  nand2 gate1564(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate1565(.a(s_145), .b(gate126inter3), .O(gate126inter10));
  nor2  gate1566(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate1567(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate1568(.a(gate126inter12), .b(gate126inter1), .O(G489));

  xor2  gate1723(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate1724(.a(gate127inter0), .b(s_168), .O(gate127inter1));
  and2  gate1725(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate1726(.a(s_168), .O(gate127inter3));
  inv1  gate1727(.a(s_169), .O(gate127inter4));
  nand2 gate1728(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate1729(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate1730(.a(G406), .O(gate127inter7));
  inv1  gate1731(.a(G407), .O(gate127inter8));
  nand2 gate1732(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate1733(.a(s_169), .b(gate127inter3), .O(gate127inter10));
  nor2  gate1734(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate1735(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate1736(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );

  xor2  gate1373(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate1374(.a(gate134inter0), .b(s_118), .O(gate134inter1));
  and2  gate1375(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate1376(.a(s_118), .O(gate134inter3));
  inv1  gate1377(.a(s_119), .O(gate134inter4));
  nand2 gate1378(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate1379(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate1380(.a(G420), .O(gate134inter7));
  inv1  gate1381(.a(G421), .O(gate134inter8));
  nand2 gate1382(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate1383(.a(s_119), .b(gate134inter3), .O(gate134inter10));
  nor2  gate1384(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate1385(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate1386(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate1009(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate1010(.a(gate143inter0), .b(s_66), .O(gate143inter1));
  and2  gate1011(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate1012(.a(s_66), .O(gate143inter3));
  inv1  gate1013(.a(s_67), .O(gate143inter4));
  nand2 gate1014(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate1015(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate1016(.a(G462), .O(gate143inter7));
  inv1  gate1017(.a(G465), .O(gate143inter8));
  nand2 gate1018(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate1019(.a(s_67), .b(gate143inter3), .O(gate143inter10));
  nor2  gate1020(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate1021(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate1022(.a(gate143inter12), .b(gate143inter1), .O(G540));
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate981(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate982(.a(gate149inter0), .b(s_62), .O(gate149inter1));
  and2  gate983(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate984(.a(s_62), .O(gate149inter3));
  inv1  gate985(.a(s_63), .O(gate149inter4));
  nand2 gate986(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate987(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate988(.a(G498), .O(gate149inter7));
  inv1  gate989(.a(G501), .O(gate149inter8));
  nand2 gate990(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate991(.a(s_63), .b(gate149inter3), .O(gate149inter10));
  nor2  gate992(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate993(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate994(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate1485(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate1486(.a(gate156inter0), .b(s_134), .O(gate156inter1));
  and2  gate1487(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate1488(.a(s_134), .O(gate156inter3));
  inv1  gate1489(.a(s_135), .O(gate156inter4));
  nand2 gate1490(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate1491(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate1492(.a(G435), .O(gate156inter7));
  inv1  gate1493(.a(G525), .O(gate156inter8));
  nand2 gate1494(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate1495(.a(s_135), .b(gate156inter3), .O(gate156inter10));
  nor2  gate1496(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate1497(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate1498(.a(gate156inter12), .b(gate156inter1), .O(G573));

  xor2  gate1583(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate1584(.a(gate157inter0), .b(s_148), .O(gate157inter1));
  and2  gate1585(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate1586(.a(s_148), .O(gate157inter3));
  inv1  gate1587(.a(s_149), .O(gate157inter4));
  nand2 gate1588(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate1589(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate1590(.a(G438), .O(gate157inter7));
  inv1  gate1591(.a(G528), .O(gate157inter8));
  nand2 gate1592(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate1593(.a(s_149), .b(gate157inter3), .O(gate157inter10));
  nor2  gate1594(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate1595(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate1596(.a(gate157inter12), .b(gate157inter1), .O(G574));

  xor2  gate813(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate814(.a(gate158inter0), .b(s_38), .O(gate158inter1));
  and2  gate815(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate816(.a(s_38), .O(gate158inter3));
  inv1  gate817(.a(s_39), .O(gate158inter4));
  nand2 gate818(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate819(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate820(.a(G441), .O(gate158inter7));
  inv1  gate821(.a(G528), .O(gate158inter8));
  nand2 gate822(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate823(.a(s_39), .b(gate158inter3), .O(gate158inter10));
  nor2  gate824(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate825(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate826(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );

  xor2  gate631(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate632(.a(gate171inter0), .b(s_12), .O(gate171inter1));
  and2  gate633(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate634(.a(s_12), .O(gate171inter3));
  inv1  gate635(.a(s_13), .O(gate171inter4));
  nand2 gate636(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate637(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate638(.a(G480), .O(gate171inter7));
  inv1  gate639(.a(G549), .O(gate171inter8));
  nand2 gate640(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate641(.a(s_13), .b(gate171inter3), .O(gate171inter10));
  nor2  gate642(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate643(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate644(.a(gate171inter12), .b(gate171inter1), .O(G588));
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate799(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate800(.a(gate186inter0), .b(s_36), .O(gate186inter1));
  and2  gate801(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate802(.a(s_36), .O(gate186inter3));
  inv1  gate803(.a(s_37), .O(gate186inter4));
  nand2 gate804(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate805(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate806(.a(G572), .O(gate186inter7));
  inv1  gate807(.a(G573), .O(gate186inter8));
  nand2 gate808(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate809(.a(s_37), .b(gate186inter3), .O(gate186inter10));
  nor2  gate810(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate811(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate812(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate995(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate996(.a(gate190inter0), .b(s_64), .O(gate190inter1));
  and2  gate997(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate998(.a(s_64), .O(gate190inter3));
  inv1  gate999(.a(s_65), .O(gate190inter4));
  nand2 gate1000(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate1001(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate1002(.a(G580), .O(gate190inter7));
  inv1  gate1003(.a(G581), .O(gate190inter8));
  nand2 gate1004(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate1005(.a(s_65), .b(gate190inter3), .O(gate190inter10));
  nor2  gate1006(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate1007(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate1008(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );

  xor2  gate883(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate884(.a(gate192inter0), .b(s_48), .O(gate192inter1));
  and2  gate885(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate886(.a(s_48), .O(gate192inter3));
  inv1  gate887(.a(s_49), .O(gate192inter4));
  nand2 gate888(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate889(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate890(.a(G584), .O(gate192inter7));
  inv1  gate891(.a(G585), .O(gate192inter8));
  nand2 gate892(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate893(.a(s_49), .b(gate192inter3), .O(gate192inter10));
  nor2  gate894(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate895(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate896(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate1345(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate1346(.a(gate195inter0), .b(s_114), .O(gate195inter1));
  and2  gate1347(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate1348(.a(s_114), .O(gate195inter3));
  inv1  gate1349(.a(s_115), .O(gate195inter4));
  nand2 gate1350(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate1351(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate1352(.a(G590), .O(gate195inter7));
  inv1  gate1353(.a(G591), .O(gate195inter8));
  nand2 gate1354(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate1355(.a(s_115), .b(gate195inter3), .O(gate195inter10));
  nor2  gate1356(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate1357(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate1358(.a(gate195inter12), .b(gate195inter1), .O(G648));

  xor2  gate1471(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate1472(.a(gate196inter0), .b(s_132), .O(gate196inter1));
  and2  gate1473(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate1474(.a(s_132), .O(gate196inter3));
  inv1  gate1475(.a(s_133), .O(gate196inter4));
  nand2 gate1476(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate1477(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate1478(.a(G592), .O(gate196inter7));
  inv1  gate1479(.a(G593), .O(gate196inter8));
  nand2 gate1480(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate1481(.a(s_133), .b(gate196inter3), .O(gate196inter10));
  nor2  gate1482(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate1483(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate1484(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );

  xor2  gate701(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate702(.a(gate202inter0), .b(s_22), .O(gate202inter1));
  and2  gate703(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate704(.a(s_22), .O(gate202inter3));
  inv1  gate705(.a(s_23), .O(gate202inter4));
  nand2 gate706(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate707(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate708(.a(G612), .O(gate202inter7));
  inv1  gate709(.a(G617), .O(gate202inter8));
  nand2 gate710(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate711(.a(s_23), .b(gate202inter3), .O(gate202inter10));
  nor2  gate712(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate713(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate714(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );

  xor2  gate939(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate940(.a(gate210inter0), .b(s_56), .O(gate210inter1));
  and2  gate941(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate942(.a(s_56), .O(gate210inter3));
  inv1  gate943(.a(s_57), .O(gate210inter4));
  nand2 gate944(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate945(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate946(.a(G607), .O(gate210inter7));
  inv1  gate947(.a(G666), .O(gate210inter8));
  nand2 gate948(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate949(.a(s_57), .b(gate210inter3), .O(gate210inter10));
  nor2  gate950(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate951(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate952(.a(gate210inter12), .b(gate210inter1), .O(G691));
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate757(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate758(.a(gate214inter0), .b(s_30), .O(gate214inter1));
  and2  gate759(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate760(.a(s_30), .O(gate214inter3));
  inv1  gate761(.a(s_31), .O(gate214inter4));
  nand2 gate762(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate763(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate764(.a(G612), .O(gate214inter7));
  inv1  gate765(.a(G672), .O(gate214inter8));
  nand2 gate766(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate767(.a(s_31), .b(gate214inter3), .O(gate214inter10));
  nor2  gate768(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate769(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate770(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );

  xor2  gate1457(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate1458(.a(gate232inter0), .b(s_130), .O(gate232inter1));
  and2  gate1459(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate1460(.a(s_130), .O(gate232inter3));
  inv1  gate1461(.a(s_131), .O(gate232inter4));
  nand2 gate1462(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate1463(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate1464(.a(G704), .O(gate232inter7));
  inv1  gate1465(.a(G705), .O(gate232inter8));
  nand2 gate1466(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate1467(.a(s_131), .b(gate232inter3), .O(gate232inter10));
  nor2  gate1468(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate1469(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate1470(.a(gate232inter12), .b(gate232inter1), .O(G727));
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );

  xor2  gate855(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate856(.a(gate246inter0), .b(s_44), .O(gate246inter1));
  and2  gate857(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate858(.a(s_44), .O(gate246inter3));
  inv1  gate859(.a(s_45), .O(gate246inter4));
  nand2 gate860(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate861(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate862(.a(G724), .O(gate246inter7));
  inv1  gate863(.a(G736), .O(gate246inter8));
  nand2 gate864(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate865(.a(s_45), .b(gate246inter3), .O(gate246inter10));
  nor2  gate866(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate867(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate868(.a(gate246inter12), .b(gate246inter1), .O(G759));

  xor2  gate1415(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate1416(.a(gate247inter0), .b(s_124), .O(gate247inter1));
  and2  gate1417(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate1418(.a(s_124), .O(gate247inter3));
  inv1  gate1419(.a(s_125), .O(gate247inter4));
  nand2 gate1420(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate1421(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate1422(.a(G251), .O(gate247inter7));
  inv1  gate1423(.a(G739), .O(gate247inter8));
  nand2 gate1424(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate1425(.a(s_125), .b(gate247inter3), .O(gate247inter10));
  nor2  gate1426(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate1427(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate1428(.a(gate247inter12), .b(gate247inter1), .O(G760));
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate1037(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate1038(.a(gate253inter0), .b(s_70), .O(gate253inter1));
  and2  gate1039(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate1040(.a(s_70), .O(gate253inter3));
  inv1  gate1041(.a(s_71), .O(gate253inter4));
  nand2 gate1042(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate1043(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate1044(.a(G260), .O(gate253inter7));
  inv1  gate1045(.a(G748), .O(gate253inter8));
  nand2 gate1046(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate1047(.a(s_71), .b(gate253inter3), .O(gate253inter10));
  nor2  gate1048(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate1049(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate1050(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate1527(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate1528(.a(gate257inter0), .b(s_140), .O(gate257inter1));
  and2  gate1529(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate1530(.a(s_140), .O(gate257inter3));
  inv1  gate1531(.a(s_141), .O(gate257inter4));
  nand2 gate1532(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate1533(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate1534(.a(G754), .O(gate257inter7));
  inv1  gate1535(.a(G755), .O(gate257inter8));
  nand2 gate1536(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate1537(.a(s_141), .b(gate257inter3), .O(gate257inter10));
  nor2  gate1538(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate1539(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate1540(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate1121(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate1122(.a(gate262inter0), .b(s_82), .O(gate262inter1));
  and2  gate1123(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate1124(.a(s_82), .O(gate262inter3));
  inv1  gate1125(.a(s_83), .O(gate262inter4));
  nand2 gate1126(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate1127(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate1128(.a(G764), .O(gate262inter7));
  inv1  gate1129(.a(G765), .O(gate262inter8));
  nand2 gate1130(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate1131(.a(s_83), .b(gate262inter3), .O(gate262inter10));
  nor2  gate1132(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate1133(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate1134(.a(gate262inter12), .b(gate262inter1), .O(G785));

  xor2  gate1359(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate1360(.a(gate263inter0), .b(s_116), .O(gate263inter1));
  and2  gate1361(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate1362(.a(s_116), .O(gate263inter3));
  inv1  gate1363(.a(s_117), .O(gate263inter4));
  nand2 gate1364(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate1365(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate1366(.a(G766), .O(gate263inter7));
  inv1  gate1367(.a(G767), .O(gate263inter8));
  nand2 gate1368(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate1369(.a(s_117), .b(gate263inter3), .O(gate263inter10));
  nor2  gate1370(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate1371(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate1372(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate715(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate716(.a(gate272inter0), .b(s_24), .O(gate272inter1));
  and2  gate717(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate718(.a(s_24), .O(gate272inter3));
  inv1  gate719(.a(s_25), .O(gate272inter4));
  nand2 gate720(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate721(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate722(.a(G663), .O(gate272inter7));
  inv1  gate723(.a(G791), .O(gate272inter8));
  nand2 gate724(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate725(.a(s_25), .b(gate272inter3), .O(gate272inter10));
  nor2  gate726(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate727(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate728(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate1317(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate1318(.a(gate283inter0), .b(s_110), .O(gate283inter1));
  and2  gate1319(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate1320(.a(s_110), .O(gate283inter3));
  inv1  gate1321(.a(s_111), .O(gate283inter4));
  nand2 gate1322(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate1323(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate1324(.a(G657), .O(gate283inter7));
  inv1  gate1325(.a(G809), .O(gate283inter8));
  nand2 gate1326(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate1327(.a(s_111), .b(gate283inter3), .O(gate283inter10));
  nor2  gate1328(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate1329(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate1330(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate1163(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate1164(.a(gate291inter0), .b(s_88), .O(gate291inter1));
  and2  gate1165(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate1166(.a(s_88), .O(gate291inter3));
  inv1  gate1167(.a(s_89), .O(gate291inter4));
  nand2 gate1168(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate1169(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate1170(.a(G822), .O(gate291inter7));
  inv1  gate1171(.a(G823), .O(gate291inter8));
  nand2 gate1172(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate1173(.a(s_89), .b(gate291inter3), .O(gate291inter10));
  nor2  gate1174(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate1175(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate1176(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate1401(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate1402(.a(gate294inter0), .b(s_122), .O(gate294inter1));
  and2  gate1403(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate1404(.a(s_122), .O(gate294inter3));
  inv1  gate1405(.a(s_123), .O(gate294inter4));
  nand2 gate1406(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate1407(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate1408(.a(G832), .O(gate294inter7));
  inv1  gate1409(.a(G833), .O(gate294inter8));
  nand2 gate1410(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate1411(.a(s_123), .b(gate294inter3), .O(gate294inter10));
  nor2  gate1412(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate1413(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate1414(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate897(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate898(.a(gate391inter0), .b(s_50), .O(gate391inter1));
  and2  gate899(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate900(.a(s_50), .O(gate391inter3));
  inv1  gate901(.a(s_51), .O(gate391inter4));
  nand2 gate902(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate903(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate904(.a(G5), .O(gate391inter7));
  inv1  gate905(.a(G1048), .O(gate391inter8));
  nand2 gate906(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate907(.a(s_51), .b(gate391inter3), .O(gate391inter10));
  nor2  gate908(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate909(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate910(.a(gate391inter12), .b(gate391inter1), .O(G1144));

  xor2  gate547(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate548(.a(gate392inter0), .b(s_0), .O(gate392inter1));
  and2  gate549(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate550(.a(s_0), .O(gate392inter3));
  inv1  gate551(.a(s_1), .O(gate392inter4));
  nand2 gate552(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate553(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate554(.a(G6), .O(gate392inter7));
  inv1  gate555(.a(G1051), .O(gate392inter8));
  nand2 gate556(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate557(.a(s_1), .b(gate392inter3), .O(gate392inter10));
  nor2  gate558(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate559(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate560(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate645(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate646(.a(gate395inter0), .b(s_14), .O(gate395inter1));
  and2  gate647(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate648(.a(s_14), .O(gate395inter3));
  inv1  gate649(.a(s_15), .O(gate395inter4));
  nand2 gate650(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate651(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate652(.a(G9), .O(gate395inter7));
  inv1  gate653(.a(G1060), .O(gate395inter8));
  nand2 gate654(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate655(.a(s_15), .b(gate395inter3), .O(gate395inter10));
  nor2  gate656(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate657(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate658(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate603(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate604(.a(gate400inter0), .b(s_8), .O(gate400inter1));
  and2  gate605(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate606(.a(s_8), .O(gate400inter3));
  inv1  gate607(.a(s_9), .O(gate400inter4));
  nand2 gate608(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate609(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate610(.a(G14), .O(gate400inter7));
  inv1  gate611(.a(G1075), .O(gate400inter8));
  nand2 gate612(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate613(.a(s_9), .b(gate400inter3), .O(gate400inter10));
  nor2  gate614(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate615(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate616(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate1695(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate1696(.a(gate413inter0), .b(s_164), .O(gate413inter1));
  and2  gate1697(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate1698(.a(s_164), .O(gate413inter3));
  inv1  gate1699(.a(s_165), .O(gate413inter4));
  nand2 gate1700(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1701(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1702(.a(G27), .O(gate413inter7));
  inv1  gate1703(.a(G1114), .O(gate413inter8));
  nand2 gate1704(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1705(.a(s_165), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1706(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1707(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1708(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );

  xor2  gate1135(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate1136(.a(gate416inter0), .b(s_84), .O(gate416inter1));
  and2  gate1137(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate1138(.a(s_84), .O(gate416inter3));
  inv1  gate1139(.a(s_85), .O(gate416inter4));
  nand2 gate1140(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate1141(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate1142(.a(G30), .O(gate416inter7));
  inv1  gate1143(.a(G1123), .O(gate416inter8));
  nand2 gate1144(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate1145(.a(s_85), .b(gate416inter3), .O(gate416inter10));
  nor2  gate1146(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate1147(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate1148(.a(gate416inter12), .b(gate416inter1), .O(G1219));

  xor2  gate1667(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate1668(.a(gate417inter0), .b(s_160), .O(gate417inter1));
  and2  gate1669(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate1670(.a(s_160), .O(gate417inter3));
  inv1  gate1671(.a(s_161), .O(gate417inter4));
  nand2 gate1672(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate1673(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate1674(.a(G31), .O(gate417inter7));
  inv1  gate1675(.a(G1126), .O(gate417inter8));
  nand2 gate1676(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate1677(.a(s_161), .b(gate417inter3), .O(gate417inter10));
  nor2  gate1678(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate1679(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate1680(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate1513(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate1514(.a(gate421inter0), .b(s_138), .O(gate421inter1));
  and2  gate1515(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate1516(.a(s_138), .O(gate421inter3));
  inv1  gate1517(.a(s_139), .O(gate421inter4));
  nand2 gate1518(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate1519(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate1520(.a(G2), .O(gate421inter7));
  inv1  gate1521(.a(G1135), .O(gate421inter8));
  nand2 gate1522(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate1523(.a(s_139), .b(gate421inter3), .O(gate421inter10));
  nor2  gate1524(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate1525(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate1526(.a(gate421inter12), .b(gate421inter1), .O(G1230));
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );

  xor2  gate1541(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate1542(.a(gate423inter0), .b(s_142), .O(gate423inter1));
  and2  gate1543(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate1544(.a(s_142), .O(gate423inter3));
  inv1  gate1545(.a(s_143), .O(gate423inter4));
  nand2 gate1546(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate1547(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate1548(.a(G3), .O(gate423inter7));
  inv1  gate1549(.a(G1138), .O(gate423inter8));
  nand2 gate1550(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate1551(.a(s_143), .b(gate423inter3), .O(gate423inter10));
  nor2  gate1552(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate1553(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate1554(.a(gate423inter12), .b(gate423inter1), .O(G1232));
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );

  xor2  gate687(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate688(.a(gate427inter0), .b(s_20), .O(gate427inter1));
  and2  gate689(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate690(.a(s_20), .O(gate427inter3));
  inv1  gate691(.a(s_21), .O(gate427inter4));
  nand2 gate692(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate693(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate694(.a(G5), .O(gate427inter7));
  inv1  gate695(.a(G1144), .O(gate427inter8));
  nand2 gate696(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate697(.a(s_21), .b(gate427inter3), .O(gate427inter10));
  nor2  gate698(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate699(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate700(.a(gate427inter12), .b(gate427inter1), .O(G1236));

  xor2  gate967(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate968(.a(gate428inter0), .b(s_60), .O(gate428inter1));
  and2  gate969(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate970(.a(s_60), .O(gate428inter3));
  inv1  gate971(.a(s_61), .O(gate428inter4));
  nand2 gate972(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate973(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate974(.a(G1048), .O(gate428inter7));
  inv1  gate975(.a(G1144), .O(gate428inter8));
  nand2 gate976(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate977(.a(s_61), .b(gate428inter3), .O(gate428inter10));
  nor2  gate978(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate979(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate980(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate1569(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate1570(.a(gate430inter0), .b(s_146), .O(gate430inter1));
  and2  gate1571(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate1572(.a(s_146), .O(gate430inter3));
  inv1  gate1573(.a(s_147), .O(gate430inter4));
  nand2 gate1574(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate1575(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate1576(.a(G1051), .O(gate430inter7));
  inv1  gate1577(.a(G1147), .O(gate430inter8));
  nand2 gate1578(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate1579(.a(s_147), .b(gate430inter3), .O(gate430inter10));
  nor2  gate1580(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate1581(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate1582(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate1653(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate1654(.a(gate432inter0), .b(s_158), .O(gate432inter1));
  and2  gate1655(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate1656(.a(s_158), .O(gate432inter3));
  inv1  gate1657(.a(s_159), .O(gate432inter4));
  nand2 gate1658(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate1659(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate1660(.a(G1054), .O(gate432inter7));
  inv1  gate1661(.a(G1150), .O(gate432inter8));
  nand2 gate1662(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate1663(.a(s_159), .b(gate432inter3), .O(gate432inter10));
  nor2  gate1664(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate1665(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate1666(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate869(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate870(.a(gate437inter0), .b(s_46), .O(gate437inter1));
  and2  gate871(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate872(.a(s_46), .O(gate437inter3));
  inv1  gate873(.a(s_47), .O(gate437inter4));
  nand2 gate874(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate875(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate876(.a(G10), .O(gate437inter7));
  inv1  gate877(.a(G1159), .O(gate437inter8));
  nand2 gate878(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate879(.a(s_47), .b(gate437inter3), .O(gate437inter10));
  nor2  gate880(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate881(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate882(.a(gate437inter12), .b(gate437inter1), .O(G1246));

  xor2  gate771(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate772(.a(gate438inter0), .b(s_32), .O(gate438inter1));
  and2  gate773(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate774(.a(s_32), .O(gate438inter3));
  inv1  gate775(.a(s_33), .O(gate438inter4));
  nand2 gate776(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate777(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate778(.a(G1063), .O(gate438inter7));
  inv1  gate779(.a(G1159), .O(gate438inter8));
  nand2 gate780(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate781(.a(s_33), .b(gate438inter3), .O(gate438inter10));
  nor2  gate782(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate783(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate784(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate1247(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate1248(.a(gate442inter0), .b(s_100), .O(gate442inter1));
  and2  gate1249(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate1250(.a(s_100), .O(gate442inter3));
  inv1  gate1251(.a(s_101), .O(gate442inter4));
  nand2 gate1252(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate1253(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate1254(.a(G1069), .O(gate442inter7));
  inv1  gate1255(.a(G1165), .O(gate442inter8));
  nand2 gate1256(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate1257(.a(s_101), .b(gate442inter3), .O(gate442inter10));
  nor2  gate1258(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate1259(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate1260(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );

  xor2  gate841(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate842(.a(gate446inter0), .b(s_42), .O(gate446inter1));
  and2  gate843(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate844(.a(s_42), .O(gate446inter3));
  inv1  gate845(.a(s_43), .O(gate446inter4));
  nand2 gate846(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate847(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate848(.a(G1075), .O(gate446inter7));
  inv1  gate849(.a(G1171), .O(gate446inter8));
  nand2 gate850(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate851(.a(s_43), .b(gate446inter3), .O(gate446inter10));
  nor2  gate852(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate853(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate854(.a(gate446inter12), .b(gate446inter1), .O(G1255));

  xor2  gate1499(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate1500(.a(gate447inter0), .b(s_136), .O(gate447inter1));
  and2  gate1501(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate1502(.a(s_136), .O(gate447inter3));
  inv1  gate1503(.a(s_137), .O(gate447inter4));
  nand2 gate1504(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate1505(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate1506(.a(G15), .O(gate447inter7));
  inv1  gate1507(.a(G1174), .O(gate447inter8));
  nand2 gate1508(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate1509(.a(s_137), .b(gate447inter3), .O(gate447inter10));
  nor2  gate1510(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate1511(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate1512(.a(gate447inter12), .b(gate447inter1), .O(G1256));
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );

  xor2  gate1177(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate1178(.a(gate449inter0), .b(s_90), .O(gate449inter1));
  and2  gate1179(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate1180(.a(s_90), .O(gate449inter3));
  inv1  gate1181(.a(s_91), .O(gate449inter4));
  nand2 gate1182(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate1183(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate1184(.a(G16), .O(gate449inter7));
  inv1  gate1185(.a(G1177), .O(gate449inter8));
  nand2 gate1186(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate1187(.a(s_91), .b(gate449inter3), .O(gate449inter10));
  nor2  gate1188(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate1189(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate1190(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate743(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate744(.a(gate465inter0), .b(s_28), .O(gate465inter1));
  and2  gate745(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate746(.a(s_28), .O(gate465inter3));
  inv1  gate747(.a(s_29), .O(gate465inter4));
  nand2 gate748(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate749(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate750(.a(G24), .O(gate465inter7));
  inv1  gate751(.a(G1201), .O(gate465inter8));
  nand2 gate752(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate753(.a(s_29), .b(gate465inter3), .O(gate465inter10));
  nor2  gate754(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate755(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate756(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate673(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate674(.a(gate472inter0), .b(s_18), .O(gate472inter1));
  and2  gate675(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate676(.a(s_18), .O(gate472inter3));
  inv1  gate677(.a(s_19), .O(gate472inter4));
  nand2 gate678(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate679(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate680(.a(G1114), .O(gate472inter7));
  inv1  gate681(.a(G1210), .O(gate472inter8));
  nand2 gate682(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate683(.a(s_19), .b(gate472inter3), .O(gate472inter10));
  nor2  gate684(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate685(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate686(.a(gate472inter12), .b(gate472inter1), .O(G1281));

  xor2  gate561(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate562(.a(gate473inter0), .b(s_2), .O(gate473inter1));
  and2  gate563(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate564(.a(s_2), .O(gate473inter3));
  inv1  gate565(.a(s_3), .O(gate473inter4));
  nand2 gate566(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate567(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate568(.a(G28), .O(gate473inter7));
  inv1  gate569(.a(G1213), .O(gate473inter8));
  nand2 gate570(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate571(.a(s_3), .b(gate473inter3), .O(gate473inter10));
  nor2  gate572(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate573(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate574(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );

  xor2  gate1275(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate1276(.a(gate478inter0), .b(s_104), .O(gate478inter1));
  and2  gate1277(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate1278(.a(s_104), .O(gate478inter3));
  inv1  gate1279(.a(s_105), .O(gate478inter4));
  nand2 gate1280(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate1281(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate1282(.a(G1123), .O(gate478inter7));
  inv1  gate1283(.a(G1219), .O(gate478inter8));
  nand2 gate1284(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate1285(.a(s_105), .b(gate478inter3), .O(gate478inter10));
  nor2  gate1286(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate1287(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate1288(.a(gate478inter12), .b(gate478inter1), .O(G1287));

  xor2  gate1737(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate1738(.a(gate479inter0), .b(s_170), .O(gate479inter1));
  and2  gate1739(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate1740(.a(s_170), .O(gate479inter3));
  inv1  gate1741(.a(s_171), .O(gate479inter4));
  nand2 gate1742(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate1743(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate1744(.a(G31), .O(gate479inter7));
  inv1  gate1745(.a(G1222), .O(gate479inter8));
  nand2 gate1746(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate1747(.a(s_171), .b(gate479inter3), .O(gate479inter10));
  nor2  gate1748(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate1749(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate1750(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );

  xor2  gate953(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate954(.a(gate484inter0), .b(s_58), .O(gate484inter1));
  and2  gate955(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate956(.a(s_58), .O(gate484inter3));
  inv1  gate957(.a(s_59), .O(gate484inter4));
  nand2 gate958(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate959(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate960(.a(G1230), .O(gate484inter7));
  inv1  gate961(.a(G1231), .O(gate484inter8));
  nand2 gate962(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate963(.a(s_59), .b(gate484inter3), .O(gate484inter10));
  nor2  gate964(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate965(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate966(.a(gate484inter12), .b(gate484inter1), .O(G1293));
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate1429(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate1430(.a(gate486inter0), .b(s_126), .O(gate486inter1));
  and2  gate1431(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate1432(.a(s_126), .O(gate486inter3));
  inv1  gate1433(.a(s_127), .O(gate486inter4));
  nand2 gate1434(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate1435(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate1436(.a(G1234), .O(gate486inter7));
  inv1  gate1437(.a(G1235), .O(gate486inter8));
  nand2 gate1438(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate1439(.a(s_127), .b(gate486inter3), .O(gate486inter10));
  nor2  gate1440(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate1441(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate1442(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate1387(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate1388(.a(gate488inter0), .b(s_120), .O(gate488inter1));
  and2  gate1389(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate1390(.a(s_120), .O(gate488inter3));
  inv1  gate1391(.a(s_121), .O(gate488inter4));
  nand2 gate1392(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate1393(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate1394(.a(G1238), .O(gate488inter7));
  inv1  gate1395(.a(G1239), .O(gate488inter8));
  nand2 gate1396(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate1397(.a(s_121), .b(gate488inter3), .O(gate488inter10));
  nor2  gate1398(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate1399(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate1400(.a(gate488inter12), .b(gate488inter1), .O(G1297));

  xor2  gate729(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate730(.a(gate489inter0), .b(s_26), .O(gate489inter1));
  and2  gate731(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate732(.a(s_26), .O(gate489inter3));
  inv1  gate733(.a(s_27), .O(gate489inter4));
  nand2 gate734(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate735(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate736(.a(G1240), .O(gate489inter7));
  inv1  gate737(.a(G1241), .O(gate489inter8));
  nand2 gate738(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate739(.a(s_27), .b(gate489inter3), .O(gate489inter10));
  nor2  gate740(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate741(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate742(.a(gate489inter12), .b(gate489inter1), .O(G1298));

  xor2  gate575(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate576(.a(gate490inter0), .b(s_4), .O(gate490inter1));
  and2  gate577(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate578(.a(s_4), .O(gate490inter3));
  inv1  gate579(.a(s_5), .O(gate490inter4));
  nand2 gate580(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate581(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate582(.a(G1242), .O(gate490inter7));
  inv1  gate583(.a(G1243), .O(gate490inter8));
  nand2 gate584(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate585(.a(s_5), .b(gate490inter3), .O(gate490inter10));
  nor2  gate586(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate587(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate588(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );

  xor2  gate1051(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate1052(.a(gate495inter0), .b(s_72), .O(gate495inter1));
  and2  gate1053(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate1054(.a(s_72), .O(gate495inter3));
  inv1  gate1055(.a(s_73), .O(gate495inter4));
  nand2 gate1056(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate1057(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate1058(.a(G1252), .O(gate495inter7));
  inv1  gate1059(.a(G1253), .O(gate495inter8));
  nand2 gate1060(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate1061(.a(s_73), .b(gate495inter3), .O(gate495inter10));
  nor2  gate1062(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate1063(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate1064(.a(gate495inter12), .b(gate495inter1), .O(G1304));

  xor2  gate925(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate926(.a(gate496inter0), .b(s_54), .O(gate496inter1));
  and2  gate927(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate928(.a(s_54), .O(gate496inter3));
  inv1  gate929(.a(s_55), .O(gate496inter4));
  nand2 gate930(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate931(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate932(.a(G1254), .O(gate496inter7));
  inv1  gate933(.a(G1255), .O(gate496inter8));
  nand2 gate934(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate935(.a(s_55), .b(gate496inter3), .O(gate496inter10));
  nor2  gate936(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate937(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate938(.a(gate496inter12), .b(gate496inter1), .O(G1305));
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate1107(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate1108(.a(gate504inter0), .b(s_80), .O(gate504inter1));
  and2  gate1109(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate1110(.a(s_80), .O(gate504inter3));
  inv1  gate1111(.a(s_81), .O(gate504inter4));
  nand2 gate1112(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate1113(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate1114(.a(G1270), .O(gate504inter7));
  inv1  gate1115(.a(G1271), .O(gate504inter8));
  nand2 gate1116(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate1117(.a(s_81), .b(gate504inter3), .O(gate504inter10));
  nor2  gate1118(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate1119(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate1120(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate659(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate660(.a(gate511inter0), .b(s_16), .O(gate511inter1));
  and2  gate661(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate662(.a(s_16), .O(gate511inter3));
  inv1  gate663(.a(s_17), .O(gate511inter4));
  nand2 gate664(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate665(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate666(.a(G1284), .O(gate511inter7));
  inv1  gate667(.a(G1285), .O(gate511inter8));
  nand2 gate668(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate669(.a(s_17), .b(gate511inter3), .O(gate511inter10));
  nor2  gate670(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate671(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate672(.a(gate511inter12), .b(gate511inter1), .O(G1320));

  xor2  gate1233(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate1234(.a(gate512inter0), .b(s_98), .O(gate512inter1));
  and2  gate1235(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate1236(.a(s_98), .O(gate512inter3));
  inv1  gate1237(.a(s_99), .O(gate512inter4));
  nand2 gate1238(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate1239(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate1240(.a(G1286), .O(gate512inter7));
  inv1  gate1241(.a(G1287), .O(gate512inter8));
  nand2 gate1242(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate1243(.a(s_99), .b(gate512inter3), .O(gate512inter10));
  nor2  gate1244(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate1245(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate1246(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule