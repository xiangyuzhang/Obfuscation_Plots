module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate715(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate716(.a(gate9inter0), .b(s_24), .O(gate9inter1));
  and2  gate717(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate718(.a(s_24), .O(gate9inter3));
  inv1  gate719(.a(s_25), .O(gate9inter4));
  nand2 gate720(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate721(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate722(.a(G1), .O(gate9inter7));
  inv1  gate723(.a(G2), .O(gate9inter8));
  nand2 gate724(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate725(.a(s_25), .b(gate9inter3), .O(gate9inter10));
  nor2  gate726(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate727(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate728(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate1289(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate1290(.a(gate13inter0), .b(s_106), .O(gate13inter1));
  and2  gate1291(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate1292(.a(s_106), .O(gate13inter3));
  inv1  gate1293(.a(s_107), .O(gate13inter4));
  nand2 gate1294(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate1295(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate1296(.a(G9), .O(gate13inter7));
  inv1  gate1297(.a(G10), .O(gate13inter8));
  nand2 gate1298(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate1299(.a(s_107), .b(gate13inter3), .O(gate13inter10));
  nor2  gate1300(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate1301(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate1302(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate1345(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate1346(.a(gate16inter0), .b(s_114), .O(gate16inter1));
  and2  gate1347(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate1348(.a(s_114), .O(gate16inter3));
  inv1  gate1349(.a(s_115), .O(gate16inter4));
  nand2 gate1350(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate1351(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate1352(.a(G15), .O(gate16inter7));
  inv1  gate1353(.a(G16), .O(gate16inter8));
  nand2 gate1354(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate1355(.a(s_115), .b(gate16inter3), .O(gate16inter10));
  nor2  gate1356(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate1357(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate1358(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate1695(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate1696(.a(gate21inter0), .b(s_164), .O(gate21inter1));
  and2  gate1697(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate1698(.a(s_164), .O(gate21inter3));
  inv1  gate1699(.a(s_165), .O(gate21inter4));
  nand2 gate1700(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate1701(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate1702(.a(G25), .O(gate21inter7));
  inv1  gate1703(.a(G26), .O(gate21inter8));
  nand2 gate1704(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate1705(.a(s_165), .b(gate21inter3), .O(gate21inter10));
  nor2  gate1706(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate1707(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate1708(.a(gate21inter12), .b(gate21inter1), .O(G302));
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate1359(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate1360(.a(gate24inter0), .b(s_116), .O(gate24inter1));
  and2  gate1361(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate1362(.a(s_116), .O(gate24inter3));
  inv1  gate1363(.a(s_117), .O(gate24inter4));
  nand2 gate1364(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate1365(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate1366(.a(G31), .O(gate24inter7));
  inv1  gate1367(.a(G32), .O(gate24inter8));
  nand2 gate1368(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate1369(.a(s_117), .b(gate24inter3), .O(gate24inter10));
  nor2  gate1370(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate1371(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate1372(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );

  xor2  gate1569(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate1570(.a(gate35inter0), .b(s_146), .O(gate35inter1));
  and2  gate1571(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate1572(.a(s_146), .O(gate35inter3));
  inv1  gate1573(.a(s_147), .O(gate35inter4));
  nand2 gate1574(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate1575(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate1576(.a(G18), .O(gate35inter7));
  inv1  gate1577(.a(G22), .O(gate35inter8));
  nand2 gate1578(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate1579(.a(s_147), .b(gate35inter3), .O(gate35inter10));
  nor2  gate1580(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate1581(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate1582(.a(gate35inter12), .b(gate35inter1), .O(G344));
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );

  xor2  gate1219(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate1220(.a(gate42inter0), .b(s_96), .O(gate42inter1));
  and2  gate1221(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate1222(.a(s_96), .O(gate42inter3));
  inv1  gate1223(.a(s_97), .O(gate42inter4));
  nand2 gate1224(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate1225(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate1226(.a(G2), .O(gate42inter7));
  inv1  gate1227(.a(G266), .O(gate42inter8));
  nand2 gate1228(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate1229(.a(s_97), .b(gate42inter3), .O(gate42inter10));
  nor2  gate1230(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate1231(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate1232(.a(gate42inter12), .b(gate42inter1), .O(G363));

  xor2  gate1429(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate1430(.a(gate43inter0), .b(s_126), .O(gate43inter1));
  and2  gate1431(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate1432(.a(s_126), .O(gate43inter3));
  inv1  gate1433(.a(s_127), .O(gate43inter4));
  nand2 gate1434(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate1435(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate1436(.a(G3), .O(gate43inter7));
  inv1  gate1437(.a(G269), .O(gate43inter8));
  nand2 gate1438(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate1439(.a(s_127), .b(gate43inter3), .O(gate43inter10));
  nor2  gate1440(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate1441(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate1442(.a(gate43inter12), .b(gate43inter1), .O(G364));
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate1751(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate1752(.a(gate46inter0), .b(s_172), .O(gate46inter1));
  and2  gate1753(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate1754(.a(s_172), .O(gate46inter3));
  inv1  gate1755(.a(s_173), .O(gate46inter4));
  nand2 gate1756(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate1757(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate1758(.a(G6), .O(gate46inter7));
  inv1  gate1759(.a(G272), .O(gate46inter8));
  nand2 gate1760(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate1761(.a(s_173), .b(gate46inter3), .O(gate46inter10));
  nor2  gate1762(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate1763(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate1764(.a(gate46inter12), .b(gate46inter1), .O(G367));

  xor2  gate1009(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate1010(.a(gate47inter0), .b(s_66), .O(gate47inter1));
  and2  gate1011(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate1012(.a(s_66), .O(gate47inter3));
  inv1  gate1013(.a(s_67), .O(gate47inter4));
  nand2 gate1014(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate1015(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate1016(.a(G7), .O(gate47inter7));
  inv1  gate1017(.a(G275), .O(gate47inter8));
  nand2 gate1018(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate1019(.a(s_67), .b(gate47inter3), .O(gate47inter10));
  nor2  gate1020(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate1021(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate1022(.a(gate47inter12), .b(gate47inter1), .O(G368));
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate1625(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate1626(.a(gate52inter0), .b(s_154), .O(gate52inter1));
  and2  gate1627(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate1628(.a(s_154), .O(gate52inter3));
  inv1  gate1629(.a(s_155), .O(gate52inter4));
  nand2 gate1630(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate1631(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate1632(.a(G12), .O(gate52inter7));
  inv1  gate1633(.a(G281), .O(gate52inter8));
  nand2 gate1634(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate1635(.a(s_155), .b(gate52inter3), .O(gate52inter10));
  nor2  gate1636(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate1637(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate1638(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );

  xor2  gate603(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate604(.a(gate61inter0), .b(s_8), .O(gate61inter1));
  and2  gate605(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate606(.a(s_8), .O(gate61inter3));
  inv1  gate607(.a(s_9), .O(gate61inter4));
  nand2 gate608(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate609(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate610(.a(G21), .O(gate61inter7));
  inv1  gate611(.a(G296), .O(gate61inter8));
  nand2 gate612(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate613(.a(s_9), .b(gate61inter3), .O(gate61inter10));
  nor2  gate614(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate615(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate616(.a(gate61inter12), .b(gate61inter1), .O(G382));

  xor2  gate967(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate968(.a(gate62inter0), .b(s_60), .O(gate62inter1));
  and2  gate969(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate970(.a(s_60), .O(gate62inter3));
  inv1  gate971(.a(s_61), .O(gate62inter4));
  nand2 gate972(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate973(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate974(.a(G22), .O(gate62inter7));
  inv1  gate975(.a(G296), .O(gate62inter8));
  nand2 gate976(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate977(.a(s_61), .b(gate62inter3), .O(gate62inter10));
  nor2  gate978(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate979(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate980(.a(gate62inter12), .b(gate62inter1), .O(G383));

  xor2  gate1499(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate1500(.a(gate63inter0), .b(s_136), .O(gate63inter1));
  and2  gate1501(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate1502(.a(s_136), .O(gate63inter3));
  inv1  gate1503(.a(s_137), .O(gate63inter4));
  nand2 gate1504(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate1505(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate1506(.a(G23), .O(gate63inter7));
  inv1  gate1507(.a(G299), .O(gate63inter8));
  nand2 gate1508(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate1509(.a(s_137), .b(gate63inter3), .O(gate63inter10));
  nor2  gate1510(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate1511(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate1512(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate1765(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate1766(.a(gate65inter0), .b(s_174), .O(gate65inter1));
  and2  gate1767(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate1768(.a(s_174), .O(gate65inter3));
  inv1  gate1769(.a(s_175), .O(gate65inter4));
  nand2 gate1770(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate1771(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate1772(.a(G25), .O(gate65inter7));
  inv1  gate1773(.a(G302), .O(gate65inter8));
  nand2 gate1774(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate1775(.a(s_175), .b(gate65inter3), .O(gate65inter10));
  nor2  gate1776(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate1777(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate1778(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate1065(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate1066(.a(gate77inter0), .b(s_74), .O(gate77inter1));
  and2  gate1067(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate1068(.a(s_74), .O(gate77inter3));
  inv1  gate1069(.a(s_75), .O(gate77inter4));
  nand2 gate1070(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate1071(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate1072(.a(G2), .O(gate77inter7));
  inv1  gate1073(.a(G320), .O(gate77inter8));
  nand2 gate1074(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate1075(.a(s_75), .b(gate77inter3), .O(gate77inter10));
  nor2  gate1076(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate1077(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate1078(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );

  xor2  gate855(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate856(.a(gate83inter0), .b(s_44), .O(gate83inter1));
  and2  gate857(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate858(.a(s_44), .O(gate83inter3));
  inv1  gate859(.a(s_45), .O(gate83inter4));
  nand2 gate860(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate861(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate862(.a(G11), .O(gate83inter7));
  inv1  gate863(.a(G329), .O(gate83inter8));
  nand2 gate864(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate865(.a(s_45), .b(gate83inter3), .O(gate83inter10));
  nor2  gate866(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate867(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate868(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate771(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate772(.a(gate85inter0), .b(s_32), .O(gate85inter1));
  and2  gate773(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate774(.a(s_32), .O(gate85inter3));
  inv1  gate775(.a(s_33), .O(gate85inter4));
  nand2 gate776(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate777(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate778(.a(G4), .O(gate85inter7));
  inv1  gate779(.a(G332), .O(gate85inter8));
  nand2 gate780(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate781(.a(s_33), .b(gate85inter3), .O(gate85inter10));
  nor2  gate782(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate783(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate784(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );

  xor2  gate925(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate926(.a(gate87inter0), .b(s_54), .O(gate87inter1));
  and2  gate927(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate928(.a(s_54), .O(gate87inter3));
  inv1  gate929(.a(s_55), .O(gate87inter4));
  nand2 gate930(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate931(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate932(.a(G12), .O(gate87inter7));
  inv1  gate933(.a(G335), .O(gate87inter8));
  nand2 gate934(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate935(.a(s_55), .b(gate87inter3), .O(gate87inter10));
  nor2  gate936(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate937(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate938(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate1107(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate1108(.a(gate90inter0), .b(s_80), .O(gate90inter1));
  and2  gate1109(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate1110(.a(s_80), .O(gate90inter3));
  inv1  gate1111(.a(s_81), .O(gate90inter4));
  nand2 gate1112(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate1113(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate1114(.a(G21), .O(gate90inter7));
  inv1  gate1115(.a(G338), .O(gate90inter8));
  nand2 gate1116(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate1117(.a(s_81), .b(gate90inter3), .O(gate90inter10));
  nor2  gate1118(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate1119(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate1120(.a(gate90inter12), .b(gate90inter1), .O(G411));
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate1415(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate1416(.a(gate96inter0), .b(s_124), .O(gate96inter1));
  and2  gate1417(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate1418(.a(s_124), .O(gate96inter3));
  inv1  gate1419(.a(s_125), .O(gate96inter4));
  nand2 gate1420(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate1421(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate1422(.a(G30), .O(gate96inter7));
  inv1  gate1423(.a(G347), .O(gate96inter8));
  nand2 gate1424(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate1425(.a(s_125), .b(gate96inter3), .O(gate96inter10));
  nor2  gate1426(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate1427(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate1428(.a(gate96inter12), .b(gate96inter1), .O(G417));
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate1149(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate1150(.a(gate100inter0), .b(s_86), .O(gate100inter1));
  and2  gate1151(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate1152(.a(s_86), .O(gate100inter3));
  inv1  gate1153(.a(s_87), .O(gate100inter4));
  nand2 gate1154(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate1155(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate1156(.a(G31), .O(gate100inter7));
  inv1  gate1157(.a(G353), .O(gate100inter8));
  nand2 gate1158(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate1159(.a(s_87), .b(gate100inter3), .O(gate100inter10));
  nor2  gate1160(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate1161(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate1162(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );

  xor2  gate1471(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate1472(.a(gate113inter0), .b(s_132), .O(gate113inter1));
  and2  gate1473(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate1474(.a(s_132), .O(gate113inter3));
  inv1  gate1475(.a(s_133), .O(gate113inter4));
  nand2 gate1476(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate1477(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate1478(.a(G378), .O(gate113inter7));
  inv1  gate1479(.a(G379), .O(gate113inter8));
  nand2 gate1480(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate1481(.a(s_133), .b(gate113inter3), .O(gate113inter10));
  nor2  gate1482(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate1483(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate1484(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );

  xor2  gate1261(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate1262(.a(gate122inter0), .b(s_102), .O(gate122inter1));
  and2  gate1263(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate1264(.a(s_102), .O(gate122inter3));
  inv1  gate1265(.a(s_103), .O(gate122inter4));
  nand2 gate1266(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate1267(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate1268(.a(G396), .O(gate122inter7));
  inv1  gate1269(.a(G397), .O(gate122inter8));
  nand2 gate1270(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate1271(.a(s_103), .b(gate122inter3), .O(gate122inter10));
  nor2  gate1272(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate1273(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate1274(.a(gate122inter12), .b(gate122inter1), .O(G477));
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate785(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate786(.a(gate131inter0), .b(s_34), .O(gate131inter1));
  and2  gate787(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate788(.a(s_34), .O(gate131inter3));
  inv1  gate789(.a(s_35), .O(gate131inter4));
  nand2 gate790(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate791(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate792(.a(G414), .O(gate131inter7));
  inv1  gate793(.a(G415), .O(gate131inter8));
  nand2 gate794(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate795(.a(s_35), .b(gate131inter3), .O(gate131inter10));
  nor2  gate796(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate797(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate798(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate1079(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate1080(.a(gate135inter0), .b(s_76), .O(gate135inter1));
  and2  gate1081(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate1082(.a(s_76), .O(gate135inter3));
  inv1  gate1083(.a(s_77), .O(gate135inter4));
  nand2 gate1084(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate1085(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate1086(.a(G422), .O(gate135inter7));
  inv1  gate1087(.a(G423), .O(gate135inter8));
  nand2 gate1088(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate1089(.a(s_77), .b(gate135inter3), .O(gate135inter10));
  nor2  gate1090(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate1091(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate1092(.a(gate135inter12), .b(gate135inter1), .O(G516));
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate1639(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1640(.a(gate148inter0), .b(s_156), .O(gate148inter1));
  and2  gate1641(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1642(.a(s_156), .O(gate148inter3));
  inv1  gate1643(.a(s_157), .O(gate148inter4));
  nand2 gate1644(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1645(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1646(.a(G492), .O(gate148inter7));
  inv1  gate1647(.a(G495), .O(gate148inter8));
  nand2 gate1648(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1649(.a(s_157), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1650(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1651(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1652(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate897(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate898(.a(gate151inter0), .b(s_50), .O(gate151inter1));
  and2  gate899(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate900(.a(s_50), .O(gate151inter3));
  inv1  gate901(.a(s_51), .O(gate151inter4));
  nand2 gate902(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate903(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate904(.a(G510), .O(gate151inter7));
  inv1  gate905(.a(G513), .O(gate151inter8));
  nand2 gate906(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate907(.a(s_51), .b(gate151inter3), .O(gate151inter10));
  nor2  gate908(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate909(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate910(.a(gate151inter12), .b(gate151inter1), .O(G564));

  xor2  gate1387(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate1388(.a(gate152inter0), .b(s_120), .O(gate152inter1));
  and2  gate1389(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate1390(.a(s_120), .O(gate152inter3));
  inv1  gate1391(.a(s_121), .O(gate152inter4));
  nand2 gate1392(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate1393(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate1394(.a(G516), .O(gate152inter7));
  inv1  gate1395(.a(G519), .O(gate152inter8));
  nand2 gate1396(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate1397(.a(s_121), .b(gate152inter3), .O(gate152inter10));
  nor2  gate1398(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate1399(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate1400(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate1723(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate1724(.a(gate157inter0), .b(s_168), .O(gate157inter1));
  and2  gate1725(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate1726(.a(s_168), .O(gate157inter3));
  inv1  gate1727(.a(s_169), .O(gate157inter4));
  nand2 gate1728(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate1729(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate1730(.a(G438), .O(gate157inter7));
  inv1  gate1731(.a(G528), .O(gate157inter8));
  nand2 gate1732(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate1733(.a(s_169), .b(gate157inter3), .O(gate157inter10));
  nor2  gate1734(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate1735(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate1736(.a(gate157inter12), .b(gate157inter1), .O(G574));

  xor2  gate995(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate996(.a(gate158inter0), .b(s_64), .O(gate158inter1));
  and2  gate997(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate998(.a(s_64), .O(gate158inter3));
  inv1  gate999(.a(s_65), .O(gate158inter4));
  nand2 gate1000(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate1001(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate1002(.a(G441), .O(gate158inter7));
  inv1  gate1003(.a(G528), .O(gate158inter8));
  nand2 gate1004(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate1005(.a(s_65), .b(gate158inter3), .O(gate158inter10));
  nor2  gate1006(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate1007(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate1008(.a(gate158inter12), .b(gate158inter1), .O(G575));

  xor2  gate757(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate758(.a(gate159inter0), .b(s_30), .O(gate159inter1));
  and2  gate759(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate760(.a(s_30), .O(gate159inter3));
  inv1  gate761(.a(s_31), .O(gate159inter4));
  nand2 gate762(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate763(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate764(.a(G444), .O(gate159inter7));
  inv1  gate765(.a(G531), .O(gate159inter8));
  nand2 gate766(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate767(.a(s_31), .b(gate159inter3), .O(gate159inter10));
  nor2  gate768(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate769(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate770(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate1205(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate1206(.a(gate161inter0), .b(s_94), .O(gate161inter1));
  and2  gate1207(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate1208(.a(s_94), .O(gate161inter3));
  inv1  gate1209(.a(s_95), .O(gate161inter4));
  nand2 gate1210(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate1211(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate1212(.a(G450), .O(gate161inter7));
  inv1  gate1213(.a(G534), .O(gate161inter8));
  nand2 gate1214(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate1215(.a(s_95), .b(gate161inter3), .O(gate161inter10));
  nor2  gate1216(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate1217(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate1218(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate561(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate562(.a(gate165inter0), .b(s_2), .O(gate165inter1));
  and2  gate563(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate564(.a(s_2), .O(gate165inter3));
  inv1  gate565(.a(s_3), .O(gate165inter4));
  nand2 gate566(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate567(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate568(.a(G462), .O(gate165inter7));
  inv1  gate569(.a(G540), .O(gate165inter8));
  nand2 gate570(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate571(.a(s_3), .b(gate165inter3), .O(gate165inter10));
  nor2  gate572(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate573(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate574(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );

  xor2  gate589(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate590(.a(gate177inter0), .b(s_6), .O(gate177inter1));
  and2  gate591(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate592(.a(s_6), .O(gate177inter3));
  inv1  gate593(.a(s_7), .O(gate177inter4));
  nand2 gate594(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate595(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate596(.a(G498), .O(gate177inter7));
  inv1  gate597(.a(G558), .O(gate177inter8));
  nand2 gate598(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate599(.a(s_7), .b(gate177inter3), .O(gate177inter10));
  nor2  gate600(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate601(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate602(.a(gate177inter12), .b(gate177inter1), .O(G594));

  xor2  gate1527(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate1528(.a(gate178inter0), .b(s_140), .O(gate178inter1));
  and2  gate1529(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate1530(.a(s_140), .O(gate178inter3));
  inv1  gate1531(.a(s_141), .O(gate178inter4));
  nand2 gate1532(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate1533(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate1534(.a(G501), .O(gate178inter7));
  inv1  gate1535(.a(G558), .O(gate178inter8));
  nand2 gate1536(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate1537(.a(s_141), .b(gate178inter3), .O(gate178inter10));
  nor2  gate1538(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate1539(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate1540(.a(gate178inter12), .b(gate178inter1), .O(G595));
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate841(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate842(.a(gate181inter0), .b(s_42), .O(gate181inter1));
  and2  gate843(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate844(.a(s_42), .O(gate181inter3));
  inv1  gate845(.a(s_43), .O(gate181inter4));
  nand2 gate846(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate847(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate848(.a(G510), .O(gate181inter7));
  inv1  gate849(.a(G564), .O(gate181inter8));
  nand2 gate850(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate851(.a(s_43), .b(gate181inter3), .O(gate181inter10));
  nor2  gate852(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate853(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate854(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate1303(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate1304(.a(gate184inter0), .b(s_108), .O(gate184inter1));
  and2  gate1305(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate1306(.a(s_108), .O(gate184inter3));
  inv1  gate1307(.a(s_109), .O(gate184inter4));
  nand2 gate1308(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate1309(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate1310(.a(G519), .O(gate184inter7));
  inv1  gate1311(.a(G567), .O(gate184inter8));
  nand2 gate1312(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate1313(.a(s_109), .b(gate184inter3), .O(gate184inter10));
  nor2  gate1314(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate1315(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate1316(.a(gate184inter12), .b(gate184inter1), .O(G601));

  xor2  gate939(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate940(.a(gate185inter0), .b(s_56), .O(gate185inter1));
  and2  gate941(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate942(.a(s_56), .O(gate185inter3));
  inv1  gate943(.a(s_57), .O(gate185inter4));
  nand2 gate944(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate945(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate946(.a(G570), .O(gate185inter7));
  inv1  gate947(.a(G571), .O(gate185inter8));
  nand2 gate948(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate949(.a(s_57), .b(gate185inter3), .O(gate185inter10));
  nor2  gate950(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate951(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate952(.a(gate185inter12), .b(gate185inter1), .O(G602));
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate1177(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate1178(.a(gate188inter0), .b(s_90), .O(gate188inter1));
  and2  gate1179(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate1180(.a(s_90), .O(gate188inter3));
  inv1  gate1181(.a(s_91), .O(gate188inter4));
  nand2 gate1182(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate1183(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate1184(.a(G576), .O(gate188inter7));
  inv1  gate1185(.a(G577), .O(gate188inter8));
  nand2 gate1186(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate1187(.a(s_91), .b(gate188inter3), .O(gate188inter10));
  nor2  gate1188(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate1189(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate1190(.a(gate188inter12), .b(gate188inter1), .O(G617));

  xor2  gate1233(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate1234(.a(gate189inter0), .b(s_98), .O(gate189inter1));
  and2  gate1235(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate1236(.a(s_98), .O(gate189inter3));
  inv1  gate1237(.a(s_99), .O(gate189inter4));
  nand2 gate1238(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate1239(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate1240(.a(G578), .O(gate189inter7));
  inv1  gate1241(.a(G579), .O(gate189inter8));
  nand2 gate1242(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate1243(.a(s_99), .b(gate189inter3), .O(gate189inter10));
  nor2  gate1244(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate1245(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate1246(.a(gate189inter12), .b(gate189inter1), .O(G622));
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );

  xor2  gate813(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate814(.a(gate192inter0), .b(s_38), .O(gate192inter1));
  and2  gate815(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate816(.a(s_38), .O(gate192inter3));
  inv1  gate817(.a(s_39), .O(gate192inter4));
  nand2 gate818(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate819(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate820(.a(G584), .O(gate192inter7));
  inv1  gate821(.a(G585), .O(gate192inter8));
  nand2 gate822(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate823(.a(s_39), .b(gate192inter3), .O(gate192inter10));
  nor2  gate824(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate825(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate826(.a(gate192inter12), .b(gate192inter1), .O(G637));

  xor2  gate729(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate730(.a(gate193inter0), .b(s_26), .O(gate193inter1));
  and2  gate731(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate732(.a(s_26), .O(gate193inter3));
  inv1  gate733(.a(s_27), .O(gate193inter4));
  nand2 gate734(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate735(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate736(.a(G586), .O(gate193inter7));
  inv1  gate737(.a(G587), .O(gate193inter8));
  nand2 gate738(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate739(.a(s_27), .b(gate193inter3), .O(gate193inter10));
  nor2  gate740(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate741(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate742(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate981(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate982(.a(gate195inter0), .b(s_62), .O(gate195inter1));
  and2  gate983(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate984(.a(s_62), .O(gate195inter3));
  inv1  gate985(.a(s_63), .O(gate195inter4));
  nand2 gate986(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate987(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate988(.a(G590), .O(gate195inter7));
  inv1  gate989(.a(G591), .O(gate195inter8));
  nand2 gate990(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate991(.a(s_63), .b(gate195inter3), .O(gate195inter10));
  nor2  gate992(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate993(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate994(.a(gate195inter12), .b(gate195inter1), .O(G648));

  xor2  gate953(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate954(.a(gate196inter0), .b(s_58), .O(gate196inter1));
  and2  gate955(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate956(.a(s_58), .O(gate196inter3));
  inv1  gate957(.a(s_59), .O(gate196inter4));
  nand2 gate958(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate959(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate960(.a(G592), .O(gate196inter7));
  inv1  gate961(.a(G593), .O(gate196inter8));
  nand2 gate962(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate963(.a(s_59), .b(gate196inter3), .O(gate196inter10));
  nor2  gate964(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate965(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate966(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );

  xor2  gate1121(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate1122(.a(gate199inter0), .b(s_82), .O(gate199inter1));
  and2  gate1123(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate1124(.a(s_82), .O(gate199inter3));
  inv1  gate1125(.a(s_83), .O(gate199inter4));
  nand2 gate1126(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate1127(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate1128(.a(G598), .O(gate199inter7));
  inv1  gate1129(.a(G599), .O(gate199inter8));
  nand2 gate1130(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate1131(.a(s_83), .b(gate199inter3), .O(gate199inter10));
  nor2  gate1132(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate1133(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate1134(.a(gate199inter12), .b(gate199inter1), .O(G660));

  xor2  gate1541(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate1542(.a(gate200inter0), .b(s_142), .O(gate200inter1));
  and2  gate1543(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate1544(.a(s_142), .O(gate200inter3));
  inv1  gate1545(.a(s_143), .O(gate200inter4));
  nand2 gate1546(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate1547(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate1548(.a(G600), .O(gate200inter7));
  inv1  gate1549(.a(G601), .O(gate200inter8));
  nand2 gate1550(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate1551(.a(s_143), .b(gate200inter3), .O(gate200inter10));
  nor2  gate1552(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate1553(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate1554(.a(gate200inter12), .b(gate200inter1), .O(G663));
nand2 gate201( .a(G602), .b(G607), .O(G666) );

  xor2  gate1331(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate1332(.a(gate202inter0), .b(s_112), .O(gate202inter1));
  and2  gate1333(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate1334(.a(s_112), .O(gate202inter3));
  inv1  gate1335(.a(s_113), .O(gate202inter4));
  nand2 gate1336(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate1337(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate1338(.a(G612), .O(gate202inter7));
  inv1  gate1339(.a(G617), .O(gate202inter8));
  nand2 gate1340(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate1341(.a(s_113), .b(gate202inter3), .O(gate202inter10));
  nor2  gate1342(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate1343(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate1344(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate1779(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate1780(.a(gate206inter0), .b(s_176), .O(gate206inter1));
  and2  gate1781(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate1782(.a(s_176), .O(gate206inter3));
  inv1  gate1783(.a(s_177), .O(gate206inter4));
  nand2 gate1784(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate1785(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate1786(.a(G632), .O(gate206inter7));
  inv1  gate1787(.a(G637), .O(gate206inter8));
  nand2 gate1788(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate1789(.a(s_177), .b(gate206inter3), .O(gate206inter10));
  nor2  gate1790(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate1791(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate1792(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate1163(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate1164(.a(gate211inter0), .b(s_88), .O(gate211inter1));
  and2  gate1165(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate1166(.a(s_88), .O(gate211inter3));
  inv1  gate1167(.a(s_89), .O(gate211inter4));
  nand2 gate1168(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate1169(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate1170(.a(G612), .O(gate211inter7));
  inv1  gate1171(.a(G669), .O(gate211inter8));
  nand2 gate1172(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate1173(.a(s_89), .b(gate211inter3), .O(gate211inter10));
  nor2  gate1174(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate1175(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate1176(.a(gate211inter12), .b(gate211inter1), .O(G692));
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate1317(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate1318(.a(gate213inter0), .b(s_110), .O(gate213inter1));
  and2  gate1319(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate1320(.a(s_110), .O(gate213inter3));
  inv1  gate1321(.a(s_111), .O(gate213inter4));
  nand2 gate1322(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate1323(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate1324(.a(G602), .O(gate213inter7));
  inv1  gate1325(.a(G672), .O(gate213inter8));
  nand2 gate1326(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate1327(.a(s_111), .b(gate213inter3), .O(gate213inter10));
  nor2  gate1328(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate1329(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate1330(.a(gate213inter12), .b(gate213inter1), .O(G694));

  xor2  gate1135(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate1136(.a(gate214inter0), .b(s_84), .O(gate214inter1));
  and2  gate1137(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate1138(.a(s_84), .O(gate214inter3));
  inv1  gate1139(.a(s_85), .O(gate214inter4));
  nand2 gate1140(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate1141(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate1142(.a(G612), .O(gate214inter7));
  inv1  gate1143(.a(G672), .O(gate214inter8));
  nand2 gate1144(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate1145(.a(s_85), .b(gate214inter3), .O(gate214inter10));
  nor2  gate1146(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate1147(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate1148(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate883(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate884(.a(gate219inter0), .b(s_48), .O(gate219inter1));
  and2  gate885(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate886(.a(s_48), .O(gate219inter3));
  inv1  gate887(.a(s_49), .O(gate219inter4));
  nand2 gate888(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate889(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate890(.a(G632), .O(gate219inter7));
  inv1  gate891(.a(G681), .O(gate219inter8));
  nand2 gate892(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate893(.a(s_49), .b(gate219inter3), .O(gate219inter10));
  nor2  gate894(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate895(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate896(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate1583(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate1584(.a(gate234inter0), .b(s_148), .O(gate234inter1));
  and2  gate1585(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate1586(.a(s_148), .O(gate234inter3));
  inv1  gate1587(.a(s_149), .O(gate234inter4));
  nand2 gate1588(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1589(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1590(.a(G245), .O(gate234inter7));
  inv1  gate1591(.a(G721), .O(gate234inter8));
  nand2 gate1592(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1593(.a(s_149), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1594(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1595(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1596(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );

  xor2  gate1247(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate1248(.a(gate238inter0), .b(s_100), .O(gate238inter1));
  and2  gate1249(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate1250(.a(s_100), .O(gate238inter3));
  inv1  gate1251(.a(s_101), .O(gate238inter4));
  nand2 gate1252(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate1253(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate1254(.a(G257), .O(gate238inter7));
  inv1  gate1255(.a(G709), .O(gate238inter8));
  nand2 gate1256(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate1257(.a(s_101), .b(gate238inter3), .O(gate238inter10));
  nor2  gate1258(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate1259(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate1260(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate827(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate828(.a(gate248inter0), .b(s_40), .O(gate248inter1));
  and2  gate829(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate830(.a(s_40), .O(gate248inter3));
  inv1  gate831(.a(s_41), .O(gate248inter4));
  nand2 gate832(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate833(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate834(.a(G727), .O(gate248inter7));
  inv1  gate835(.a(G739), .O(gate248inter8));
  nand2 gate836(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate837(.a(s_41), .b(gate248inter3), .O(gate248inter10));
  nor2  gate838(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate839(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate840(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );

  xor2  gate911(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate912(.a(gate251inter0), .b(s_52), .O(gate251inter1));
  and2  gate913(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate914(.a(s_52), .O(gate251inter3));
  inv1  gate915(.a(s_53), .O(gate251inter4));
  nand2 gate916(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate917(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate918(.a(G257), .O(gate251inter7));
  inv1  gate919(.a(G745), .O(gate251inter8));
  nand2 gate920(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate921(.a(s_53), .b(gate251inter3), .O(gate251inter10));
  nor2  gate922(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate923(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate924(.a(gate251inter12), .b(gate251inter1), .O(G764));
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );

  xor2  gate631(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate632(.a(gate260inter0), .b(s_12), .O(gate260inter1));
  and2  gate633(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate634(.a(s_12), .O(gate260inter3));
  inv1  gate635(.a(s_13), .O(gate260inter4));
  nand2 gate636(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate637(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate638(.a(G760), .O(gate260inter7));
  inv1  gate639(.a(G761), .O(gate260inter8));
  nand2 gate640(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate641(.a(s_13), .b(gate260inter3), .O(gate260inter10));
  nor2  gate642(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate643(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate644(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate1191(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate1192(.a(gate262inter0), .b(s_92), .O(gate262inter1));
  and2  gate1193(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate1194(.a(s_92), .O(gate262inter3));
  inv1  gate1195(.a(s_93), .O(gate262inter4));
  nand2 gate1196(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate1197(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate1198(.a(G764), .O(gate262inter7));
  inv1  gate1199(.a(G765), .O(gate262inter8));
  nand2 gate1200(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate1201(.a(s_93), .b(gate262inter3), .O(gate262inter10));
  nor2  gate1202(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate1203(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate1204(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate743(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate744(.a(gate270inter0), .b(s_28), .O(gate270inter1));
  and2  gate745(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate746(.a(s_28), .O(gate270inter3));
  inv1  gate747(.a(s_29), .O(gate270inter4));
  nand2 gate748(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate749(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate750(.a(G657), .O(gate270inter7));
  inv1  gate751(.a(G785), .O(gate270inter8));
  nand2 gate752(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate753(.a(s_29), .b(gate270inter3), .O(gate270inter10));
  nor2  gate754(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate755(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate756(.a(gate270inter12), .b(gate270inter1), .O(G809));
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );

  xor2  gate1401(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate1402(.a(gate273inter0), .b(s_122), .O(gate273inter1));
  and2  gate1403(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate1404(.a(s_122), .O(gate273inter3));
  inv1  gate1405(.a(s_123), .O(gate273inter4));
  nand2 gate1406(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate1407(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate1408(.a(G642), .O(gate273inter7));
  inv1  gate1409(.a(G794), .O(gate273inter8));
  nand2 gate1410(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate1411(.a(s_123), .b(gate273inter3), .O(gate273inter10));
  nor2  gate1412(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate1413(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate1414(.a(gate273inter12), .b(gate273inter1), .O(G818));
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate1667(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate1668(.a(gate278inter0), .b(s_160), .O(gate278inter1));
  and2  gate1669(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate1670(.a(s_160), .O(gate278inter3));
  inv1  gate1671(.a(s_161), .O(gate278inter4));
  nand2 gate1672(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate1673(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate1674(.a(G776), .O(gate278inter7));
  inv1  gate1675(.a(G800), .O(gate278inter8));
  nand2 gate1676(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate1677(.a(s_161), .b(gate278inter3), .O(gate278inter10));
  nor2  gate1678(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate1679(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate1680(.a(gate278inter12), .b(gate278inter1), .O(G823));

  xor2  gate1597(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate1598(.a(gate279inter0), .b(s_150), .O(gate279inter1));
  and2  gate1599(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate1600(.a(s_150), .O(gate279inter3));
  inv1  gate1601(.a(s_151), .O(gate279inter4));
  nand2 gate1602(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate1603(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate1604(.a(G651), .O(gate279inter7));
  inv1  gate1605(.a(G803), .O(gate279inter8));
  nand2 gate1606(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate1607(.a(s_151), .b(gate279inter3), .O(gate279inter10));
  nor2  gate1608(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate1609(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate1610(.a(gate279inter12), .b(gate279inter1), .O(G824));

  xor2  gate799(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate800(.a(gate280inter0), .b(s_36), .O(gate280inter1));
  and2  gate801(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate802(.a(s_36), .O(gate280inter3));
  inv1  gate803(.a(s_37), .O(gate280inter4));
  nand2 gate804(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate805(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate806(.a(G779), .O(gate280inter7));
  inv1  gate807(.a(G803), .O(gate280inter8));
  nand2 gate808(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate809(.a(s_37), .b(gate280inter3), .O(gate280inter10));
  nor2  gate810(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate811(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate812(.a(gate280inter12), .b(gate280inter1), .O(G825));

  xor2  gate659(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate660(.a(gate281inter0), .b(s_16), .O(gate281inter1));
  and2  gate661(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate662(.a(s_16), .O(gate281inter3));
  inv1  gate663(.a(s_17), .O(gate281inter4));
  nand2 gate664(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate665(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate666(.a(G654), .O(gate281inter7));
  inv1  gate667(.a(G806), .O(gate281inter8));
  nand2 gate668(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate669(.a(s_17), .b(gate281inter3), .O(gate281inter10));
  nor2  gate670(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate671(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate672(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate645(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate646(.a(gate283inter0), .b(s_14), .O(gate283inter1));
  and2  gate647(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate648(.a(s_14), .O(gate283inter3));
  inv1  gate649(.a(s_15), .O(gate283inter4));
  nand2 gate650(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate651(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate652(.a(G657), .O(gate283inter7));
  inv1  gate653(.a(G809), .O(gate283inter8));
  nand2 gate654(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate655(.a(s_15), .b(gate283inter3), .O(gate283inter10));
  nor2  gate656(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate657(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate658(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate1023(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate1024(.a(gate290inter0), .b(s_68), .O(gate290inter1));
  and2  gate1025(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate1026(.a(s_68), .O(gate290inter3));
  inv1  gate1027(.a(s_69), .O(gate290inter4));
  nand2 gate1028(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate1029(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate1030(.a(G820), .O(gate290inter7));
  inv1  gate1031(.a(G821), .O(gate290inter8));
  nand2 gate1032(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate1033(.a(s_69), .b(gate290inter3), .O(gate290inter10));
  nor2  gate1034(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate1035(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate1036(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate1373(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate1374(.a(gate393inter0), .b(s_118), .O(gate393inter1));
  and2  gate1375(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate1376(.a(s_118), .O(gate393inter3));
  inv1  gate1377(.a(s_119), .O(gate393inter4));
  nand2 gate1378(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate1379(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate1380(.a(G7), .O(gate393inter7));
  inv1  gate1381(.a(G1054), .O(gate393inter8));
  nand2 gate1382(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate1383(.a(s_119), .b(gate393inter3), .O(gate393inter10));
  nor2  gate1384(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate1385(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate1386(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );

  xor2  gate1443(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate1444(.a(gate401inter0), .b(s_128), .O(gate401inter1));
  and2  gate1445(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate1446(.a(s_128), .O(gate401inter3));
  inv1  gate1447(.a(s_129), .O(gate401inter4));
  nand2 gate1448(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate1449(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate1450(.a(G15), .O(gate401inter7));
  inv1  gate1451(.a(G1078), .O(gate401inter8));
  nand2 gate1452(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate1453(.a(s_129), .b(gate401inter3), .O(gate401inter10));
  nor2  gate1454(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate1455(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate1456(.a(gate401inter12), .b(gate401inter1), .O(G1174));

  xor2  gate869(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate870(.a(gate402inter0), .b(s_46), .O(gate402inter1));
  and2  gate871(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate872(.a(s_46), .O(gate402inter3));
  inv1  gate873(.a(s_47), .O(gate402inter4));
  nand2 gate874(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate875(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate876(.a(G16), .O(gate402inter7));
  inv1  gate877(.a(G1081), .O(gate402inter8));
  nand2 gate878(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate879(.a(s_47), .b(gate402inter3), .O(gate402inter10));
  nor2  gate880(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate881(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate882(.a(gate402inter12), .b(gate402inter1), .O(G1177));
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate1611(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate1612(.a(gate415inter0), .b(s_152), .O(gate415inter1));
  and2  gate1613(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate1614(.a(s_152), .O(gate415inter3));
  inv1  gate1615(.a(s_153), .O(gate415inter4));
  nand2 gate1616(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate1617(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate1618(.a(G29), .O(gate415inter7));
  inv1  gate1619(.a(G1120), .O(gate415inter8));
  nand2 gate1620(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate1621(.a(s_153), .b(gate415inter3), .O(gate415inter10));
  nor2  gate1622(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate1623(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate1624(.a(gate415inter12), .b(gate415inter1), .O(G1216));

  xor2  gate1681(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate1682(.a(gate416inter0), .b(s_162), .O(gate416inter1));
  and2  gate1683(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate1684(.a(s_162), .O(gate416inter3));
  inv1  gate1685(.a(s_163), .O(gate416inter4));
  nand2 gate1686(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate1687(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate1688(.a(G30), .O(gate416inter7));
  inv1  gate1689(.a(G1123), .O(gate416inter8));
  nand2 gate1690(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate1691(.a(s_163), .b(gate416inter3), .O(gate416inter10));
  nor2  gate1692(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate1693(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate1694(.a(gate416inter12), .b(gate416inter1), .O(G1219));
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );

  xor2  gate1737(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate1738(.a(gate426inter0), .b(s_170), .O(gate426inter1));
  and2  gate1739(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate1740(.a(s_170), .O(gate426inter3));
  inv1  gate1741(.a(s_171), .O(gate426inter4));
  nand2 gate1742(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate1743(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate1744(.a(G1045), .O(gate426inter7));
  inv1  gate1745(.a(G1141), .O(gate426inter8));
  nand2 gate1746(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate1747(.a(s_171), .b(gate426inter3), .O(gate426inter10));
  nor2  gate1748(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate1749(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate1750(.a(gate426inter12), .b(gate426inter1), .O(G1235));

  xor2  gate1793(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate1794(.a(gate427inter0), .b(s_178), .O(gate427inter1));
  and2  gate1795(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate1796(.a(s_178), .O(gate427inter3));
  inv1  gate1797(.a(s_179), .O(gate427inter4));
  nand2 gate1798(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate1799(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate1800(.a(G5), .O(gate427inter7));
  inv1  gate1801(.a(G1144), .O(gate427inter8));
  nand2 gate1802(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate1803(.a(s_179), .b(gate427inter3), .O(gate427inter10));
  nor2  gate1804(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate1805(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate1806(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );

  xor2  gate617(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate618(.a(gate429inter0), .b(s_10), .O(gate429inter1));
  and2  gate619(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate620(.a(s_10), .O(gate429inter3));
  inv1  gate621(.a(s_11), .O(gate429inter4));
  nand2 gate622(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate623(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate624(.a(G6), .O(gate429inter7));
  inv1  gate625(.a(G1147), .O(gate429inter8));
  nand2 gate626(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate627(.a(s_11), .b(gate429inter3), .O(gate429inter10));
  nor2  gate628(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate629(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate630(.a(gate429inter12), .b(gate429inter1), .O(G1238));
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate1807(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate1808(.a(gate433inter0), .b(s_180), .O(gate433inter1));
  and2  gate1809(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate1810(.a(s_180), .O(gate433inter3));
  inv1  gate1811(.a(s_181), .O(gate433inter4));
  nand2 gate1812(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate1813(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate1814(.a(G8), .O(gate433inter7));
  inv1  gate1815(.a(G1153), .O(gate433inter8));
  nand2 gate1816(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate1817(.a(s_181), .b(gate433inter3), .O(gate433inter10));
  nor2  gate1818(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate1819(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate1820(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate1051(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate1052(.a(gate441inter0), .b(s_72), .O(gate441inter1));
  and2  gate1053(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate1054(.a(s_72), .O(gate441inter3));
  inv1  gate1055(.a(s_73), .O(gate441inter4));
  nand2 gate1056(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate1057(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate1058(.a(G12), .O(gate441inter7));
  inv1  gate1059(.a(G1165), .O(gate441inter8));
  nand2 gate1060(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate1061(.a(s_73), .b(gate441inter3), .O(gate441inter10));
  nor2  gate1062(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate1063(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate1064(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate1485(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate1486(.a(gate444inter0), .b(s_134), .O(gate444inter1));
  and2  gate1487(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate1488(.a(s_134), .O(gate444inter3));
  inv1  gate1489(.a(s_135), .O(gate444inter4));
  nand2 gate1490(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate1491(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate1492(.a(G1072), .O(gate444inter7));
  inv1  gate1493(.a(G1168), .O(gate444inter8));
  nand2 gate1494(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate1495(.a(s_135), .b(gate444inter3), .O(gate444inter10));
  nor2  gate1496(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate1497(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate1498(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );

  xor2  gate1037(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate1038(.a(gate450inter0), .b(s_70), .O(gate450inter1));
  and2  gate1039(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate1040(.a(s_70), .O(gate450inter3));
  inv1  gate1041(.a(s_71), .O(gate450inter4));
  nand2 gate1042(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate1043(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate1044(.a(G1081), .O(gate450inter7));
  inv1  gate1045(.a(G1177), .O(gate450inter8));
  nand2 gate1046(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate1047(.a(s_71), .b(gate450inter3), .O(gate450inter10));
  nor2  gate1048(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate1049(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate1050(.a(gate450inter12), .b(gate450inter1), .O(G1259));
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );

  xor2  gate687(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate688(.a(gate452inter0), .b(s_20), .O(gate452inter1));
  and2  gate689(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate690(.a(s_20), .O(gate452inter3));
  inv1  gate691(.a(s_21), .O(gate452inter4));
  nand2 gate692(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate693(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate694(.a(G1084), .O(gate452inter7));
  inv1  gate695(.a(G1180), .O(gate452inter8));
  nand2 gate696(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate697(.a(s_21), .b(gate452inter3), .O(gate452inter10));
  nor2  gate698(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate699(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate700(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );

  xor2  gate1457(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate1458(.a(gate454inter0), .b(s_130), .O(gate454inter1));
  and2  gate1459(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate1460(.a(s_130), .O(gate454inter3));
  inv1  gate1461(.a(s_131), .O(gate454inter4));
  nand2 gate1462(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate1463(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate1464(.a(G1087), .O(gate454inter7));
  inv1  gate1465(.a(G1183), .O(gate454inter8));
  nand2 gate1466(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate1467(.a(s_131), .b(gate454inter3), .O(gate454inter10));
  nor2  gate1468(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate1469(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate1470(.a(gate454inter12), .b(gate454inter1), .O(G1263));
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate701(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate702(.a(gate456inter0), .b(s_22), .O(gate456inter1));
  and2  gate703(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate704(.a(s_22), .O(gate456inter3));
  inv1  gate705(.a(s_23), .O(gate456inter4));
  nand2 gate706(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate707(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate708(.a(G1090), .O(gate456inter7));
  inv1  gate709(.a(G1186), .O(gate456inter8));
  nand2 gate710(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate711(.a(s_23), .b(gate456inter3), .O(gate456inter10));
  nor2  gate712(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate713(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate714(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate1275(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate1276(.a(gate459inter0), .b(s_104), .O(gate459inter1));
  and2  gate1277(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate1278(.a(s_104), .O(gate459inter3));
  inv1  gate1279(.a(s_105), .O(gate459inter4));
  nand2 gate1280(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate1281(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate1282(.a(G21), .O(gate459inter7));
  inv1  gate1283(.a(G1192), .O(gate459inter8));
  nand2 gate1284(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate1285(.a(s_105), .b(gate459inter3), .O(gate459inter10));
  nor2  gate1286(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate1287(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate1288(.a(gate459inter12), .b(gate459inter1), .O(G1268));

  xor2  gate1653(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate1654(.a(gate460inter0), .b(s_158), .O(gate460inter1));
  and2  gate1655(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate1656(.a(s_158), .O(gate460inter3));
  inv1  gate1657(.a(s_159), .O(gate460inter4));
  nand2 gate1658(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate1659(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate1660(.a(G1096), .O(gate460inter7));
  inv1  gate1661(.a(G1192), .O(gate460inter8));
  nand2 gate1662(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate1663(.a(s_159), .b(gate460inter3), .O(gate460inter10));
  nor2  gate1664(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate1665(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate1666(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate1555(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate1556(.a(gate463inter0), .b(s_144), .O(gate463inter1));
  and2  gate1557(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate1558(.a(s_144), .O(gate463inter3));
  inv1  gate1559(.a(s_145), .O(gate463inter4));
  nand2 gate1560(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate1561(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate1562(.a(G23), .O(gate463inter7));
  inv1  gate1563(.a(G1198), .O(gate463inter8));
  nand2 gate1564(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate1565(.a(s_145), .b(gate463inter3), .O(gate463inter10));
  nor2  gate1566(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate1567(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate1568(.a(gate463inter12), .b(gate463inter1), .O(G1272));

  xor2  gate1513(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate1514(.a(gate464inter0), .b(s_138), .O(gate464inter1));
  and2  gate1515(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate1516(.a(s_138), .O(gate464inter3));
  inv1  gate1517(.a(s_139), .O(gate464inter4));
  nand2 gate1518(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate1519(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate1520(.a(G1102), .O(gate464inter7));
  inv1  gate1521(.a(G1198), .O(gate464inter8));
  nand2 gate1522(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate1523(.a(s_139), .b(gate464inter3), .O(gate464inter10));
  nor2  gate1524(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate1525(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate1526(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate1093(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate1094(.a(gate480inter0), .b(s_78), .O(gate480inter1));
  and2  gate1095(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate1096(.a(s_78), .O(gate480inter3));
  inv1  gate1097(.a(s_79), .O(gate480inter4));
  nand2 gate1098(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate1099(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate1100(.a(G1126), .O(gate480inter7));
  inv1  gate1101(.a(G1222), .O(gate480inter8));
  nand2 gate1102(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate1103(.a(s_79), .b(gate480inter3), .O(gate480inter10));
  nor2  gate1104(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate1105(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate1106(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate575(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate576(.a(gate486inter0), .b(s_4), .O(gate486inter1));
  and2  gate577(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate578(.a(s_4), .O(gate486inter3));
  inv1  gate579(.a(s_5), .O(gate486inter4));
  nand2 gate580(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate581(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate582(.a(G1234), .O(gate486inter7));
  inv1  gate583(.a(G1235), .O(gate486inter8));
  nand2 gate584(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate585(.a(s_5), .b(gate486inter3), .O(gate486inter10));
  nor2  gate586(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate587(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate588(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate547(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate548(.a(gate510inter0), .b(s_0), .O(gate510inter1));
  and2  gate549(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate550(.a(s_0), .O(gate510inter3));
  inv1  gate551(.a(s_1), .O(gate510inter4));
  nand2 gate552(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate553(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate554(.a(G1282), .O(gate510inter7));
  inv1  gate555(.a(G1283), .O(gate510inter8));
  nand2 gate556(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate557(.a(s_1), .b(gate510inter3), .O(gate510inter10));
  nor2  gate558(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate559(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate560(.a(gate510inter12), .b(gate510inter1), .O(G1319));

  xor2  gate673(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate674(.a(gate511inter0), .b(s_18), .O(gate511inter1));
  and2  gate675(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate676(.a(s_18), .O(gate511inter3));
  inv1  gate677(.a(s_19), .O(gate511inter4));
  nand2 gate678(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate679(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate680(.a(G1284), .O(gate511inter7));
  inv1  gate681(.a(G1285), .O(gate511inter8));
  nand2 gate682(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate683(.a(s_19), .b(gate511inter3), .O(gate511inter10));
  nor2  gate684(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate685(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate686(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate1709(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate1710(.a(gate514inter0), .b(s_166), .O(gate514inter1));
  and2  gate1711(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate1712(.a(s_166), .O(gate514inter3));
  inv1  gate1713(.a(s_167), .O(gate514inter4));
  nand2 gate1714(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate1715(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate1716(.a(G1290), .O(gate514inter7));
  inv1  gate1717(.a(G1291), .O(gate514inter8));
  nand2 gate1718(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate1719(.a(s_167), .b(gate514inter3), .O(gate514inter10));
  nor2  gate1720(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate1721(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate1722(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule