module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate799(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate800(.a(gate11inter0), .b(s_36), .O(gate11inter1));
  and2  gate801(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate802(.a(s_36), .O(gate11inter3));
  inv1  gate803(.a(s_37), .O(gate11inter4));
  nand2 gate804(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate805(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate806(.a(G5), .O(gate11inter7));
  inv1  gate807(.a(G6), .O(gate11inter8));
  nand2 gate808(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate809(.a(s_37), .b(gate11inter3), .O(gate11inter10));
  nor2  gate810(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate811(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate812(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate1107(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate1108(.a(gate13inter0), .b(s_80), .O(gate13inter1));
  and2  gate1109(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate1110(.a(s_80), .O(gate13inter3));
  inv1  gate1111(.a(s_81), .O(gate13inter4));
  nand2 gate1112(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate1113(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate1114(.a(G9), .O(gate13inter7));
  inv1  gate1115(.a(G10), .O(gate13inter8));
  nand2 gate1116(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate1117(.a(s_81), .b(gate13inter3), .O(gate13inter10));
  nor2  gate1118(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate1119(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate1120(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate841(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate842(.a(gate16inter0), .b(s_42), .O(gate16inter1));
  and2  gate843(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate844(.a(s_42), .O(gate16inter3));
  inv1  gate845(.a(s_43), .O(gate16inter4));
  nand2 gate846(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate847(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate848(.a(G15), .O(gate16inter7));
  inv1  gate849(.a(G16), .O(gate16inter8));
  nand2 gate850(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate851(.a(s_43), .b(gate16inter3), .O(gate16inter10));
  nor2  gate852(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate853(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate854(.a(gate16inter12), .b(gate16inter1), .O(G287));

  xor2  gate785(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate786(.a(gate17inter0), .b(s_34), .O(gate17inter1));
  and2  gate787(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate788(.a(s_34), .O(gate17inter3));
  inv1  gate789(.a(s_35), .O(gate17inter4));
  nand2 gate790(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate791(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate792(.a(G17), .O(gate17inter7));
  inv1  gate793(.a(G18), .O(gate17inter8));
  nand2 gate794(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate795(.a(s_35), .b(gate17inter3), .O(gate17inter10));
  nor2  gate796(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate797(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate798(.a(gate17inter12), .b(gate17inter1), .O(G290));

  xor2  gate1877(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate1878(.a(gate18inter0), .b(s_190), .O(gate18inter1));
  and2  gate1879(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate1880(.a(s_190), .O(gate18inter3));
  inv1  gate1881(.a(s_191), .O(gate18inter4));
  nand2 gate1882(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate1883(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate1884(.a(G19), .O(gate18inter7));
  inv1  gate1885(.a(G20), .O(gate18inter8));
  nand2 gate1886(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate1887(.a(s_191), .b(gate18inter3), .O(gate18inter10));
  nor2  gate1888(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate1889(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate1890(.a(gate18inter12), .b(gate18inter1), .O(G293));

  xor2  gate1121(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate1122(.a(gate19inter0), .b(s_82), .O(gate19inter1));
  and2  gate1123(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate1124(.a(s_82), .O(gate19inter3));
  inv1  gate1125(.a(s_83), .O(gate19inter4));
  nand2 gate1126(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate1127(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate1128(.a(G21), .O(gate19inter7));
  inv1  gate1129(.a(G22), .O(gate19inter8));
  nand2 gate1130(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate1131(.a(s_83), .b(gate19inter3), .O(gate19inter10));
  nor2  gate1132(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate1133(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate1134(.a(gate19inter12), .b(gate19inter1), .O(G296));

  xor2  gate1653(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate1654(.a(gate20inter0), .b(s_158), .O(gate20inter1));
  and2  gate1655(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate1656(.a(s_158), .O(gate20inter3));
  inv1  gate1657(.a(s_159), .O(gate20inter4));
  nand2 gate1658(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate1659(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate1660(.a(G23), .O(gate20inter7));
  inv1  gate1661(.a(G24), .O(gate20inter8));
  nand2 gate1662(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate1663(.a(s_159), .b(gate20inter3), .O(gate20inter10));
  nor2  gate1664(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate1665(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate1666(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate1583(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate1584(.a(gate23inter0), .b(s_148), .O(gate23inter1));
  and2  gate1585(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate1586(.a(s_148), .O(gate23inter3));
  inv1  gate1587(.a(s_149), .O(gate23inter4));
  nand2 gate1588(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate1589(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate1590(.a(G29), .O(gate23inter7));
  inv1  gate1591(.a(G30), .O(gate23inter8));
  nand2 gate1592(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate1593(.a(s_149), .b(gate23inter3), .O(gate23inter10));
  nor2  gate1594(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate1595(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate1596(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate925(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate926(.a(gate29inter0), .b(s_54), .O(gate29inter1));
  and2  gate927(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate928(.a(s_54), .O(gate29inter3));
  inv1  gate929(.a(s_55), .O(gate29inter4));
  nand2 gate930(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate931(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate932(.a(G3), .O(gate29inter7));
  inv1  gate933(.a(G7), .O(gate29inter8));
  nand2 gate934(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate935(.a(s_55), .b(gate29inter3), .O(gate29inter10));
  nor2  gate936(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate937(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate938(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate855(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate856(.a(gate37inter0), .b(s_44), .O(gate37inter1));
  and2  gate857(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate858(.a(s_44), .O(gate37inter3));
  inv1  gate859(.a(s_45), .O(gate37inter4));
  nand2 gate860(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate861(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate862(.a(G19), .O(gate37inter7));
  inv1  gate863(.a(G23), .O(gate37inter8));
  nand2 gate864(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate865(.a(s_45), .b(gate37inter3), .O(gate37inter10));
  nor2  gate866(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate867(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate868(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate813(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate814(.a(gate39inter0), .b(s_38), .O(gate39inter1));
  and2  gate815(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate816(.a(s_38), .O(gate39inter3));
  inv1  gate817(.a(s_39), .O(gate39inter4));
  nand2 gate818(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate819(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate820(.a(G20), .O(gate39inter7));
  inv1  gate821(.a(G24), .O(gate39inter8));
  nand2 gate822(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate823(.a(s_39), .b(gate39inter3), .O(gate39inter10));
  nor2  gate824(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate825(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate826(.a(gate39inter12), .b(gate39inter1), .O(G356));

  xor2  gate1345(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate1346(.a(gate40inter0), .b(s_114), .O(gate40inter1));
  and2  gate1347(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate1348(.a(s_114), .O(gate40inter3));
  inv1  gate1349(.a(s_115), .O(gate40inter4));
  nand2 gate1350(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate1351(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate1352(.a(G28), .O(gate40inter7));
  inv1  gate1353(.a(G32), .O(gate40inter8));
  nand2 gate1354(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate1355(.a(s_115), .b(gate40inter3), .O(gate40inter10));
  nor2  gate1356(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate1357(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate1358(.a(gate40inter12), .b(gate40inter1), .O(G359));
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate1387(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate1388(.a(gate46inter0), .b(s_120), .O(gate46inter1));
  and2  gate1389(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate1390(.a(s_120), .O(gate46inter3));
  inv1  gate1391(.a(s_121), .O(gate46inter4));
  nand2 gate1392(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate1393(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate1394(.a(G6), .O(gate46inter7));
  inv1  gate1395(.a(G272), .O(gate46inter8));
  nand2 gate1396(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate1397(.a(s_121), .b(gate46inter3), .O(gate46inter10));
  nor2  gate1398(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate1399(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate1400(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );

  xor2  gate1975(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate1976(.a(gate50inter0), .b(s_204), .O(gate50inter1));
  and2  gate1977(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate1978(.a(s_204), .O(gate50inter3));
  inv1  gate1979(.a(s_205), .O(gate50inter4));
  nand2 gate1980(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate1981(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate1982(.a(G10), .O(gate50inter7));
  inv1  gate1983(.a(G278), .O(gate50inter8));
  nand2 gate1984(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate1985(.a(s_205), .b(gate50inter3), .O(gate50inter10));
  nor2  gate1986(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate1987(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate1988(.a(gate50inter12), .b(gate50inter1), .O(G371));
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );

  xor2  gate589(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate590(.a(gate56inter0), .b(s_6), .O(gate56inter1));
  and2  gate591(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate592(.a(s_6), .O(gate56inter3));
  inv1  gate593(.a(s_7), .O(gate56inter4));
  nand2 gate594(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate595(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate596(.a(G16), .O(gate56inter7));
  inv1  gate597(.a(G287), .O(gate56inter8));
  nand2 gate598(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate599(.a(s_7), .b(gate56inter3), .O(gate56inter10));
  nor2  gate600(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate601(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate602(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate981(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate982(.a(gate59inter0), .b(s_62), .O(gate59inter1));
  and2  gate983(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate984(.a(s_62), .O(gate59inter3));
  inv1  gate985(.a(s_63), .O(gate59inter4));
  nand2 gate986(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate987(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate988(.a(G19), .O(gate59inter7));
  inv1  gate989(.a(G293), .O(gate59inter8));
  nand2 gate990(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate991(.a(s_63), .b(gate59inter3), .O(gate59inter10));
  nor2  gate992(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate993(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate994(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate1863(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate1864(.a(gate63inter0), .b(s_188), .O(gate63inter1));
  and2  gate1865(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate1866(.a(s_188), .O(gate63inter3));
  inv1  gate1867(.a(s_189), .O(gate63inter4));
  nand2 gate1868(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate1869(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate1870(.a(G23), .O(gate63inter7));
  inv1  gate1871(.a(G299), .O(gate63inter8));
  nand2 gate1872(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate1873(.a(s_189), .b(gate63inter3), .O(gate63inter10));
  nor2  gate1874(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate1875(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate1876(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate1891(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate1892(.a(gate66inter0), .b(s_192), .O(gate66inter1));
  and2  gate1893(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate1894(.a(s_192), .O(gate66inter3));
  inv1  gate1895(.a(s_193), .O(gate66inter4));
  nand2 gate1896(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate1897(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate1898(.a(G26), .O(gate66inter7));
  inv1  gate1899(.a(G302), .O(gate66inter8));
  nand2 gate1900(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate1901(.a(s_193), .b(gate66inter3), .O(gate66inter10));
  nor2  gate1902(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate1903(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate1904(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );

  xor2  gate1709(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate1710(.a(gate84inter0), .b(s_166), .O(gate84inter1));
  and2  gate1711(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate1712(.a(s_166), .O(gate84inter3));
  inv1  gate1713(.a(s_167), .O(gate84inter4));
  nand2 gate1714(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate1715(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate1716(.a(G15), .O(gate84inter7));
  inv1  gate1717(.a(G329), .O(gate84inter8));
  nand2 gate1718(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate1719(.a(s_167), .b(gate84inter3), .O(gate84inter10));
  nor2  gate1720(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate1721(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate1722(.a(gate84inter12), .b(gate84inter1), .O(G405));
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );

  xor2  gate1723(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate1724(.a(gate93inter0), .b(s_168), .O(gate93inter1));
  and2  gate1725(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate1726(.a(s_168), .O(gate93inter3));
  inv1  gate1727(.a(s_169), .O(gate93inter4));
  nand2 gate1728(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate1729(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate1730(.a(G18), .O(gate93inter7));
  inv1  gate1731(.a(G344), .O(gate93inter8));
  nand2 gate1732(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate1733(.a(s_169), .b(gate93inter3), .O(gate93inter10));
  nor2  gate1734(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate1735(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate1736(.a(gate93inter12), .b(gate93inter1), .O(G414));
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate1233(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate1234(.a(gate95inter0), .b(s_98), .O(gate95inter1));
  and2  gate1235(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate1236(.a(s_98), .O(gate95inter3));
  inv1  gate1237(.a(s_99), .O(gate95inter4));
  nand2 gate1238(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate1239(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate1240(.a(G26), .O(gate95inter7));
  inv1  gate1241(.a(G347), .O(gate95inter8));
  nand2 gate1242(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate1243(.a(s_99), .b(gate95inter3), .O(gate95inter10));
  nor2  gate1244(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate1245(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate1246(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate715(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate716(.a(gate98inter0), .b(s_24), .O(gate98inter1));
  and2  gate717(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate718(.a(s_24), .O(gate98inter3));
  inv1  gate719(.a(s_25), .O(gate98inter4));
  nand2 gate720(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate721(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate722(.a(G23), .O(gate98inter7));
  inv1  gate723(.a(G350), .O(gate98inter8));
  nand2 gate724(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate725(.a(s_25), .b(gate98inter3), .O(gate98inter10));
  nor2  gate726(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate727(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate728(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate911(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate912(.a(gate107inter0), .b(s_52), .O(gate107inter1));
  and2  gate913(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate914(.a(s_52), .O(gate107inter3));
  inv1  gate915(.a(s_53), .O(gate107inter4));
  nand2 gate916(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate917(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate918(.a(G366), .O(gate107inter7));
  inv1  gate919(.a(G367), .O(gate107inter8));
  nand2 gate920(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate921(.a(s_53), .b(gate107inter3), .O(gate107inter10));
  nor2  gate922(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate923(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate924(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );

  xor2  gate1079(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate1080(.a(gate111inter0), .b(s_76), .O(gate111inter1));
  and2  gate1081(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate1082(.a(s_76), .O(gate111inter3));
  inv1  gate1083(.a(s_77), .O(gate111inter4));
  nand2 gate1084(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate1085(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate1086(.a(G374), .O(gate111inter7));
  inv1  gate1087(.a(G375), .O(gate111inter8));
  nand2 gate1088(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate1089(.a(s_77), .b(gate111inter3), .O(gate111inter10));
  nor2  gate1090(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate1091(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate1092(.a(gate111inter12), .b(gate111inter1), .O(G444));

  xor2  gate1205(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate1206(.a(gate112inter0), .b(s_94), .O(gate112inter1));
  and2  gate1207(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate1208(.a(s_94), .O(gate112inter3));
  inv1  gate1209(.a(s_95), .O(gate112inter4));
  nand2 gate1210(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate1211(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate1212(.a(G376), .O(gate112inter7));
  inv1  gate1213(.a(G377), .O(gate112inter8));
  nand2 gate1214(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate1215(.a(s_95), .b(gate112inter3), .O(gate112inter10));
  nor2  gate1216(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate1217(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate1218(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate1023(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate1024(.a(gate115inter0), .b(s_68), .O(gate115inter1));
  and2  gate1025(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate1026(.a(s_68), .O(gate115inter3));
  inv1  gate1027(.a(s_69), .O(gate115inter4));
  nand2 gate1028(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate1029(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate1030(.a(G382), .O(gate115inter7));
  inv1  gate1031(.a(G383), .O(gate115inter8));
  nand2 gate1032(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate1033(.a(s_69), .b(gate115inter3), .O(gate115inter10));
  nor2  gate1034(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate1035(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate1036(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate1905(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate1906(.a(gate124inter0), .b(s_194), .O(gate124inter1));
  and2  gate1907(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate1908(.a(s_194), .O(gate124inter3));
  inv1  gate1909(.a(s_195), .O(gate124inter4));
  nand2 gate1910(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate1911(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate1912(.a(G400), .O(gate124inter7));
  inv1  gate1913(.a(G401), .O(gate124inter8));
  nand2 gate1914(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate1915(.a(s_195), .b(gate124inter3), .O(gate124inter10));
  nor2  gate1916(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate1917(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate1918(.a(gate124inter12), .b(gate124inter1), .O(G483));

  xor2  gate1835(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate1836(.a(gate125inter0), .b(s_184), .O(gate125inter1));
  and2  gate1837(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate1838(.a(s_184), .O(gate125inter3));
  inv1  gate1839(.a(s_185), .O(gate125inter4));
  nand2 gate1840(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate1841(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate1842(.a(G402), .O(gate125inter7));
  inv1  gate1843(.a(G403), .O(gate125inter8));
  nand2 gate1844(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate1845(.a(s_185), .b(gate125inter3), .O(gate125inter10));
  nor2  gate1846(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate1847(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate1848(.a(gate125inter12), .b(gate125inter1), .O(G486));

  xor2  gate1499(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate1500(.a(gate126inter0), .b(s_136), .O(gate126inter1));
  and2  gate1501(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate1502(.a(s_136), .O(gate126inter3));
  inv1  gate1503(.a(s_137), .O(gate126inter4));
  nand2 gate1504(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate1505(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate1506(.a(G404), .O(gate126inter7));
  inv1  gate1507(.a(G405), .O(gate126inter8));
  nand2 gate1508(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate1509(.a(s_137), .b(gate126inter3), .O(gate126inter10));
  nor2  gate1510(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate1511(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate1512(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate883(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate884(.a(gate135inter0), .b(s_48), .O(gate135inter1));
  and2  gate885(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate886(.a(s_48), .O(gate135inter3));
  inv1  gate887(.a(s_49), .O(gate135inter4));
  nand2 gate888(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate889(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate890(.a(G422), .O(gate135inter7));
  inv1  gate891(.a(G423), .O(gate135inter8));
  nand2 gate892(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate893(.a(s_49), .b(gate135inter3), .O(gate135inter10));
  nor2  gate894(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate895(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate896(.a(gate135inter12), .b(gate135inter1), .O(G516));
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate1611(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate1612(.a(gate144inter0), .b(s_152), .O(gate144inter1));
  and2  gate1613(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate1614(.a(s_152), .O(gate144inter3));
  inv1  gate1615(.a(s_153), .O(gate144inter4));
  nand2 gate1616(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate1617(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate1618(.a(G468), .O(gate144inter7));
  inv1  gate1619(.a(G471), .O(gate144inter8));
  nand2 gate1620(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate1621(.a(s_153), .b(gate144inter3), .O(gate144inter10));
  nor2  gate1622(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate1623(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate1624(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate1625(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate1626(.a(gate147inter0), .b(s_154), .O(gate147inter1));
  and2  gate1627(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate1628(.a(s_154), .O(gate147inter3));
  inv1  gate1629(.a(s_155), .O(gate147inter4));
  nand2 gate1630(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate1631(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate1632(.a(G486), .O(gate147inter7));
  inv1  gate1633(.a(G489), .O(gate147inter8));
  nand2 gate1634(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate1635(.a(s_155), .b(gate147inter3), .O(gate147inter10));
  nor2  gate1636(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate1637(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate1638(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate1807(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate1808(.a(gate151inter0), .b(s_180), .O(gate151inter1));
  and2  gate1809(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate1810(.a(s_180), .O(gate151inter3));
  inv1  gate1811(.a(s_181), .O(gate151inter4));
  nand2 gate1812(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate1813(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate1814(.a(G510), .O(gate151inter7));
  inv1  gate1815(.a(G513), .O(gate151inter8));
  nand2 gate1816(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate1817(.a(s_181), .b(gate151inter3), .O(gate151inter10));
  nor2  gate1818(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate1819(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate1820(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate603(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate604(.a(gate157inter0), .b(s_8), .O(gate157inter1));
  and2  gate605(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate606(.a(s_8), .O(gate157inter3));
  inv1  gate607(.a(s_9), .O(gate157inter4));
  nand2 gate608(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate609(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate610(.a(G438), .O(gate157inter7));
  inv1  gate611(.a(G528), .O(gate157inter8));
  nand2 gate612(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate613(.a(s_9), .b(gate157inter3), .O(gate157inter10));
  nor2  gate614(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate615(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate616(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate1009(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate1010(.a(gate161inter0), .b(s_66), .O(gate161inter1));
  and2  gate1011(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate1012(.a(s_66), .O(gate161inter3));
  inv1  gate1013(.a(s_67), .O(gate161inter4));
  nand2 gate1014(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate1015(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate1016(.a(G450), .O(gate161inter7));
  inv1  gate1017(.a(G534), .O(gate161inter8));
  nand2 gate1018(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate1019(.a(s_67), .b(gate161inter3), .O(gate161inter10));
  nor2  gate1020(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate1021(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate1022(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );

  xor2  gate1373(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate1374(.a(gate163inter0), .b(s_118), .O(gate163inter1));
  and2  gate1375(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate1376(.a(s_118), .O(gate163inter3));
  inv1  gate1377(.a(s_119), .O(gate163inter4));
  nand2 gate1378(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate1379(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate1380(.a(G456), .O(gate163inter7));
  inv1  gate1381(.a(G537), .O(gate163inter8));
  nand2 gate1382(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate1383(.a(s_119), .b(gate163inter3), .O(gate163inter10));
  nor2  gate1384(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate1385(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate1386(.a(gate163inter12), .b(gate163inter1), .O(G580));
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );

  xor2  gate1415(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate1416(.a(gate168inter0), .b(s_124), .O(gate168inter1));
  and2  gate1417(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate1418(.a(s_124), .O(gate168inter3));
  inv1  gate1419(.a(s_125), .O(gate168inter4));
  nand2 gate1420(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate1421(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate1422(.a(G471), .O(gate168inter7));
  inv1  gate1423(.a(G543), .O(gate168inter8));
  nand2 gate1424(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate1425(.a(s_125), .b(gate168inter3), .O(gate168inter10));
  nor2  gate1426(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate1427(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate1428(.a(gate168inter12), .b(gate168inter1), .O(G585));
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );

  xor2  gate1289(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate1290(.a(gate171inter0), .b(s_106), .O(gate171inter1));
  and2  gate1291(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate1292(.a(s_106), .O(gate171inter3));
  inv1  gate1293(.a(s_107), .O(gate171inter4));
  nand2 gate1294(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate1295(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate1296(.a(G480), .O(gate171inter7));
  inv1  gate1297(.a(G549), .O(gate171inter8));
  nand2 gate1298(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate1299(.a(s_107), .b(gate171inter3), .O(gate171inter10));
  nor2  gate1300(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate1301(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate1302(.a(gate171inter12), .b(gate171inter1), .O(G588));
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );

  xor2  gate659(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate660(.a(gate176inter0), .b(s_16), .O(gate176inter1));
  and2  gate661(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate662(.a(s_16), .O(gate176inter3));
  inv1  gate663(.a(s_17), .O(gate176inter4));
  nand2 gate664(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate665(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate666(.a(G495), .O(gate176inter7));
  inv1  gate667(.a(G555), .O(gate176inter8));
  nand2 gate668(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate669(.a(s_17), .b(gate176inter3), .O(gate176inter10));
  nor2  gate670(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate671(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate672(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );

  xor2  gate701(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate702(.a(gate179inter0), .b(s_22), .O(gate179inter1));
  and2  gate703(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate704(.a(s_22), .O(gate179inter3));
  inv1  gate705(.a(s_23), .O(gate179inter4));
  nand2 gate706(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate707(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate708(.a(G504), .O(gate179inter7));
  inv1  gate709(.a(G561), .O(gate179inter8));
  nand2 gate710(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate711(.a(s_23), .b(gate179inter3), .O(gate179inter10));
  nor2  gate712(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate713(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate714(.a(gate179inter12), .b(gate179inter1), .O(G596));
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate1639(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate1640(.a(gate181inter0), .b(s_156), .O(gate181inter1));
  and2  gate1641(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate1642(.a(s_156), .O(gate181inter3));
  inv1  gate1643(.a(s_157), .O(gate181inter4));
  nand2 gate1644(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate1645(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate1646(.a(G510), .O(gate181inter7));
  inv1  gate1647(.a(G564), .O(gate181inter8));
  nand2 gate1648(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate1649(.a(s_157), .b(gate181inter3), .O(gate181inter10));
  nor2  gate1650(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate1651(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate1652(.a(gate181inter12), .b(gate181inter1), .O(G598));

  xor2  gate1177(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate1178(.a(gate182inter0), .b(s_90), .O(gate182inter1));
  and2  gate1179(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate1180(.a(s_90), .O(gate182inter3));
  inv1  gate1181(.a(s_91), .O(gate182inter4));
  nand2 gate1182(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate1183(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate1184(.a(G513), .O(gate182inter7));
  inv1  gate1185(.a(G564), .O(gate182inter8));
  nand2 gate1186(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate1187(.a(s_91), .b(gate182inter3), .O(gate182inter10));
  nor2  gate1188(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate1189(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate1190(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate1569(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate1570(.a(gate184inter0), .b(s_146), .O(gate184inter1));
  and2  gate1571(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate1572(.a(s_146), .O(gate184inter3));
  inv1  gate1573(.a(s_147), .O(gate184inter4));
  nand2 gate1574(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate1575(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate1576(.a(G519), .O(gate184inter7));
  inv1  gate1577(.a(G567), .O(gate184inter8));
  nand2 gate1578(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate1579(.a(s_147), .b(gate184inter3), .O(gate184inter10));
  nor2  gate1580(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate1581(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate1582(.a(gate184inter12), .b(gate184inter1), .O(G601));

  xor2  gate1247(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate1248(.a(gate185inter0), .b(s_100), .O(gate185inter1));
  and2  gate1249(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate1250(.a(s_100), .O(gate185inter3));
  inv1  gate1251(.a(s_101), .O(gate185inter4));
  nand2 gate1252(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate1253(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate1254(.a(G570), .O(gate185inter7));
  inv1  gate1255(.a(G571), .O(gate185inter8));
  nand2 gate1256(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate1257(.a(s_101), .b(gate185inter3), .O(gate185inter10));
  nor2  gate1258(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate1259(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate1260(.a(gate185inter12), .b(gate185inter1), .O(G602));

  xor2  gate1261(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1262(.a(gate186inter0), .b(s_102), .O(gate186inter1));
  and2  gate1263(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1264(.a(s_102), .O(gate186inter3));
  inv1  gate1265(.a(s_103), .O(gate186inter4));
  nand2 gate1266(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1267(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1268(.a(G572), .O(gate186inter7));
  inv1  gate1269(.a(G573), .O(gate186inter8));
  nand2 gate1270(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1271(.a(s_103), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1272(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1273(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1274(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate1751(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate1752(.a(gate188inter0), .b(s_172), .O(gate188inter1));
  and2  gate1753(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate1754(.a(s_172), .O(gate188inter3));
  inv1  gate1755(.a(s_173), .O(gate188inter4));
  nand2 gate1756(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate1757(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate1758(.a(G576), .O(gate188inter7));
  inv1  gate1759(.a(G577), .O(gate188inter8));
  nand2 gate1760(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate1761(.a(s_173), .b(gate188inter3), .O(gate188inter10));
  nor2  gate1762(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate1763(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate1764(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate1303(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate1304(.a(gate193inter0), .b(s_108), .O(gate193inter1));
  and2  gate1305(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate1306(.a(s_108), .O(gate193inter3));
  inv1  gate1307(.a(s_109), .O(gate193inter4));
  nand2 gate1308(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate1309(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate1310(.a(G586), .O(gate193inter7));
  inv1  gate1311(.a(G587), .O(gate193inter8));
  nand2 gate1312(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate1313(.a(s_109), .b(gate193inter3), .O(gate193inter10));
  nor2  gate1314(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate1315(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate1316(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate547(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate548(.a(gate195inter0), .b(s_0), .O(gate195inter1));
  and2  gate549(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate550(.a(s_0), .O(gate195inter3));
  inv1  gate551(.a(s_1), .O(gate195inter4));
  nand2 gate552(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate553(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate554(.a(G590), .O(gate195inter7));
  inv1  gate555(.a(G591), .O(gate195inter8));
  nand2 gate556(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate557(.a(s_1), .b(gate195inter3), .O(gate195inter10));
  nor2  gate558(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate559(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate560(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );

  xor2  gate1541(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate1542(.a(gate199inter0), .b(s_142), .O(gate199inter1));
  and2  gate1543(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate1544(.a(s_142), .O(gate199inter3));
  inv1  gate1545(.a(s_143), .O(gate199inter4));
  nand2 gate1546(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate1547(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate1548(.a(G598), .O(gate199inter7));
  inv1  gate1549(.a(G599), .O(gate199inter8));
  nand2 gate1550(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate1551(.a(s_143), .b(gate199inter3), .O(gate199inter10));
  nor2  gate1552(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate1553(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate1554(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );

  xor2  gate1037(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate1038(.a(gate202inter0), .b(s_70), .O(gate202inter1));
  and2  gate1039(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate1040(.a(s_70), .O(gate202inter3));
  inv1  gate1041(.a(s_71), .O(gate202inter4));
  nand2 gate1042(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate1043(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate1044(.a(G612), .O(gate202inter7));
  inv1  gate1045(.a(G617), .O(gate202inter8));
  nand2 gate1046(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate1047(.a(s_71), .b(gate202inter3), .O(gate202inter10));
  nor2  gate1048(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate1049(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate1050(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );

  xor2  gate631(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate632(.a(gate204inter0), .b(s_12), .O(gate204inter1));
  and2  gate633(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate634(.a(s_12), .O(gate204inter3));
  inv1  gate635(.a(s_13), .O(gate204inter4));
  nand2 gate636(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate637(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate638(.a(G607), .O(gate204inter7));
  inv1  gate639(.a(G617), .O(gate204inter8));
  nand2 gate640(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate641(.a(s_13), .b(gate204inter3), .O(gate204inter10));
  nor2  gate642(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate643(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate644(.a(gate204inter12), .b(gate204inter1), .O(G675));

  xor2  gate1695(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate1696(.a(gate205inter0), .b(s_164), .O(gate205inter1));
  and2  gate1697(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate1698(.a(s_164), .O(gate205inter3));
  inv1  gate1699(.a(s_165), .O(gate205inter4));
  nand2 gate1700(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate1701(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate1702(.a(G622), .O(gate205inter7));
  inv1  gate1703(.a(G627), .O(gate205inter8));
  nand2 gate1704(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate1705(.a(s_165), .b(gate205inter3), .O(gate205inter10));
  nor2  gate1706(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate1707(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate1708(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );

  xor2  gate1359(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate1360(.a(gate207inter0), .b(s_116), .O(gate207inter1));
  and2  gate1361(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate1362(.a(s_116), .O(gate207inter3));
  inv1  gate1363(.a(s_117), .O(gate207inter4));
  nand2 gate1364(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate1365(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate1366(.a(G622), .O(gate207inter7));
  inv1  gate1367(.a(G632), .O(gate207inter8));
  nand2 gate1368(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate1369(.a(s_117), .b(gate207inter3), .O(gate207inter10));
  nor2  gate1370(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate1371(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate1372(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate1135(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate1136(.a(gate213inter0), .b(s_84), .O(gate213inter1));
  and2  gate1137(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate1138(.a(s_84), .O(gate213inter3));
  inv1  gate1139(.a(s_85), .O(gate213inter4));
  nand2 gate1140(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate1141(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate1142(.a(G602), .O(gate213inter7));
  inv1  gate1143(.a(G672), .O(gate213inter8));
  nand2 gate1144(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate1145(.a(s_85), .b(gate213inter3), .O(gate213inter10));
  nor2  gate1146(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate1147(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate1148(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate771(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate772(.a(gate215inter0), .b(s_32), .O(gate215inter1));
  and2  gate773(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate774(.a(s_32), .O(gate215inter3));
  inv1  gate775(.a(s_33), .O(gate215inter4));
  nand2 gate776(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate777(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate778(.a(G607), .O(gate215inter7));
  inv1  gate779(.a(G675), .O(gate215inter8));
  nand2 gate780(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate781(.a(s_33), .b(gate215inter3), .O(gate215inter10));
  nor2  gate782(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate783(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate784(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate1555(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate1556(.a(gate219inter0), .b(s_144), .O(gate219inter1));
  and2  gate1557(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate1558(.a(s_144), .O(gate219inter3));
  inv1  gate1559(.a(s_145), .O(gate219inter4));
  nand2 gate1560(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate1561(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate1562(.a(G632), .O(gate219inter7));
  inv1  gate1563(.a(G681), .O(gate219inter8));
  nand2 gate1564(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate1565(.a(s_145), .b(gate219inter3), .O(gate219inter10));
  nor2  gate1566(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate1567(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate1568(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );

  xor2  gate1065(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate1066(.a(gate225inter0), .b(s_74), .O(gate225inter1));
  and2  gate1067(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate1068(.a(s_74), .O(gate225inter3));
  inv1  gate1069(.a(s_75), .O(gate225inter4));
  nand2 gate1070(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate1071(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate1072(.a(G690), .O(gate225inter7));
  inv1  gate1073(.a(G691), .O(gate225inter8));
  nand2 gate1074(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate1075(.a(s_75), .b(gate225inter3), .O(gate225inter10));
  nor2  gate1076(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate1077(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate1078(.a(gate225inter12), .b(gate225inter1), .O(G706));

  xor2  gate1443(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate1444(.a(gate226inter0), .b(s_128), .O(gate226inter1));
  and2  gate1445(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate1446(.a(s_128), .O(gate226inter3));
  inv1  gate1447(.a(s_129), .O(gate226inter4));
  nand2 gate1448(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate1449(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate1450(.a(G692), .O(gate226inter7));
  inv1  gate1451(.a(G693), .O(gate226inter8));
  nand2 gate1452(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate1453(.a(s_129), .b(gate226inter3), .O(gate226inter10));
  nor2  gate1454(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate1455(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate1456(.a(gate226inter12), .b(gate226inter1), .O(G709));

  xor2  gate1849(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate1850(.a(gate227inter0), .b(s_186), .O(gate227inter1));
  and2  gate1851(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate1852(.a(s_186), .O(gate227inter3));
  inv1  gate1853(.a(s_187), .O(gate227inter4));
  nand2 gate1854(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate1855(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate1856(.a(G694), .O(gate227inter7));
  inv1  gate1857(.a(G695), .O(gate227inter8));
  nand2 gate1858(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate1859(.a(s_187), .b(gate227inter3), .O(gate227inter10));
  nor2  gate1860(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate1861(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate1862(.a(gate227inter12), .b(gate227inter1), .O(G712));
nand2 gate228( .a(G696), .b(G697), .O(G715) );

  xor2  gate1779(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate1780(.a(gate229inter0), .b(s_176), .O(gate229inter1));
  and2  gate1781(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate1782(.a(s_176), .O(gate229inter3));
  inv1  gate1783(.a(s_177), .O(gate229inter4));
  nand2 gate1784(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate1785(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate1786(.a(G698), .O(gate229inter7));
  inv1  gate1787(.a(G699), .O(gate229inter8));
  nand2 gate1788(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate1789(.a(s_177), .b(gate229inter3), .O(gate229inter10));
  nor2  gate1790(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate1791(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate1792(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );

  xor2  gate1275(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate1276(.a(gate232inter0), .b(s_104), .O(gate232inter1));
  and2  gate1277(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate1278(.a(s_104), .O(gate232inter3));
  inv1  gate1279(.a(s_105), .O(gate232inter4));
  nand2 gate1280(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate1281(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate1282(.a(G704), .O(gate232inter7));
  inv1  gate1283(.a(G705), .O(gate232inter8));
  nand2 gate1284(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate1285(.a(s_105), .b(gate232inter3), .O(gate232inter10));
  nor2  gate1286(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate1287(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate1288(.a(gate232inter12), .b(gate232inter1), .O(G727));
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );

  xor2  gate939(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate940(.a(gate238inter0), .b(s_56), .O(gate238inter1));
  and2  gate941(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate942(.a(s_56), .O(gate238inter3));
  inv1  gate943(.a(s_57), .O(gate238inter4));
  nand2 gate944(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate945(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate946(.a(G257), .O(gate238inter7));
  inv1  gate947(.a(G709), .O(gate238inter8));
  nand2 gate948(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate949(.a(s_57), .b(gate238inter3), .O(gate238inter10));
  nor2  gate950(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate951(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate952(.a(gate238inter12), .b(gate238inter1), .O(G745));

  xor2  gate1597(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate1598(.a(gate239inter0), .b(s_150), .O(gate239inter1));
  and2  gate1599(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate1600(.a(s_150), .O(gate239inter3));
  inv1  gate1601(.a(s_151), .O(gate239inter4));
  nand2 gate1602(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate1603(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate1604(.a(G260), .O(gate239inter7));
  inv1  gate1605(.a(G712), .O(gate239inter8));
  nand2 gate1606(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate1607(.a(s_151), .b(gate239inter3), .O(gate239inter10));
  nor2  gate1608(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate1609(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate1610(.a(gate239inter12), .b(gate239inter1), .O(G748));

  xor2  gate1331(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate1332(.a(gate240inter0), .b(s_112), .O(gate240inter1));
  and2  gate1333(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate1334(.a(s_112), .O(gate240inter3));
  inv1  gate1335(.a(s_113), .O(gate240inter4));
  nand2 gate1336(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate1337(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate1338(.a(G263), .O(gate240inter7));
  inv1  gate1339(.a(G715), .O(gate240inter8));
  nand2 gate1340(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate1341(.a(s_113), .b(gate240inter3), .O(gate240inter10));
  nor2  gate1342(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate1343(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate1344(.a(gate240inter12), .b(gate240inter1), .O(G751));

  xor2  gate687(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate688(.a(gate241inter0), .b(s_20), .O(gate241inter1));
  and2  gate689(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate690(.a(s_20), .O(gate241inter3));
  inv1  gate691(.a(s_21), .O(gate241inter4));
  nand2 gate692(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate693(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate694(.a(G242), .O(gate241inter7));
  inv1  gate695(.a(G730), .O(gate241inter8));
  nand2 gate696(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate697(.a(s_21), .b(gate241inter3), .O(gate241inter10));
  nor2  gate698(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate699(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate700(.a(gate241inter12), .b(gate241inter1), .O(G754));

  xor2  gate1989(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate1990(.a(gate242inter0), .b(s_206), .O(gate242inter1));
  and2  gate1991(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate1992(.a(s_206), .O(gate242inter3));
  inv1  gate1993(.a(s_207), .O(gate242inter4));
  nand2 gate1994(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate1995(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate1996(.a(G718), .O(gate242inter7));
  inv1  gate1997(.a(G730), .O(gate242inter8));
  nand2 gate1998(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate1999(.a(s_207), .b(gate242inter3), .O(gate242inter10));
  nor2  gate2000(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate2001(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate2002(.a(gate242inter12), .b(gate242inter1), .O(G755));
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate1821(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate1822(.a(gate245inter0), .b(s_182), .O(gate245inter1));
  and2  gate1823(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate1824(.a(s_182), .O(gate245inter3));
  inv1  gate1825(.a(s_183), .O(gate245inter4));
  nand2 gate1826(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate1827(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate1828(.a(G248), .O(gate245inter7));
  inv1  gate1829(.a(G736), .O(gate245inter8));
  nand2 gate1830(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate1831(.a(s_183), .b(gate245inter3), .O(gate245inter10));
  nor2  gate1832(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate1833(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate1834(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );

  xor2  gate673(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate674(.a(gate247inter0), .b(s_18), .O(gate247inter1));
  and2  gate675(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate676(.a(s_18), .O(gate247inter3));
  inv1  gate677(.a(s_19), .O(gate247inter4));
  nand2 gate678(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate679(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate680(.a(G251), .O(gate247inter7));
  inv1  gate681(.a(G739), .O(gate247inter8));
  nand2 gate682(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate683(.a(s_19), .b(gate247inter3), .O(gate247inter10));
  nor2  gate684(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate685(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate686(.a(gate247inter12), .b(gate247inter1), .O(G760));
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate1793(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate1794(.a(gate249inter0), .b(s_178), .O(gate249inter1));
  and2  gate1795(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate1796(.a(s_178), .O(gate249inter3));
  inv1  gate1797(.a(s_179), .O(gate249inter4));
  nand2 gate1798(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate1799(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate1800(.a(G254), .O(gate249inter7));
  inv1  gate1801(.a(G742), .O(gate249inter8));
  nand2 gate1802(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate1803(.a(s_179), .b(gate249inter3), .O(gate249inter10));
  nor2  gate1804(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate1805(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate1806(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate1919(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate1920(.a(gate263inter0), .b(s_196), .O(gate263inter1));
  and2  gate1921(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate1922(.a(s_196), .O(gate263inter3));
  inv1  gate1923(.a(s_197), .O(gate263inter4));
  nand2 gate1924(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate1925(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate1926(.a(G766), .O(gate263inter7));
  inv1  gate1927(.a(G767), .O(gate263inter8));
  nand2 gate1928(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate1929(.a(s_197), .b(gate263inter3), .O(gate263inter10));
  nor2  gate1930(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate1931(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate1932(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate1527(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate1528(.a(gate268inter0), .b(s_140), .O(gate268inter1));
  and2  gate1529(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate1530(.a(s_140), .O(gate268inter3));
  inv1  gate1531(.a(s_141), .O(gate268inter4));
  nand2 gate1532(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1533(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1534(.a(G651), .O(gate268inter7));
  inv1  gate1535(.a(G779), .O(gate268inter8));
  nand2 gate1536(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1537(.a(s_141), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1538(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1539(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1540(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate1149(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate1150(.a(gate272inter0), .b(s_86), .O(gate272inter1));
  and2  gate1151(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate1152(.a(s_86), .O(gate272inter3));
  inv1  gate1153(.a(s_87), .O(gate272inter4));
  nand2 gate1154(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate1155(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate1156(.a(G663), .O(gate272inter7));
  inv1  gate1157(.a(G791), .O(gate272inter8));
  nand2 gate1158(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate1159(.a(s_87), .b(gate272inter3), .O(gate272inter10));
  nor2  gate1160(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate1161(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate1162(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate645(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate646(.a(gate276inter0), .b(s_14), .O(gate276inter1));
  and2  gate647(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate648(.a(s_14), .O(gate276inter3));
  inv1  gate649(.a(s_15), .O(gate276inter4));
  nand2 gate650(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate651(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate652(.a(G773), .O(gate276inter7));
  inv1  gate653(.a(G797), .O(gate276inter8));
  nand2 gate654(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate655(.a(s_15), .b(gate276inter3), .O(gate276inter10));
  nor2  gate656(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate657(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate658(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate1429(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate1430(.a(gate278inter0), .b(s_126), .O(gate278inter1));
  and2  gate1431(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate1432(.a(s_126), .O(gate278inter3));
  inv1  gate1433(.a(s_127), .O(gate278inter4));
  nand2 gate1434(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate1435(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate1436(.a(G776), .O(gate278inter7));
  inv1  gate1437(.a(G800), .O(gate278inter8));
  nand2 gate1438(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate1439(.a(s_127), .b(gate278inter3), .O(gate278inter10));
  nor2  gate1440(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate1441(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate1442(.a(gate278inter12), .b(gate278inter1), .O(G823));

  xor2  gate575(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate576(.a(gate279inter0), .b(s_4), .O(gate279inter1));
  and2  gate577(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate578(.a(s_4), .O(gate279inter3));
  inv1  gate579(.a(s_5), .O(gate279inter4));
  nand2 gate580(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate581(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate582(.a(G651), .O(gate279inter7));
  inv1  gate583(.a(G803), .O(gate279inter8));
  nand2 gate584(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate585(.a(s_5), .b(gate279inter3), .O(gate279inter10));
  nor2  gate586(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate587(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate588(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate1401(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate1402(.a(gate283inter0), .b(s_122), .O(gate283inter1));
  and2  gate1403(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate1404(.a(s_122), .O(gate283inter3));
  inv1  gate1405(.a(s_123), .O(gate283inter4));
  nand2 gate1406(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate1407(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate1408(.a(G657), .O(gate283inter7));
  inv1  gate1409(.a(G809), .O(gate283inter8));
  nand2 gate1410(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate1411(.a(s_123), .b(gate283inter3), .O(gate283inter10));
  nor2  gate1412(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate1413(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate1414(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate729(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate730(.a(gate289inter0), .b(s_26), .O(gate289inter1));
  and2  gate731(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate732(.a(s_26), .O(gate289inter3));
  inv1  gate733(.a(s_27), .O(gate289inter4));
  nand2 gate734(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate735(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate736(.a(G818), .O(gate289inter7));
  inv1  gate737(.a(G819), .O(gate289inter8));
  nand2 gate738(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate739(.a(s_27), .b(gate289inter3), .O(gate289inter10));
  nor2  gate740(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate741(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate742(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate1457(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate1458(.a(gate293inter0), .b(s_130), .O(gate293inter1));
  and2  gate1459(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate1460(.a(s_130), .O(gate293inter3));
  inv1  gate1461(.a(s_131), .O(gate293inter4));
  nand2 gate1462(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate1463(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate1464(.a(G828), .O(gate293inter7));
  inv1  gate1465(.a(G829), .O(gate293inter8));
  nand2 gate1466(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate1467(.a(s_131), .b(gate293inter3), .O(gate293inter10));
  nor2  gate1468(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate1469(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate1470(.a(gate293inter12), .b(gate293inter1), .O(G886));

  xor2  gate1765(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate1766(.a(gate294inter0), .b(s_174), .O(gate294inter1));
  and2  gate1767(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate1768(.a(s_174), .O(gate294inter3));
  inv1  gate1769(.a(s_175), .O(gate294inter4));
  nand2 gate1770(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate1771(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate1772(.a(G832), .O(gate294inter7));
  inv1  gate1773(.a(G833), .O(gate294inter8));
  nand2 gate1774(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate1775(.a(s_175), .b(gate294inter3), .O(gate294inter10));
  nor2  gate1776(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate1777(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate1778(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate1667(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate1668(.a(gate391inter0), .b(s_160), .O(gate391inter1));
  and2  gate1669(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate1670(.a(s_160), .O(gate391inter3));
  inv1  gate1671(.a(s_161), .O(gate391inter4));
  nand2 gate1672(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate1673(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate1674(.a(G5), .O(gate391inter7));
  inv1  gate1675(.a(G1048), .O(gate391inter8));
  nand2 gate1676(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate1677(.a(s_161), .b(gate391inter3), .O(gate391inter10));
  nor2  gate1678(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate1679(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate1680(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate2017(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate2018(.a(gate395inter0), .b(s_210), .O(gate395inter1));
  and2  gate2019(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate2020(.a(s_210), .O(gate395inter3));
  inv1  gate2021(.a(s_211), .O(gate395inter4));
  nand2 gate2022(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate2023(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate2024(.a(G9), .O(gate395inter7));
  inv1  gate2025(.a(G1060), .O(gate395inter8));
  nand2 gate2026(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate2027(.a(s_211), .b(gate395inter3), .O(gate395inter10));
  nor2  gate2028(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate2029(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate2030(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );

  xor2  gate1471(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate1472(.a(gate404inter0), .b(s_132), .O(gate404inter1));
  and2  gate1473(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate1474(.a(s_132), .O(gate404inter3));
  inv1  gate1475(.a(s_133), .O(gate404inter4));
  nand2 gate1476(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate1477(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate1478(.a(G18), .O(gate404inter7));
  inv1  gate1479(.a(G1087), .O(gate404inter8));
  nand2 gate1480(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate1481(.a(s_133), .b(gate404inter3), .O(gate404inter10));
  nor2  gate1482(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate1483(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate1484(.a(gate404inter12), .b(gate404inter1), .O(G1183));
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate1681(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate1682(.a(gate411inter0), .b(s_162), .O(gate411inter1));
  and2  gate1683(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate1684(.a(s_162), .O(gate411inter3));
  inv1  gate1685(.a(s_163), .O(gate411inter4));
  nand2 gate1686(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate1687(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate1688(.a(G25), .O(gate411inter7));
  inv1  gate1689(.a(G1108), .O(gate411inter8));
  nand2 gate1690(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate1691(.a(s_163), .b(gate411inter3), .O(gate411inter10));
  nor2  gate1692(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate1693(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate1694(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );

  xor2  gate1317(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate1318(.a(gate416inter0), .b(s_110), .O(gate416inter1));
  and2  gate1319(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate1320(.a(s_110), .O(gate416inter3));
  inv1  gate1321(.a(s_111), .O(gate416inter4));
  nand2 gate1322(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate1323(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate1324(.a(G30), .O(gate416inter7));
  inv1  gate1325(.a(G1123), .O(gate416inter8));
  nand2 gate1326(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate1327(.a(s_111), .b(gate416inter3), .O(gate416inter10));
  nor2  gate1328(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate1329(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate1330(.a(gate416inter12), .b(gate416inter1), .O(G1219));
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );

  xor2  gate1051(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate1052(.a(gate418inter0), .b(s_72), .O(gate418inter1));
  and2  gate1053(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate1054(.a(s_72), .O(gate418inter3));
  inv1  gate1055(.a(s_73), .O(gate418inter4));
  nand2 gate1056(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate1057(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate1058(.a(G32), .O(gate418inter7));
  inv1  gate1059(.a(G1129), .O(gate418inter8));
  nand2 gate1060(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate1061(.a(s_73), .b(gate418inter3), .O(gate418inter10));
  nor2  gate1062(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate1063(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate1064(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate1947(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate1948(.a(gate421inter0), .b(s_200), .O(gate421inter1));
  and2  gate1949(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate1950(.a(s_200), .O(gate421inter3));
  inv1  gate1951(.a(s_201), .O(gate421inter4));
  nand2 gate1952(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate1953(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate1954(.a(G2), .O(gate421inter7));
  inv1  gate1955(.a(G1135), .O(gate421inter8));
  nand2 gate1956(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate1957(.a(s_201), .b(gate421inter3), .O(gate421inter10));
  nor2  gate1958(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate1959(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate1960(.a(gate421inter12), .b(gate421inter1), .O(G1230));
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );

  xor2  gate1219(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate1220(.a(gate427inter0), .b(s_96), .O(gate427inter1));
  and2  gate1221(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate1222(.a(s_96), .O(gate427inter3));
  inv1  gate1223(.a(s_97), .O(gate427inter4));
  nand2 gate1224(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate1225(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate1226(.a(G5), .O(gate427inter7));
  inv1  gate1227(.a(G1144), .O(gate427inter8));
  nand2 gate1228(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate1229(.a(s_97), .b(gate427inter3), .O(gate427inter10));
  nor2  gate1230(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate1231(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate1232(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate995(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate996(.a(gate430inter0), .b(s_64), .O(gate430inter1));
  and2  gate997(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate998(.a(s_64), .O(gate430inter3));
  inv1  gate999(.a(s_65), .O(gate430inter4));
  nand2 gate1000(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate1001(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate1002(.a(G1051), .O(gate430inter7));
  inv1  gate1003(.a(G1147), .O(gate430inter8));
  nand2 gate1004(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate1005(.a(s_65), .b(gate430inter3), .O(gate430inter10));
  nor2  gate1006(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate1007(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate1008(.a(gate430inter12), .b(gate430inter1), .O(G1239));

  xor2  gate2003(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate2004(.a(gate431inter0), .b(s_208), .O(gate431inter1));
  and2  gate2005(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate2006(.a(s_208), .O(gate431inter3));
  inv1  gate2007(.a(s_209), .O(gate431inter4));
  nand2 gate2008(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate2009(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate2010(.a(G7), .O(gate431inter7));
  inv1  gate2011(.a(G1150), .O(gate431inter8));
  nand2 gate2012(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate2013(.a(s_209), .b(gate431inter3), .O(gate431inter10));
  nor2  gate2014(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate2015(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate2016(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate1737(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate1738(.a(gate438inter0), .b(s_170), .O(gate438inter1));
  and2  gate1739(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate1740(.a(s_170), .O(gate438inter3));
  inv1  gate1741(.a(s_171), .O(gate438inter4));
  nand2 gate1742(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate1743(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate1744(.a(G1063), .O(gate438inter7));
  inv1  gate1745(.a(G1159), .O(gate438inter8));
  nand2 gate1746(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate1747(.a(s_171), .b(gate438inter3), .O(gate438inter10));
  nor2  gate1748(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate1749(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate1750(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate1485(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate1486(.a(gate444inter0), .b(s_134), .O(gate444inter1));
  and2  gate1487(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate1488(.a(s_134), .O(gate444inter3));
  inv1  gate1489(.a(s_135), .O(gate444inter4));
  nand2 gate1490(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate1491(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate1492(.a(G1072), .O(gate444inter7));
  inv1  gate1493(.a(G1168), .O(gate444inter8));
  nand2 gate1494(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate1495(.a(s_135), .b(gate444inter3), .O(gate444inter10));
  nor2  gate1496(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate1497(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate1498(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate1513(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate1514(.a(gate448inter0), .b(s_138), .O(gate448inter1));
  and2  gate1515(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate1516(.a(s_138), .O(gate448inter3));
  inv1  gate1517(.a(s_139), .O(gate448inter4));
  nand2 gate1518(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate1519(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate1520(.a(G1078), .O(gate448inter7));
  inv1  gate1521(.a(G1174), .O(gate448inter8));
  nand2 gate1522(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate1523(.a(s_139), .b(gate448inter3), .O(gate448inter10));
  nor2  gate1524(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate1525(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate1526(.a(gate448inter12), .b(gate448inter1), .O(G1257));

  xor2  gate1163(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate1164(.a(gate449inter0), .b(s_88), .O(gate449inter1));
  and2  gate1165(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate1166(.a(s_88), .O(gate449inter3));
  inv1  gate1167(.a(s_89), .O(gate449inter4));
  nand2 gate1168(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate1169(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate1170(.a(G16), .O(gate449inter7));
  inv1  gate1171(.a(G1177), .O(gate449inter8));
  nand2 gate1172(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate1173(.a(s_89), .b(gate449inter3), .O(gate449inter10));
  nor2  gate1174(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate1175(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate1176(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate617(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate618(.a(gate461inter0), .b(s_10), .O(gate461inter1));
  and2  gate619(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate620(.a(s_10), .O(gate461inter3));
  inv1  gate621(.a(s_11), .O(gate461inter4));
  nand2 gate622(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate623(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate624(.a(G22), .O(gate461inter7));
  inv1  gate625(.a(G1195), .O(gate461inter8));
  nand2 gate626(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate627(.a(s_11), .b(gate461inter3), .O(gate461inter10));
  nor2  gate628(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate629(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate630(.a(gate461inter12), .b(gate461inter1), .O(G1270));
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate897(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate898(.a(gate464inter0), .b(s_50), .O(gate464inter1));
  and2  gate899(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate900(.a(s_50), .O(gate464inter3));
  inv1  gate901(.a(s_51), .O(gate464inter4));
  nand2 gate902(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate903(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate904(.a(G1102), .O(gate464inter7));
  inv1  gate905(.a(G1198), .O(gate464inter8));
  nand2 gate906(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate907(.a(s_51), .b(gate464inter3), .O(gate464inter10));
  nor2  gate908(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate909(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate910(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate561(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate562(.a(gate467inter0), .b(s_2), .O(gate467inter1));
  and2  gate563(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate564(.a(s_2), .O(gate467inter3));
  inv1  gate565(.a(s_3), .O(gate467inter4));
  nand2 gate566(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate567(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate568(.a(G25), .O(gate467inter7));
  inv1  gate569(.a(G1204), .O(gate467inter8));
  nand2 gate570(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate571(.a(s_3), .b(gate467inter3), .O(gate467inter10));
  nor2  gate572(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate573(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate574(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate827(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate828(.a(gate475inter0), .b(s_40), .O(gate475inter1));
  and2  gate829(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate830(.a(s_40), .O(gate475inter3));
  inv1  gate831(.a(s_41), .O(gate475inter4));
  nand2 gate832(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate833(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate834(.a(G29), .O(gate475inter7));
  inv1  gate835(.a(G1216), .O(gate475inter8));
  nand2 gate836(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate837(.a(s_41), .b(gate475inter3), .O(gate475inter10));
  nor2  gate838(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate839(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate840(.a(gate475inter12), .b(gate475inter1), .O(G1284));

  xor2  gate1961(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate1962(.a(gate476inter0), .b(s_202), .O(gate476inter1));
  and2  gate1963(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate1964(.a(s_202), .O(gate476inter3));
  inv1  gate1965(.a(s_203), .O(gate476inter4));
  nand2 gate1966(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate1967(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate1968(.a(G1120), .O(gate476inter7));
  inv1  gate1969(.a(G1216), .O(gate476inter8));
  nand2 gate1970(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate1971(.a(s_203), .b(gate476inter3), .O(gate476inter10));
  nor2  gate1972(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate1973(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate1974(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );

  xor2  gate743(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate744(.a(gate483inter0), .b(s_28), .O(gate483inter1));
  and2  gate745(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate746(.a(s_28), .O(gate483inter3));
  inv1  gate747(.a(s_29), .O(gate483inter4));
  nand2 gate748(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate749(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate750(.a(G1228), .O(gate483inter7));
  inv1  gate751(.a(G1229), .O(gate483inter8));
  nand2 gate752(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate753(.a(s_29), .b(gate483inter3), .O(gate483inter10));
  nor2  gate754(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate755(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate756(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate967(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate968(.a(gate486inter0), .b(s_60), .O(gate486inter1));
  and2  gate969(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate970(.a(s_60), .O(gate486inter3));
  inv1  gate971(.a(s_61), .O(gate486inter4));
  nand2 gate972(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate973(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate974(.a(G1234), .O(gate486inter7));
  inv1  gate975(.a(G1235), .O(gate486inter8));
  nand2 gate976(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate977(.a(s_61), .b(gate486inter3), .O(gate486inter10));
  nor2  gate978(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate979(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate980(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate953(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate954(.a(gate488inter0), .b(s_58), .O(gate488inter1));
  and2  gate955(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate956(.a(s_58), .O(gate488inter3));
  inv1  gate957(.a(s_59), .O(gate488inter4));
  nand2 gate958(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate959(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate960(.a(G1238), .O(gate488inter7));
  inv1  gate961(.a(G1239), .O(gate488inter8));
  nand2 gate962(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate963(.a(s_59), .b(gate488inter3), .O(gate488inter10));
  nor2  gate964(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate965(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate966(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate1093(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate1094(.a(gate492inter0), .b(s_78), .O(gate492inter1));
  and2  gate1095(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate1096(.a(s_78), .O(gate492inter3));
  inv1  gate1097(.a(s_79), .O(gate492inter4));
  nand2 gate1098(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate1099(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate1100(.a(G1246), .O(gate492inter7));
  inv1  gate1101(.a(G1247), .O(gate492inter8));
  nand2 gate1102(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate1103(.a(s_79), .b(gate492inter3), .O(gate492inter10));
  nor2  gate1104(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate1105(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate1106(.a(gate492inter12), .b(gate492inter1), .O(G1301));
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate1933(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate1934(.a(gate499inter0), .b(s_198), .O(gate499inter1));
  and2  gate1935(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate1936(.a(s_198), .O(gate499inter3));
  inv1  gate1937(.a(s_199), .O(gate499inter4));
  nand2 gate1938(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate1939(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate1940(.a(G1260), .O(gate499inter7));
  inv1  gate1941(.a(G1261), .O(gate499inter8));
  nand2 gate1942(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate1943(.a(s_199), .b(gate499inter3), .O(gate499inter10));
  nor2  gate1944(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate1945(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate1946(.a(gate499inter12), .b(gate499inter1), .O(G1308));

  xor2  gate869(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate870(.a(gate500inter0), .b(s_46), .O(gate500inter1));
  and2  gate871(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate872(.a(s_46), .O(gate500inter3));
  inv1  gate873(.a(s_47), .O(gate500inter4));
  nand2 gate874(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate875(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate876(.a(G1262), .O(gate500inter7));
  inv1  gate877(.a(G1263), .O(gate500inter8));
  nand2 gate878(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate879(.a(s_47), .b(gate500inter3), .O(gate500inter10));
  nor2  gate880(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate881(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate882(.a(gate500inter12), .b(gate500inter1), .O(G1309));
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );

  xor2  gate757(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate758(.a(gate513inter0), .b(s_30), .O(gate513inter1));
  and2  gate759(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate760(.a(s_30), .O(gate513inter3));
  inv1  gate761(.a(s_31), .O(gate513inter4));
  nand2 gate762(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate763(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate764(.a(G1288), .O(gate513inter7));
  inv1  gate765(.a(G1289), .O(gate513inter8));
  nand2 gate766(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate767(.a(s_31), .b(gate513inter3), .O(gate513inter10));
  nor2  gate768(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate769(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate770(.a(gate513inter12), .b(gate513inter1), .O(G1322));

  xor2  gate1191(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate1192(.a(gate514inter0), .b(s_92), .O(gate514inter1));
  and2  gate1193(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate1194(.a(s_92), .O(gate514inter3));
  inv1  gate1195(.a(s_93), .O(gate514inter4));
  nand2 gate1196(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate1197(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate1198(.a(G1290), .O(gate514inter7));
  inv1  gate1199(.a(G1291), .O(gate514inter8));
  nand2 gate1200(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate1201(.a(s_93), .b(gate514inter3), .O(gate514inter10));
  nor2  gate1202(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate1203(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate1204(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule