module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281, s_282, s_283, s_284, s_285, s_286, s_287, s_288, s_289, s_290, s_291, s_292, s_293, s_294, s_295, s_296, s_297, s_298, s_299, s_300, s_301, s_302, s_303, s_304, s_305, s_306, s_307, s_308, s_309, s_310, s_311, s_312, s_313, s_314, s_315, s_316, s_317, s_318, s_319, s_320, s_321, s_322, s_323, s_324, s_325, s_326, s_327, s_328, s_329, s_330, s_331, s_332, s_333, s_334, s_335, s_336, s_337, s_338, s_339, s_340, s_341, s_342, s_343, s_344, s_345, s_346, s_347, s_348, s_349, s_350, s_351, s_352, s_353, s_354, s_355, s_356, s_357, s_358, s_359, s_360, s_361;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate2003(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate2004(.a(gate9inter0), .b(s_208), .O(gate9inter1));
  and2  gate2005(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate2006(.a(s_208), .O(gate9inter3));
  inv1  gate2007(.a(s_209), .O(gate9inter4));
  nand2 gate2008(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate2009(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate2010(.a(G1), .O(gate9inter7));
  inv1  gate2011(.a(G2), .O(gate9inter8));
  nand2 gate2012(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate2013(.a(s_209), .b(gate9inter3), .O(gate9inter10));
  nor2  gate2014(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate2015(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate2016(.a(gate9inter12), .b(gate9inter1), .O(G266));

  xor2  gate2311(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate2312(.a(gate10inter0), .b(s_252), .O(gate10inter1));
  and2  gate2313(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate2314(.a(s_252), .O(gate10inter3));
  inv1  gate2315(.a(s_253), .O(gate10inter4));
  nand2 gate2316(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate2317(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate2318(.a(G3), .O(gate10inter7));
  inv1  gate2319(.a(G4), .O(gate10inter8));
  nand2 gate2320(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate2321(.a(s_253), .b(gate10inter3), .O(gate10inter10));
  nor2  gate2322(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate2323(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate2324(.a(gate10inter12), .b(gate10inter1), .O(G269));

  xor2  gate2017(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate2018(.a(gate11inter0), .b(s_210), .O(gate11inter1));
  and2  gate2019(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate2020(.a(s_210), .O(gate11inter3));
  inv1  gate2021(.a(s_211), .O(gate11inter4));
  nand2 gate2022(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate2023(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate2024(.a(G5), .O(gate11inter7));
  inv1  gate2025(.a(G6), .O(gate11inter8));
  nand2 gate2026(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate2027(.a(s_211), .b(gate11inter3), .O(gate11inter10));
  nor2  gate2028(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate2029(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate2030(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );

  xor2  gate1961(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate1962(.a(gate14inter0), .b(s_202), .O(gate14inter1));
  and2  gate1963(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate1964(.a(s_202), .O(gate14inter3));
  inv1  gate1965(.a(s_203), .O(gate14inter4));
  nand2 gate1966(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate1967(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate1968(.a(G11), .O(gate14inter7));
  inv1  gate1969(.a(G12), .O(gate14inter8));
  nand2 gate1970(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate1971(.a(s_203), .b(gate14inter3), .O(gate14inter10));
  nor2  gate1972(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate1973(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate1974(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate1989(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate1990(.a(gate17inter0), .b(s_206), .O(gate17inter1));
  and2  gate1991(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate1992(.a(s_206), .O(gate17inter3));
  inv1  gate1993(.a(s_207), .O(gate17inter4));
  nand2 gate1994(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate1995(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate1996(.a(G17), .O(gate17inter7));
  inv1  gate1997(.a(G18), .O(gate17inter8));
  nand2 gate1998(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate1999(.a(s_207), .b(gate17inter3), .O(gate17inter10));
  nor2  gate2000(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate2001(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate2002(.a(gate17inter12), .b(gate17inter1), .O(G290));

  xor2  gate883(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate884(.a(gate18inter0), .b(s_48), .O(gate18inter1));
  and2  gate885(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate886(.a(s_48), .O(gate18inter3));
  inv1  gate887(.a(s_49), .O(gate18inter4));
  nand2 gate888(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate889(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate890(.a(G19), .O(gate18inter7));
  inv1  gate891(.a(G20), .O(gate18inter8));
  nand2 gate892(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate893(.a(s_49), .b(gate18inter3), .O(gate18inter10));
  nor2  gate894(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate895(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate896(.a(gate18inter12), .b(gate18inter1), .O(G293));

  xor2  gate785(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate786(.a(gate19inter0), .b(s_34), .O(gate19inter1));
  and2  gate787(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate788(.a(s_34), .O(gate19inter3));
  inv1  gate789(.a(s_35), .O(gate19inter4));
  nand2 gate790(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate791(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate792(.a(G21), .O(gate19inter7));
  inv1  gate793(.a(G22), .O(gate19inter8));
  nand2 gate794(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate795(.a(s_35), .b(gate19inter3), .O(gate19inter10));
  nor2  gate796(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate797(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate798(.a(gate19inter12), .b(gate19inter1), .O(G296));

  xor2  gate2885(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate2886(.a(gate20inter0), .b(s_334), .O(gate20inter1));
  and2  gate2887(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate2888(.a(s_334), .O(gate20inter3));
  inv1  gate2889(.a(s_335), .O(gate20inter4));
  nand2 gate2890(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate2891(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate2892(.a(G23), .O(gate20inter7));
  inv1  gate2893(.a(G24), .O(gate20inter8));
  nand2 gate2894(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate2895(.a(s_335), .b(gate20inter3), .O(gate20inter10));
  nor2  gate2896(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate2897(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate2898(.a(gate20inter12), .b(gate20inter1), .O(G299));

  xor2  gate1457(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate1458(.a(gate21inter0), .b(s_130), .O(gate21inter1));
  and2  gate1459(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate1460(.a(s_130), .O(gate21inter3));
  inv1  gate1461(.a(s_131), .O(gate21inter4));
  nand2 gate1462(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate1463(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate1464(.a(G25), .O(gate21inter7));
  inv1  gate1465(.a(G26), .O(gate21inter8));
  nand2 gate1466(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate1467(.a(s_131), .b(gate21inter3), .O(gate21inter10));
  nor2  gate1468(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate1469(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate1470(.a(gate21inter12), .b(gate21inter1), .O(G302));
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate1345(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate1346(.a(gate23inter0), .b(s_114), .O(gate23inter1));
  and2  gate1347(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate1348(.a(s_114), .O(gate23inter3));
  inv1  gate1349(.a(s_115), .O(gate23inter4));
  nand2 gate1350(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate1351(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate1352(.a(G29), .O(gate23inter7));
  inv1  gate1353(.a(G30), .O(gate23inter8));
  nand2 gate1354(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate1355(.a(s_115), .b(gate23inter3), .O(gate23inter10));
  nor2  gate1356(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate1357(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate1358(.a(gate23inter12), .b(gate23inter1), .O(G308));

  xor2  gate2171(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate2172(.a(gate24inter0), .b(s_232), .O(gate24inter1));
  and2  gate2173(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate2174(.a(s_232), .O(gate24inter3));
  inv1  gate2175(.a(s_233), .O(gate24inter4));
  nand2 gate2176(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate2177(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate2178(.a(G31), .O(gate24inter7));
  inv1  gate2179(.a(G32), .O(gate24inter8));
  nand2 gate2180(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate2181(.a(s_233), .b(gate24inter3), .O(gate24inter10));
  nor2  gate2182(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate2183(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate2184(.a(gate24inter12), .b(gate24inter1), .O(G311));

  xor2  gate2269(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate2270(.a(gate25inter0), .b(s_246), .O(gate25inter1));
  and2  gate2271(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate2272(.a(s_246), .O(gate25inter3));
  inv1  gate2273(.a(s_247), .O(gate25inter4));
  nand2 gate2274(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate2275(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate2276(.a(G1), .O(gate25inter7));
  inv1  gate2277(.a(G5), .O(gate25inter8));
  nand2 gate2278(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate2279(.a(s_247), .b(gate25inter3), .O(gate25inter10));
  nor2  gate2280(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate2281(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate2282(.a(gate25inter12), .b(gate25inter1), .O(G314));

  xor2  gate1415(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate1416(.a(gate26inter0), .b(s_124), .O(gate26inter1));
  and2  gate1417(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate1418(.a(s_124), .O(gate26inter3));
  inv1  gate1419(.a(s_125), .O(gate26inter4));
  nand2 gate1420(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate1421(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate1422(.a(G9), .O(gate26inter7));
  inv1  gate1423(.a(G13), .O(gate26inter8));
  nand2 gate1424(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate1425(.a(s_125), .b(gate26inter3), .O(gate26inter10));
  nor2  gate1426(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate1427(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate1428(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate1443(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate1444(.a(gate28inter0), .b(s_128), .O(gate28inter1));
  and2  gate1445(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate1446(.a(s_128), .O(gate28inter3));
  inv1  gate1447(.a(s_129), .O(gate28inter4));
  nand2 gate1448(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate1449(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate1450(.a(G10), .O(gate28inter7));
  inv1  gate1451(.a(G14), .O(gate28inter8));
  nand2 gate1452(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate1453(.a(s_129), .b(gate28inter3), .O(gate28inter10));
  nor2  gate1454(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate1455(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate1456(.a(gate28inter12), .b(gate28inter1), .O(G323));

  xor2  gate2899(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate2900(.a(gate29inter0), .b(s_336), .O(gate29inter1));
  and2  gate2901(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate2902(.a(s_336), .O(gate29inter3));
  inv1  gate2903(.a(s_337), .O(gate29inter4));
  nand2 gate2904(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate2905(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate2906(.a(G3), .O(gate29inter7));
  inv1  gate2907(.a(G7), .O(gate29inter8));
  nand2 gate2908(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate2909(.a(s_337), .b(gate29inter3), .O(gate29inter10));
  nor2  gate2910(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate2911(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate2912(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );

  xor2  gate2073(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate2074(.a(gate32inter0), .b(s_218), .O(gate32inter1));
  and2  gate2075(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate2076(.a(s_218), .O(gate32inter3));
  inv1  gate2077(.a(s_219), .O(gate32inter4));
  nand2 gate2078(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate2079(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate2080(.a(G12), .O(gate32inter7));
  inv1  gate2081(.a(G16), .O(gate32inter8));
  nand2 gate2082(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate2083(.a(s_219), .b(gate32inter3), .O(gate32inter10));
  nor2  gate2084(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate2085(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate2086(.a(gate32inter12), .b(gate32inter1), .O(G335));

  xor2  gate1667(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate1668(.a(gate33inter0), .b(s_160), .O(gate33inter1));
  and2  gate1669(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate1670(.a(s_160), .O(gate33inter3));
  inv1  gate1671(.a(s_161), .O(gate33inter4));
  nand2 gate1672(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate1673(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate1674(.a(G17), .O(gate33inter7));
  inv1  gate1675(.a(G21), .O(gate33inter8));
  nand2 gate1676(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate1677(.a(s_161), .b(gate33inter3), .O(gate33inter10));
  nor2  gate1678(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate1679(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate1680(.a(gate33inter12), .b(gate33inter1), .O(G338));
nand2 gate34( .a(G25), .b(G29), .O(G341) );

  xor2  gate743(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate744(.a(gate35inter0), .b(s_28), .O(gate35inter1));
  and2  gate745(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate746(.a(s_28), .O(gate35inter3));
  inv1  gate747(.a(s_29), .O(gate35inter4));
  nand2 gate748(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate749(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate750(.a(G18), .O(gate35inter7));
  inv1  gate751(.a(G22), .O(gate35inter8));
  nand2 gate752(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate753(.a(s_29), .b(gate35inter3), .O(gate35inter10));
  nor2  gate754(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate755(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate756(.a(gate35inter12), .b(gate35inter1), .O(G344));
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate1821(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate1822(.a(gate37inter0), .b(s_182), .O(gate37inter1));
  and2  gate1823(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate1824(.a(s_182), .O(gate37inter3));
  inv1  gate1825(.a(s_183), .O(gate37inter4));
  nand2 gate1826(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate1827(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate1828(.a(G19), .O(gate37inter7));
  inv1  gate1829(.a(G23), .O(gate37inter8));
  nand2 gate1830(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate1831(.a(s_183), .b(gate37inter3), .O(gate37inter10));
  nor2  gate1832(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate1833(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate1834(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate2605(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate2606(.a(gate39inter0), .b(s_294), .O(gate39inter1));
  and2  gate2607(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate2608(.a(s_294), .O(gate39inter3));
  inv1  gate2609(.a(s_295), .O(gate39inter4));
  nand2 gate2610(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate2611(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate2612(.a(G20), .O(gate39inter7));
  inv1  gate2613(.a(G24), .O(gate39inter8));
  nand2 gate2614(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate2615(.a(s_295), .b(gate39inter3), .O(gate39inter10));
  nor2  gate2616(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate2617(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate2618(.a(gate39inter12), .b(gate39inter1), .O(G356));

  xor2  gate2549(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate2550(.a(gate40inter0), .b(s_286), .O(gate40inter1));
  and2  gate2551(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate2552(.a(s_286), .O(gate40inter3));
  inv1  gate2553(.a(s_287), .O(gate40inter4));
  nand2 gate2554(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate2555(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate2556(.a(G28), .O(gate40inter7));
  inv1  gate2557(.a(G32), .O(gate40inter8));
  nand2 gate2558(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate2559(.a(s_287), .b(gate40inter3), .O(gate40inter10));
  nor2  gate2560(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate2561(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate2562(.a(gate40inter12), .b(gate40inter1), .O(G359));

  xor2  gate2689(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate2690(.a(gate41inter0), .b(s_306), .O(gate41inter1));
  and2  gate2691(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate2692(.a(s_306), .O(gate41inter3));
  inv1  gate2693(.a(s_307), .O(gate41inter4));
  nand2 gate2694(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate2695(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate2696(.a(G1), .O(gate41inter7));
  inv1  gate2697(.a(G266), .O(gate41inter8));
  nand2 gate2698(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate2699(.a(s_307), .b(gate41inter3), .O(gate41inter10));
  nor2  gate2700(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate2701(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate2702(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate1261(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate1262(.a(gate43inter0), .b(s_102), .O(gate43inter1));
  and2  gate1263(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate1264(.a(s_102), .O(gate43inter3));
  inv1  gate1265(.a(s_103), .O(gate43inter4));
  nand2 gate1266(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate1267(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate1268(.a(G3), .O(gate43inter7));
  inv1  gate1269(.a(G269), .O(gate43inter8));
  nand2 gate1270(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate1271(.a(s_103), .b(gate43inter3), .O(gate43inter10));
  nor2  gate1272(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate1273(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate1274(.a(gate43inter12), .b(gate43inter1), .O(G364));

  xor2  gate1513(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate1514(.a(gate44inter0), .b(s_138), .O(gate44inter1));
  and2  gate1515(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate1516(.a(s_138), .O(gate44inter3));
  inv1  gate1517(.a(s_139), .O(gate44inter4));
  nand2 gate1518(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate1519(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate1520(.a(G4), .O(gate44inter7));
  inv1  gate1521(.a(G269), .O(gate44inter8));
  nand2 gate1522(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate1523(.a(s_139), .b(gate44inter3), .O(gate44inter10));
  nor2  gate1524(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate1525(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate1526(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );

  xor2  gate2997(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate2998(.a(gate47inter0), .b(s_350), .O(gate47inter1));
  and2  gate2999(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate3000(.a(s_350), .O(gate47inter3));
  inv1  gate3001(.a(s_351), .O(gate47inter4));
  nand2 gate3002(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate3003(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate3004(.a(G7), .O(gate47inter7));
  inv1  gate3005(.a(G275), .O(gate47inter8));
  nand2 gate3006(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate3007(.a(s_351), .b(gate47inter3), .O(gate47inter10));
  nor2  gate3008(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate3009(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate3010(.a(gate47inter12), .b(gate47inter1), .O(G368));

  xor2  gate2815(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate2816(.a(gate48inter0), .b(s_324), .O(gate48inter1));
  and2  gate2817(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate2818(.a(s_324), .O(gate48inter3));
  inv1  gate2819(.a(s_325), .O(gate48inter4));
  nand2 gate2820(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate2821(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate2822(.a(G8), .O(gate48inter7));
  inv1  gate2823(.a(G275), .O(gate48inter8));
  nand2 gate2824(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate2825(.a(s_325), .b(gate48inter3), .O(gate48inter10));
  nor2  gate2826(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate2827(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate2828(.a(gate48inter12), .b(gate48inter1), .O(G369));

  xor2  gate1779(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate1780(.a(gate49inter0), .b(s_176), .O(gate49inter1));
  and2  gate1781(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate1782(.a(s_176), .O(gate49inter3));
  inv1  gate1783(.a(s_177), .O(gate49inter4));
  nand2 gate1784(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate1785(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate1786(.a(G9), .O(gate49inter7));
  inv1  gate1787(.a(G278), .O(gate49inter8));
  nand2 gate1788(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate1789(.a(s_177), .b(gate49inter3), .O(gate49inter10));
  nor2  gate1790(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate1791(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate1792(.a(gate49inter12), .b(gate49inter1), .O(G370));

  xor2  gate2115(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate2116(.a(gate50inter0), .b(s_224), .O(gate50inter1));
  and2  gate2117(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate2118(.a(s_224), .O(gate50inter3));
  inv1  gate2119(.a(s_225), .O(gate50inter4));
  nand2 gate2120(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate2121(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate2122(.a(G10), .O(gate50inter7));
  inv1  gate2123(.a(G278), .O(gate50inter8));
  nand2 gate2124(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate2125(.a(s_225), .b(gate50inter3), .O(gate50inter10));
  nor2  gate2126(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate2127(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate2128(.a(gate50inter12), .b(gate50inter1), .O(G371));
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate2129(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate2130(.a(gate52inter0), .b(s_226), .O(gate52inter1));
  and2  gate2131(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate2132(.a(s_226), .O(gate52inter3));
  inv1  gate2133(.a(s_227), .O(gate52inter4));
  nand2 gate2134(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate2135(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate2136(.a(G12), .O(gate52inter7));
  inv1  gate2137(.a(G281), .O(gate52inter8));
  nand2 gate2138(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate2139(.a(s_227), .b(gate52inter3), .O(gate52inter10));
  nor2  gate2140(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate2141(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate2142(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate1891(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate1892(.a(gate55inter0), .b(s_192), .O(gate55inter1));
  and2  gate1893(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate1894(.a(s_192), .O(gate55inter3));
  inv1  gate1895(.a(s_193), .O(gate55inter4));
  nand2 gate1896(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate1897(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate1898(.a(G15), .O(gate55inter7));
  inv1  gate1899(.a(G287), .O(gate55inter8));
  nand2 gate1900(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate1901(.a(s_193), .b(gate55inter3), .O(gate55inter10));
  nor2  gate1902(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate1903(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate1904(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate827(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate828(.a(gate57inter0), .b(s_40), .O(gate57inter1));
  and2  gate829(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate830(.a(s_40), .O(gate57inter3));
  inv1  gate831(.a(s_41), .O(gate57inter4));
  nand2 gate832(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate833(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate834(.a(G17), .O(gate57inter7));
  inv1  gate835(.a(G290), .O(gate57inter8));
  nand2 gate836(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate837(.a(s_41), .b(gate57inter3), .O(gate57inter10));
  nor2  gate838(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate839(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate840(.a(gate57inter12), .b(gate57inter1), .O(G378));
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate1653(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate1654(.a(gate59inter0), .b(s_158), .O(gate59inter1));
  and2  gate1655(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate1656(.a(s_158), .O(gate59inter3));
  inv1  gate1657(.a(s_159), .O(gate59inter4));
  nand2 gate1658(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate1659(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate1660(.a(G19), .O(gate59inter7));
  inv1  gate1661(.a(G293), .O(gate59inter8));
  nand2 gate1662(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate1663(.a(s_159), .b(gate59inter3), .O(gate59inter10));
  nor2  gate1664(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate1665(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate1666(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate1051(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate1052(.a(gate63inter0), .b(s_72), .O(gate63inter1));
  and2  gate1053(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate1054(.a(s_72), .O(gate63inter3));
  inv1  gate1055(.a(s_73), .O(gate63inter4));
  nand2 gate1056(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate1057(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate1058(.a(G23), .O(gate63inter7));
  inv1  gate1059(.a(G299), .O(gate63inter8));
  nand2 gate1060(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate1061(.a(s_73), .b(gate63inter3), .O(gate63inter10));
  nor2  gate1062(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate1063(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate1064(.a(gate63inter12), .b(gate63inter1), .O(G384));

  xor2  gate1401(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate1402(.a(gate64inter0), .b(s_122), .O(gate64inter1));
  and2  gate1403(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate1404(.a(s_122), .O(gate64inter3));
  inv1  gate1405(.a(s_123), .O(gate64inter4));
  nand2 gate1406(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate1407(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate1408(.a(G24), .O(gate64inter7));
  inv1  gate1409(.a(G299), .O(gate64inter8));
  nand2 gate1410(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate1411(.a(s_123), .b(gate64inter3), .O(gate64inter10));
  nor2  gate1412(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate1413(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate1414(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate2787(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate2788(.a(gate67inter0), .b(s_320), .O(gate67inter1));
  and2  gate2789(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate2790(.a(s_320), .O(gate67inter3));
  inv1  gate2791(.a(s_321), .O(gate67inter4));
  nand2 gate2792(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate2793(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate2794(.a(G27), .O(gate67inter7));
  inv1  gate2795(.a(G305), .O(gate67inter8));
  nand2 gate2796(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate2797(.a(s_321), .b(gate67inter3), .O(gate67inter10));
  nor2  gate2798(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate2799(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate2800(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate1275(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate1276(.a(gate69inter0), .b(s_104), .O(gate69inter1));
  and2  gate1277(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate1278(.a(s_104), .O(gate69inter3));
  inv1  gate1279(.a(s_105), .O(gate69inter4));
  nand2 gate1280(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate1281(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate1282(.a(G29), .O(gate69inter7));
  inv1  gate1283(.a(G308), .O(gate69inter8));
  nand2 gate1284(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate1285(.a(s_105), .b(gate69inter3), .O(gate69inter10));
  nor2  gate1286(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate1287(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate1288(.a(gate69inter12), .b(gate69inter1), .O(G390));

  xor2  gate2661(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate2662(.a(gate70inter0), .b(s_302), .O(gate70inter1));
  and2  gate2663(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate2664(.a(s_302), .O(gate70inter3));
  inv1  gate2665(.a(s_303), .O(gate70inter4));
  nand2 gate2666(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate2667(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate2668(.a(G30), .O(gate70inter7));
  inv1  gate2669(.a(G308), .O(gate70inter8));
  nand2 gate2670(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate2671(.a(s_303), .b(gate70inter3), .O(gate70inter10));
  nor2  gate2672(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate2673(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate2674(.a(gate70inter12), .b(gate70inter1), .O(G391));

  xor2  gate575(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate576(.a(gate71inter0), .b(s_4), .O(gate71inter1));
  and2  gate577(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate578(.a(s_4), .O(gate71inter3));
  inv1  gate579(.a(s_5), .O(gate71inter4));
  nand2 gate580(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate581(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate582(.a(G31), .O(gate71inter7));
  inv1  gate583(.a(G311), .O(gate71inter8));
  nand2 gate584(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate585(.a(s_5), .b(gate71inter3), .O(gate71inter10));
  nor2  gate586(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate587(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate588(.a(gate71inter12), .b(gate71inter1), .O(G392));

  xor2  gate1317(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate1318(.a(gate72inter0), .b(s_110), .O(gate72inter1));
  and2  gate1319(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate1320(.a(s_110), .O(gate72inter3));
  inv1  gate1321(.a(s_111), .O(gate72inter4));
  nand2 gate1322(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate1323(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate1324(.a(G32), .O(gate72inter7));
  inv1  gate1325(.a(G311), .O(gate72inter8));
  nand2 gate1326(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate1327(.a(s_111), .b(gate72inter3), .O(gate72inter10));
  nor2  gate1328(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate1329(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate1330(.a(gate72inter12), .b(gate72inter1), .O(G393));
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate2745(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate2746(.a(gate74inter0), .b(s_314), .O(gate74inter1));
  and2  gate2747(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate2748(.a(s_314), .O(gate74inter3));
  inv1  gate2749(.a(s_315), .O(gate74inter4));
  nand2 gate2750(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate2751(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate2752(.a(G5), .O(gate74inter7));
  inv1  gate2753(.a(G314), .O(gate74inter8));
  nand2 gate2754(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate2755(.a(s_315), .b(gate74inter3), .O(gate74inter10));
  nor2  gate2756(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate2757(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate2758(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );

  xor2  gate2927(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate2928(.a(gate76inter0), .b(s_340), .O(gate76inter1));
  and2  gate2929(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate2930(.a(s_340), .O(gate76inter3));
  inv1  gate2931(.a(s_341), .O(gate76inter4));
  nand2 gate2932(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate2933(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate2934(.a(G13), .O(gate76inter7));
  inv1  gate2935(.a(G317), .O(gate76inter8));
  nand2 gate2936(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate2937(.a(s_341), .b(gate76inter3), .O(gate76inter10));
  nor2  gate2938(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate2939(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate2940(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate2507(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate2508(.a(gate78inter0), .b(s_280), .O(gate78inter1));
  and2  gate2509(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate2510(.a(s_280), .O(gate78inter3));
  inv1  gate2511(.a(s_281), .O(gate78inter4));
  nand2 gate2512(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate2513(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate2514(.a(G6), .O(gate78inter7));
  inv1  gate2515(.a(G320), .O(gate78inter8));
  nand2 gate2516(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate2517(.a(s_281), .b(gate78inter3), .O(gate78inter10));
  nor2  gate2518(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate2519(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate2520(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate1149(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate1150(.a(gate81inter0), .b(s_86), .O(gate81inter1));
  and2  gate1151(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate1152(.a(s_86), .O(gate81inter3));
  inv1  gate1153(.a(s_87), .O(gate81inter4));
  nand2 gate1154(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate1155(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate1156(.a(G3), .O(gate81inter7));
  inv1  gate1157(.a(G326), .O(gate81inter8));
  nand2 gate1158(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate1159(.a(s_87), .b(gate81inter3), .O(gate81inter10));
  nor2  gate1160(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate1161(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate1162(.a(gate81inter12), .b(gate81inter1), .O(G402));

  xor2  gate2675(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate2676(.a(gate82inter0), .b(s_304), .O(gate82inter1));
  and2  gate2677(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate2678(.a(s_304), .O(gate82inter3));
  inv1  gate2679(.a(s_305), .O(gate82inter4));
  nand2 gate2680(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate2681(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate2682(.a(G7), .O(gate82inter7));
  inv1  gate2683(.a(G326), .O(gate82inter8));
  nand2 gate2684(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate2685(.a(s_305), .b(gate82inter3), .O(gate82inter10));
  nor2  gate2686(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate2687(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate2688(.a(gate82inter12), .b(gate82inter1), .O(G403));

  xor2  gate2451(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate2452(.a(gate83inter0), .b(s_272), .O(gate83inter1));
  and2  gate2453(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate2454(.a(s_272), .O(gate83inter3));
  inv1  gate2455(.a(s_273), .O(gate83inter4));
  nand2 gate2456(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate2457(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate2458(.a(G11), .O(gate83inter7));
  inv1  gate2459(.a(G329), .O(gate83inter8));
  nand2 gate2460(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate2461(.a(s_273), .b(gate83inter3), .O(gate83inter10));
  nor2  gate2462(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate2463(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate2464(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate1737(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate1738(.a(gate85inter0), .b(s_170), .O(gate85inter1));
  and2  gate1739(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate1740(.a(s_170), .O(gate85inter3));
  inv1  gate1741(.a(s_171), .O(gate85inter4));
  nand2 gate1742(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate1743(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate1744(.a(G4), .O(gate85inter7));
  inv1  gate1745(.a(G332), .O(gate85inter8));
  nand2 gate1746(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate1747(.a(s_171), .b(gate85inter3), .O(gate85inter10));
  nor2  gate1748(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate1749(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate1750(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );

  xor2  gate2087(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate2088(.a(gate89inter0), .b(s_220), .O(gate89inter1));
  and2  gate2089(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate2090(.a(s_220), .O(gate89inter3));
  inv1  gate2091(.a(s_221), .O(gate89inter4));
  nand2 gate2092(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate2093(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate2094(.a(G17), .O(gate89inter7));
  inv1  gate2095(.a(G338), .O(gate89inter8));
  nand2 gate2096(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate2097(.a(s_221), .b(gate89inter3), .O(gate89inter10));
  nor2  gate2098(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate2099(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate2100(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate1597(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate1598(.a(gate91inter0), .b(s_150), .O(gate91inter1));
  and2  gate1599(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate1600(.a(s_150), .O(gate91inter3));
  inv1  gate1601(.a(s_151), .O(gate91inter4));
  nand2 gate1602(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate1603(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate1604(.a(G25), .O(gate91inter7));
  inv1  gate1605(.a(G341), .O(gate91inter8));
  nand2 gate1606(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate1607(.a(s_151), .b(gate91inter3), .O(gate91inter10));
  nor2  gate1608(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate1609(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate1610(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );

  xor2  gate2871(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate2872(.a(gate93inter0), .b(s_332), .O(gate93inter1));
  and2  gate2873(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate2874(.a(s_332), .O(gate93inter3));
  inv1  gate2875(.a(s_333), .O(gate93inter4));
  nand2 gate2876(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate2877(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate2878(.a(G18), .O(gate93inter7));
  inv1  gate2879(.a(G344), .O(gate93inter8));
  nand2 gate2880(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate2881(.a(s_333), .b(gate93inter3), .O(gate93inter10));
  nor2  gate2882(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate2883(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate2884(.a(gate93inter12), .b(gate93inter1), .O(G414));
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate2101(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate2102(.a(gate95inter0), .b(s_222), .O(gate95inter1));
  and2  gate2103(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate2104(.a(s_222), .O(gate95inter3));
  inv1  gate2105(.a(s_223), .O(gate95inter4));
  nand2 gate2106(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate2107(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate2108(.a(G26), .O(gate95inter7));
  inv1  gate2109(.a(G347), .O(gate95inter8));
  nand2 gate2110(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate2111(.a(s_223), .b(gate95inter3), .O(gate95inter10));
  nor2  gate2112(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate2113(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate2114(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate2633(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate2634(.a(gate100inter0), .b(s_298), .O(gate100inter1));
  and2  gate2635(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate2636(.a(s_298), .O(gate100inter3));
  inv1  gate2637(.a(s_299), .O(gate100inter4));
  nand2 gate2638(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate2639(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate2640(.a(G31), .O(gate100inter7));
  inv1  gate2641(.a(G353), .O(gate100inter8));
  nand2 gate2642(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate2643(.a(s_299), .b(gate100inter3), .O(gate100inter10));
  nor2  gate2644(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate2645(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate2646(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );

  xor2  gate1877(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate1878(.a(gate103inter0), .b(s_190), .O(gate103inter1));
  and2  gate1879(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate1880(.a(s_190), .O(gate103inter3));
  inv1  gate1881(.a(s_191), .O(gate103inter4));
  nand2 gate1882(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate1883(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate1884(.a(G28), .O(gate103inter7));
  inv1  gate1885(.a(G359), .O(gate103inter8));
  nand2 gate1886(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate1887(.a(s_191), .b(gate103inter3), .O(gate103inter10));
  nor2  gate1888(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate1889(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate1890(.a(gate103inter12), .b(gate103inter1), .O(G424));
nand2 gate104( .a(G32), .b(G359), .O(G425) );

  xor2  gate1219(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate1220(.a(gate105inter0), .b(s_96), .O(gate105inter1));
  and2  gate1221(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate1222(.a(s_96), .O(gate105inter3));
  inv1  gate1223(.a(s_97), .O(gate105inter4));
  nand2 gate1224(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate1225(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate1226(.a(G362), .O(gate105inter7));
  inv1  gate1227(.a(G363), .O(gate105inter8));
  nand2 gate1228(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate1229(.a(s_97), .b(gate105inter3), .O(gate105inter10));
  nor2  gate1230(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate1231(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate1232(.a(gate105inter12), .b(gate105inter1), .O(G426));

  xor2  gate1527(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate1528(.a(gate106inter0), .b(s_140), .O(gate106inter1));
  and2  gate1529(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate1530(.a(s_140), .O(gate106inter3));
  inv1  gate1531(.a(s_141), .O(gate106inter4));
  nand2 gate1532(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate1533(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate1534(.a(G364), .O(gate106inter7));
  inv1  gate1535(.a(G365), .O(gate106inter8));
  nand2 gate1536(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate1537(.a(s_141), .b(gate106inter3), .O(gate106inter10));
  nor2  gate1538(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate1539(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate1540(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate2843(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate2844(.a(gate108inter0), .b(s_328), .O(gate108inter1));
  and2  gate2845(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate2846(.a(s_328), .O(gate108inter3));
  inv1  gate2847(.a(s_329), .O(gate108inter4));
  nand2 gate2848(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate2849(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate2850(.a(G368), .O(gate108inter7));
  inv1  gate2851(.a(G369), .O(gate108inter8));
  nand2 gate2852(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate2853(.a(s_329), .b(gate108inter3), .O(gate108inter10));
  nor2  gate2854(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate2855(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate2856(.a(gate108inter12), .b(gate108inter1), .O(G435));
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );

  xor2  gate1555(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate1556(.a(gate111inter0), .b(s_144), .O(gate111inter1));
  and2  gate1557(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate1558(.a(s_144), .O(gate111inter3));
  inv1  gate1559(.a(s_145), .O(gate111inter4));
  nand2 gate1560(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate1561(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate1562(.a(G374), .O(gate111inter7));
  inv1  gate1563(.a(G375), .O(gate111inter8));
  nand2 gate1564(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate1565(.a(s_145), .b(gate111inter3), .O(gate111inter10));
  nor2  gate1566(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate1567(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate1568(.a(gate111inter12), .b(gate111inter1), .O(G444));

  xor2  gate2367(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate2368(.a(gate112inter0), .b(s_260), .O(gate112inter1));
  and2  gate2369(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate2370(.a(s_260), .O(gate112inter3));
  inv1  gate2371(.a(s_261), .O(gate112inter4));
  nand2 gate2372(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate2373(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate2374(.a(G376), .O(gate112inter7));
  inv1  gate2375(.a(G377), .O(gate112inter8));
  nand2 gate2376(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate2377(.a(s_261), .b(gate112inter3), .O(gate112inter10));
  nor2  gate2378(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate2379(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate2380(.a(gate112inter12), .b(gate112inter1), .O(G447));

  xor2  gate3053(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate3054(.a(gate113inter0), .b(s_358), .O(gate113inter1));
  and2  gate3055(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate3056(.a(s_358), .O(gate113inter3));
  inv1  gate3057(.a(s_359), .O(gate113inter4));
  nand2 gate3058(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate3059(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate3060(.a(G378), .O(gate113inter7));
  inv1  gate3061(.a(G379), .O(gate113inter8));
  nand2 gate3062(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate3063(.a(s_359), .b(gate113inter3), .O(gate113inter10));
  nor2  gate3064(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate3065(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate3066(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate2395(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate2396(.a(gate121inter0), .b(s_264), .O(gate121inter1));
  and2  gate2397(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate2398(.a(s_264), .O(gate121inter3));
  inv1  gate2399(.a(s_265), .O(gate121inter4));
  nand2 gate2400(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate2401(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate2402(.a(G394), .O(gate121inter7));
  inv1  gate2403(.a(G395), .O(gate121inter8));
  nand2 gate2404(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate2405(.a(s_265), .b(gate121inter3), .O(gate121inter10));
  nor2  gate2406(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate2407(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate2408(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate1695(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate1696(.a(gate128inter0), .b(s_164), .O(gate128inter1));
  and2  gate1697(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate1698(.a(s_164), .O(gate128inter3));
  inv1  gate1699(.a(s_165), .O(gate128inter4));
  nand2 gate1700(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate1701(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate1702(.a(G408), .O(gate128inter7));
  inv1  gate1703(.a(G409), .O(gate128inter8));
  nand2 gate1704(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate1705(.a(s_165), .b(gate128inter3), .O(gate128inter10));
  nor2  gate1706(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate1707(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate1708(.a(gate128inter12), .b(gate128inter1), .O(G495));
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate561(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate562(.a(gate130inter0), .b(s_2), .O(gate130inter1));
  and2  gate563(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate564(.a(s_2), .O(gate130inter3));
  inv1  gate565(.a(s_3), .O(gate130inter4));
  nand2 gate566(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate567(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate568(.a(G412), .O(gate130inter7));
  inv1  gate569(.a(G413), .O(gate130inter8));
  nand2 gate570(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate571(.a(s_3), .b(gate130inter3), .O(gate130inter10));
  nor2  gate572(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate573(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate574(.a(gate130inter12), .b(gate130inter1), .O(G501));
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );

  xor2  gate645(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate646(.a(gate133inter0), .b(s_14), .O(gate133inter1));
  and2  gate647(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate648(.a(s_14), .O(gate133inter3));
  inv1  gate649(.a(s_15), .O(gate133inter4));
  nand2 gate650(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate651(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate652(.a(G418), .O(gate133inter7));
  inv1  gate653(.a(G419), .O(gate133inter8));
  nand2 gate654(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate655(.a(s_15), .b(gate133inter3), .O(gate133inter10));
  nor2  gate656(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate657(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate658(.a(gate133inter12), .b(gate133inter1), .O(G510));
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate1429(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate1430(.a(gate136inter0), .b(s_126), .O(gate136inter1));
  and2  gate1431(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate1432(.a(s_126), .O(gate136inter3));
  inv1  gate1433(.a(s_127), .O(gate136inter4));
  nand2 gate1434(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate1435(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate1436(.a(G424), .O(gate136inter7));
  inv1  gate1437(.a(G425), .O(gate136inter8));
  nand2 gate1438(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate1439(.a(s_127), .b(gate136inter3), .O(gate136inter10));
  nor2  gate1440(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate1441(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate1442(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate981(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate982(.a(gate138inter0), .b(s_62), .O(gate138inter1));
  and2  gate983(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate984(.a(s_62), .O(gate138inter3));
  inv1  gate985(.a(s_63), .O(gate138inter4));
  nand2 gate986(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate987(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate988(.a(G432), .O(gate138inter7));
  inv1  gate989(.a(G435), .O(gate138inter8));
  nand2 gate990(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate991(.a(s_63), .b(gate138inter3), .O(gate138inter10));
  nor2  gate992(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate993(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate994(.a(gate138inter12), .b(gate138inter1), .O(G525));

  xor2  gate2437(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate2438(.a(gate139inter0), .b(s_270), .O(gate139inter1));
  and2  gate2439(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate2440(.a(s_270), .O(gate139inter3));
  inv1  gate2441(.a(s_271), .O(gate139inter4));
  nand2 gate2442(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate2443(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate2444(.a(G438), .O(gate139inter7));
  inv1  gate2445(.a(G441), .O(gate139inter8));
  nand2 gate2446(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate2447(.a(s_271), .b(gate139inter3), .O(gate139inter10));
  nor2  gate2448(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate2449(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate2450(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate939(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate940(.a(gate141inter0), .b(s_56), .O(gate141inter1));
  and2  gate941(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate942(.a(s_56), .O(gate141inter3));
  inv1  gate943(.a(s_57), .O(gate141inter4));
  nand2 gate944(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate945(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate946(.a(G450), .O(gate141inter7));
  inv1  gate947(.a(G453), .O(gate141inter8));
  nand2 gate948(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate949(.a(s_57), .b(gate141inter3), .O(gate141inter10));
  nor2  gate950(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate951(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate952(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate2703(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate2704(.a(gate147inter0), .b(s_308), .O(gate147inter1));
  and2  gate2705(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate2706(.a(s_308), .O(gate147inter3));
  inv1  gate2707(.a(s_309), .O(gate147inter4));
  nand2 gate2708(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate2709(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate2710(.a(G486), .O(gate147inter7));
  inv1  gate2711(.a(G489), .O(gate147inter8));
  nand2 gate2712(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate2713(.a(s_309), .b(gate147inter3), .O(gate147inter10));
  nor2  gate2714(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate2715(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate2716(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate1583(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate1584(.a(gate149inter0), .b(s_148), .O(gate149inter1));
  and2  gate1585(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate1586(.a(s_148), .O(gate149inter3));
  inv1  gate1587(.a(s_149), .O(gate149inter4));
  nand2 gate1588(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate1589(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate1590(.a(G498), .O(gate149inter7));
  inv1  gate1591(.a(G501), .O(gate149inter8));
  nand2 gate1592(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate1593(.a(s_149), .b(gate149inter3), .O(gate149inter10));
  nor2  gate1594(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate1595(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate1596(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate589(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate590(.a(gate153inter0), .b(s_6), .O(gate153inter1));
  and2  gate591(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate592(.a(s_6), .O(gate153inter3));
  inv1  gate593(.a(s_7), .O(gate153inter4));
  nand2 gate594(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate595(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate596(.a(G426), .O(gate153inter7));
  inv1  gate597(.a(G522), .O(gate153inter8));
  nand2 gate598(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate599(.a(s_7), .b(gate153inter3), .O(gate153inter10));
  nor2  gate600(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate601(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate602(.a(gate153inter12), .b(gate153inter1), .O(G570));
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate2829(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate2830(.a(gate159inter0), .b(s_326), .O(gate159inter1));
  and2  gate2831(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate2832(.a(s_326), .O(gate159inter3));
  inv1  gate2833(.a(s_327), .O(gate159inter4));
  nand2 gate2834(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate2835(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate2836(.a(G444), .O(gate159inter7));
  inv1  gate2837(.a(G531), .O(gate159inter8));
  nand2 gate2838(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate2839(.a(s_327), .b(gate159inter3), .O(gate159inter10));
  nor2  gate2840(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate2841(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate2842(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate2227(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate2228(.a(gate161inter0), .b(s_240), .O(gate161inter1));
  and2  gate2229(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate2230(.a(s_240), .O(gate161inter3));
  inv1  gate2231(.a(s_241), .O(gate161inter4));
  nand2 gate2232(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate2233(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate2234(.a(G450), .O(gate161inter7));
  inv1  gate2235(.a(G534), .O(gate161inter8));
  nand2 gate2236(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate2237(.a(s_241), .b(gate161inter3), .O(gate161inter10));
  nor2  gate2238(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate2239(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate2240(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate673(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate674(.a(gate165inter0), .b(s_18), .O(gate165inter1));
  and2  gate675(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate676(.a(s_18), .O(gate165inter3));
  inv1  gate677(.a(s_19), .O(gate165inter4));
  nand2 gate678(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate679(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate680(.a(G462), .O(gate165inter7));
  inv1  gate681(.a(G540), .O(gate165inter8));
  nand2 gate682(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate683(.a(s_19), .b(gate165inter3), .O(gate165inter10));
  nor2  gate684(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate685(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate686(.a(gate165inter12), .b(gate165inter1), .O(G582));

  xor2  gate1849(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate1850(.a(gate166inter0), .b(s_186), .O(gate166inter1));
  and2  gate1851(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate1852(.a(s_186), .O(gate166inter3));
  inv1  gate1853(.a(s_187), .O(gate166inter4));
  nand2 gate1854(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate1855(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate1856(.a(G465), .O(gate166inter7));
  inv1  gate1857(.a(G540), .O(gate166inter8));
  nand2 gate1858(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate1859(.a(s_187), .b(gate166inter3), .O(gate166inter10));
  nor2  gate1860(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate1861(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate1862(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );

  xor2  gate687(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate688(.a(gate169inter0), .b(s_20), .O(gate169inter1));
  and2  gate689(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate690(.a(s_20), .O(gate169inter3));
  inv1  gate691(.a(s_21), .O(gate169inter4));
  nand2 gate692(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate693(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate694(.a(G474), .O(gate169inter7));
  inv1  gate695(.a(G546), .O(gate169inter8));
  nand2 gate696(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate697(.a(s_21), .b(gate169inter3), .O(gate169inter10));
  nor2  gate698(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate699(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate700(.a(gate169inter12), .b(gate169inter1), .O(G586));
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate631(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate632(.a(gate172inter0), .b(s_12), .O(gate172inter1));
  and2  gate633(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate634(.a(s_12), .O(gate172inter3));
  inv1  gate635(.a(s_13), .O(gate172inter4));
  nand2 gate636(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate637(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate638(.a(G483), .O(gate172inter7));
  inv1  gate639(.a(G549), .O(gate172inter8));
  nand2 gate640(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate641(.a(s_13), .b(gate172inter3), .O(gate172inter10));
  nor2  gate642(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate643(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate644(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate757(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate758(.a(gate183inter0), .b(s_30), .O(gate183inter1));
  and2  gate759(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate760(.a(s_30), .O(gate183inter3));
  inv1  gate761(.a(s_31), .O(gate183inter4));
  nand2 gate762(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate763(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate764(.a(G516), .O(gate183inter7));
  inv1  gate765(.a(G567), .O(gate183inter8));
  nand2 gate766(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate767(.a(s_31), .b(gate183inter3), .O(gate183inter10));
  nor2  gate768(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate769(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate770(.a(gate183inter12), .b(gate183inter1), .O(G600));

  xor2  gate2185(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate2186(.a(gate184inter0), .b(s_234), .O(gate184inter1));
  and2  gate2187(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate2188(.a(s_234), .O(gate184inter3));
  inv1  gate2189(.a(s_235), .O(gate184inter4));
  nand2 gate2190(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate2191(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate2192(.a(G519), .O(gate184inter7));
  inv1  gate2193(.a(G567), .O(gate184inter8));
  nand2 gate2194(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate2195(.a(s_235), .b(gate184inter3), .O(gate184inter10));
  nor2  gate2196(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate2197(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate2198(.a(gate184inter12), .b(gate184inter1), .O(G601));

  xor2  gate3011(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate3012(.a(gate185inter0), .b(s_352), .O(gate185inter1));
  and2  gate3013(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate3014(.a(s_352), .O(gate185inter3));
  inv1  gate3015(.a(s_353), .O(gate185inter4));
  nand2 gate3016(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate3017(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate3018(.a(G570), .O(gate185inter7));
  inv1  gate3019(.a(G571), .O(gate185inter8));
  nand2 gate3020(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate3021(.a(s_353), .b(gate185inter3), .O(gate185inter10));
  nor2  gate3022(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate3023(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate3024(.a(gate185inter12), .b(gate185inter1), .O(G602));
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate2983(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate2984(.a(gate190inter0), .b(s_348), .O(gate190inter1));
  and2  gate2985(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate2986(.a(s_348), .O(gate190inter3));
  inv1  gate2987(.a(s_349), .O(gate190inter4));
  nand2 gate2988(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate2989(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate2990(.a(G580), .O(gate190inter7));
  inv1  gate2991(.a(G581), .O(gate190inter8));
  nand2 gate2992(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate2993(.a(s_349), .b(gate190inter3), .O(gate190inter10));
  nor2  gate2994(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate2995(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate2996(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate2717(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate2718(.a(gate195inter0), .b(s_310), .O(gate195inter1));
  and2  gate2719(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate2720(.a(s_310), .O(gate195inter3));
  inv1  gate2721(.a(s_311), .O(gate195inter4));
  nand2 gate2722(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate2723(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate2724(.a(G590), .O(gate195inter7));
  inv1  gate2725(.a(G591), .O(gate195inter8));
  nand2 gate2726(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate2727(.a(s_311), .b(gate195inter3), .O(gate195inter10));
  nor2  gate2728(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate2729(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate2730(.a(gate195inter12), .b(gate195inter1), .O(G648));

  xor2  gate2955(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate2956(.a(gate196inter0), .b(s_344), .O(gate196inter1));
  and2  gate2957(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate2958(.a(s_344), .O(gate196inter3));
  inv1  gate2959(.a(s_345), .O(gate196inter4));
  nand2 gate2960(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate2961(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate2962(.a(G592), .O(gate196inter7));
  inv1  gate2963(.a(G593), .O(gate196inter8));
  nand2 gate2964(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate2965(.a(s_345), .b(gate196inter3), .O(gate196inter10));
  nor2  gate2966(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate2967(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate2968(.a(gate196inter12), .b(gate196inter1), .O(G651));

  xor2  gate1233(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate1234(.a(gate197inter0), .b(s_98), .O(gate197inter1));
  and2  gate1235(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate1236(.a(s_98), .O(gate197inter3));
  inv1  gate1237(.a(s_99), .O(gate197inter4));
  nand2 gate1238(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate1239(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate1240(.a(G594), .O(gate197inter7));
  inv1  gate1241(.a(G595), .O(gate197inter8));
  nand2 gate1242(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate1243(.a(s_99), .b(gate197inter3), .O(gate197inter10));
  nor2  gate1244(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate1245(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate1246(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );

  xor2  gate2255(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate2256(.a(gate199inter0), .b(s_244), .O(gate199inter1));
  and2  gate2257(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate2258(.a(s_244), .O(gate199inter3));
  inv1  gate2259(.a(s_245), .O(gate199inter4));
  nand2 gate2260(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate2261(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate2262(.a(G598), .O(gate199inter7));
  inv1  gate2263(.a(G599), .O(gate199inter8));
  nand2 gate2264(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate2265(.a(s_245), .b(gate199inter3), .O(gate199inter10));
  nor2  gate2266(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate2267(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate2268(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate995(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate996(.a(gate201inter0), .b(s_64), .O(gate201inter1));
  and2  gate997(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate998(.a(s_64), .O(gate201inter3));
  inv1  gate999(.a(s_65), .O(gate201inter4));
  nand2 gate1000(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate1001(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate1002(.a(G602), .O(gate201inter7));
  inv1  gate1003(.a(G607), .O(gate201inter8));
  nand2 gate1004(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate1005(.a(s_65), .b(gate201inter3), .O(gate201inter10));
  nor2  gate1006(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate1007(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate1008(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate2647(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate2648(.a(gate205inter0), .b(s_300), .O(gate205inter1));
  and2  gate2649(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate2650(.a(s_300), .O(gate205inter3));
  inv1  gate2651(.a(s_301), .O(gate205inter4));
  nand2 gate2652(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate2653(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate2654(.a(G622), .O(gate205inter7));
  inv1  gate2655(.a(G627), .O(gate205inter8));
  nand2 gate2656(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate2657(.a(s_301), .b(gate205inter3), .O(gate205inter10));
  nor2  gate2658(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate2659(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate2660(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );

  xor2  gate1541(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate1542(.a(gate209inter0), .b(s_142), .O(gate209inter1));
  and2  gate1543(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate1544(.a(s_142), .O(gate209inter3));
  inv1  gate1545(.a(s_143), .O(gate209inter4));
  nand2 gate1546(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate1547(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate1548(.a(G602), .O(gate209inter7));
  inv1  gate1549(.a(G666), .O(gate209inter8));
  nand2 gate1550(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate1551(.a(s_143), .b(gate209inter3), .O(gate209inter10));
  nor2  gate1552(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate1553(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate1554(.a(gate209inter12), .b(gate209inter1), .O(G690));
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );

  xor2  gate2353(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate2354(.a(gate212inter0), .b(s_258), .O(gate212inter1));
  and2  gate2355(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate2356(.a(s_258), .O(gate212inter3));
  inv1  gate2357(.a(s_259), .O(gate212inter4));
  nand2 gate2358(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate2359(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate2360(.a(G617), .O(gate212inter7));
  inv1  gate2361(.a(G669), .O(gate212inter8));
  nand2 gate2362(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate2363(.a(s_259), .b(gate212inter3), .O(gate212inter10));
  nor2  gate2364(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate2365(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate2366(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate1807(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate1808(.a(gate215inter0), .b(s_180), .O(gate215inter1));
  and2  gate1809(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate1810(.a(s_180), .O(gate215inter3));
  inv1  gate1811(.a(s_181), .O(gate215inter4));
  nand2 gate1812(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate1813(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate1814(.a(G607), .O(gate215inter7));
  inv1  gate1815(.a(G675), .O(gate215inter8));
  nand2 gate1816(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate1817(.a(s_181), .b(gate215inter3), .O(gate215inter10));
  nor2  gate1818(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate1819(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate1820(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate1205(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate1206(.a(gate219inter0), .b(s_94), .O(gate219inter1));
  and2  gate1207(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate1208(.a(s_94), .O(gate219inter3));
  inv1  gate1209(.a(s_95), .O(gate219inter4));
  nand2 gate1210(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate1211(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate1212(.a(G632), .O(gate219inter7));
  inv1  gate1213(.a(G681), .O(gate219inter8));
  nand2 gate1214(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate1215(.a(s_95), .b(gate219inter3), .O(gate219inter10));
  nor2  gate1216(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate1217(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate1218(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate2045(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate2046(.a(gate223inter0), .b(s_214), .O(gate223inter1));
  and2  gate2047(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate2048(.a(s_214), .O(gate223inter3));
  inv1  gate2049(.a(s_215), .O(gate223inter4));
  nand2 gate2050(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate2051(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate2052(.a(G627), .O(gate223inter7));
  inv1  gate2053(.a(G687), .O(gate223inter8));
  nand2 gate2054(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate2055(.a(s_215), .b(gate223inter3), .O(gate223inter10));
  nor2  gate2056(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate2057(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate2058(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate2059(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate2060(.a(gate227inter0), .b(s_216), .O(gate227inter1));
  and2  gate2061(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate2062(.a(s_216), .O(gate227inter3));
  inv1  gate2063(.a(s_217), .O(gate227inter4));
  nand2 gate2064(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate2065(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate2066(.a(G694), .O(gate227inter7));
  inv1  gate2067(.a(G695), .O(gate227inter8));
  nand2 gate2068(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate2069(.a(s_217), .b(gate227inter3), .O(gate227inter10));
  nor2  gate2070(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate2071(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate2072(.a(gate227inter12), .b(gate227inter1), .O(G712));
nand2 gate228( .a(G696), .b(G697), .O(G715) );

  xor2  gate2591(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate2592(.a(gate229inter0), .b(s_292), .O(gate229inter1));
  and2  gate2593(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate2594(.a(s_292), .O(gate229inter3));
  inv1  gate2595(.a(s_293), .O(gate229inter4));
  nand2 gate2596(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate2597(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate2598(.a(G698), .O(gate229inter7));
  inv1  gate2599(.a(G699), .O(gate229inter8));
  nand2 gate2600(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate2601(.a(s_293), .b(gate229inter3), .O(gate229inter10));
  nor2  gate2602(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate2603(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate2604(.a(gate229inter12), .b(gate229inter1), .O(G718));

  xor2  gate1793(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate1794(.a(gate230inter0), .b(s_178), .O(gate230inter1));
  and2  gate1795(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate1796(.a(s_178), .O(gate230inter3));
  inv1  gate1797(.a(s_179), .O(gate230inter4));
  nand2 gate1798(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate1799(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate1800(.a(G700), .O(gate230inter7));
  inv1  gate1801(.a(G701), .O(gate230inter8));
  nand2 gate1802(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate1803(.a(s_179), .b(gate230inter3), .O(gate230inter10));
  nor2  gate1804(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate1805(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate1806(.a(gate230inter12), .b(gate230inter1), .O(G721));

  xor2  gate659(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate660(.a(gate231inter0), .b(s_16), .O(gate231inter1));
  and2  gate661(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate662(.a(s_16), .O(gate231inter3));
  inv1  gate663(.a(s_17), .O(gate231inter4));
  nand2 gate664(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate665(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate666(.a(G702), .O(gate231inter7));
  inv1  gate667(.a(G703), .O(gate231inter8));
  nand2 gate668(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate669(.a(s_17), .b(gate231inter3), .O(gate231inter10));
  nor2  gate670(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate671(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate672(.a(gate231inter12), .b(gate231inter1), .O(G724));

  xor2  gate1569(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate1570(.a(gate232inter0), .b(s_146), .O(gate232inter1));
  and2  gate1571(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate1572(.a(s_146), .O(gate232inter3));
  inv1  gate1573(.a(s_147), .O(gate232inter4));
  nand2 gate1574(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate1575(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate1576(.a(G704), .O(gate232inter7));
  inv1  gate1577(.a(G705), .O(gate232inter8));
  nand2 gate1578(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate1579(.a(s_147), .b(gate232inter3), .O(gate232inter10));
  nor2  gate1580(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate1581(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate1582(.a(gate232inter12), .b(gate232inter1), .O(G727));

  xor2  gate2969(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate2970(.a(gate233inter0), .b(s_346), .O(gate233inter1));
  and2  gate2971(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate2972(.a(s_346), .O(gate233inter3));
  inv1  gate2973(.a(s_347), .O(gate233inter4));
  nand2 gate2974(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate2975(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate2976(.a(G242), .O(gate233inter7));
  inv1  gate2977(.a(G718), .O(gate233inter8));
  nand2 gate2978(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate2979(.a(s_347), .b(gate233inter3), .O(gate233inter10));
  nor2  gate2980(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate2981(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate2982(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );

  xor2  gate2409(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate2410(.a(gate235inter0), .b(s_266), .O(gate235inter1));
  and2  gate2411(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate2412(.a(s_266), .O(gate235inter3));
  inv1  gate2413(.a(s_267), .O(gate235inter4));
  nand2 gate2414(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate2415(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate2416(.a(G248), .O(gate235inter7));
  inv1  gate2417(.a(G724), .O(gate235inter8));
  nand2 gate2418(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate2419(.a(s_267), .b(gate235inter3), .O(gate235inter10));
  nor2  gate2420(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate2421(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate2422(.a(gate235inter12), .b(gate235inter1), .O(G736));

  xor2  gate2325(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate2326(.a(gate236inter0), .b(s_254), .O(gate236inter1));
  and2  gate2327(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate2328(.a(s_254), .O(gate236inter3));
  inv1  gate2329(.a(s_255), .O(gate236inter4));
  nand2 gate2330(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate2331(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate2332(.a(G251), .O(gate236inter7));
  inv1  gate2333(.a(G727), .O(gate236inter8));
  nand2 gate2334(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate2335(.a(s_255), .b(gate236inter3), .O(gate236inter10));
  nor2  gate2336(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate2337(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate2338(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );

  xor2  gate967(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate968(.a(gate238inter0), .b(s_60), .O(gate238inter1));
  and2  gate969(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate970(.a(s_60), .O(gate238inter3));
  inv1  gate971(.a(s_61), .O(gate238inter4));
  nand2 gate972(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate973(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate974(.a(G257), .O(gate238inter7));
  inv1  gate975(.a(G709), .O(gate238inter8));
  nand2 gate976(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate977(.a(s_61), .b(gate238inter3), .O(gate238inter10));
  nor2  gate978(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate979(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate980(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate1331(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate1332(.a(gate240inter0), .b(s_112), .O(gate240inter1));
  and2  gate1333(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate1334(.a(s_112), .O(gate240inter3));
  inv1  gate1335(.a(s_113), .O(gate240inter4));
  nand2 gate1336(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate1337(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate1338(.a(G263), .O(gate240inter7));
  inv1  gate1339(.a(G715), .O(gate240inter8));
  nand2 gate1340(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate1341(.a(s_113), .b(gate240inter3), .O(gate240inter10));
  nor2  gate1342(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate1343(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate1344(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate1485(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1486(.a(gate243inter0), .b(s_134), .O(gate243inter1));
  and2  gate1487(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1488(.a(s_134), .O(gate243inter3));
  inv1  gate1489(.a(s_135), .O(gate243inter4));
  nand2 gate1490(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1491(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1492(.a(G245), .O(gate243inter7));
  inv1  gate1493(.a(G733), .O(gate243inter8));
  nand2 gate1494(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1495(.a(s_135), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1496(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1497(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1498(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );

  xor2  gate701(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate702(.a(gate247inter0), .b(s_22), .O(gate247inter1));
  and2  gate703(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate704(.a(s_22), .O(gate247inter3));
  inv1  gate705(.a(s_23), .O(gate247inter4));
  nand2 gate706(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate707(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate708(.a(G251), .O(gate247inter7));
  inv1  gate709(.a(G739), .O(gate247inter8));
  nand2 gate710(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate711(.a(s_23), .b(gate247inter3), .O(gate247inter10));
  nor2  gate712(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate713(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate714(.a(gate247inter12), .b(gate247inter1), .O(G760));
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate603(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate604(.a(gate250inter0), .b(s_8), .O(gate250inter1));
  and2  gate605(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate606(.a(s_8), .O(gate250inter3));
  inv1  gate607(.a(s_9), .O(gate250inter4));
  nand2 gate608(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate609(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate610(.a(G706), .O(gate250inter7));
  inv1  gate611(.a(G742), .O(gate250inter8));
  nand2 gate612(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate613(.a(s_9), .b(gate250inter3), .O(gate250inter10));
  nor2  gate614(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate615(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate616(.a(gate250inter12), .b(gate250inter1), .O(G763));

  xor2  gate2619(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate2620(.a(gate251inter0), .b(s_296), .O(gate251inter1));
  and2  gate2621(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate2622(.a(s_296), .O(gate251inter3));
  inv1  gate2623(.a(s_297), .O(gate251inter4));
  nand2 gate2624(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate2625(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate2626(.a(G257), .O(gate251inter7));
  inv1  gate2627(.a(G745), .O(gate251inter8));
  nand2 gate2628(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate2629(.a(s_297), .b(gate251inter3), .O(gate251inter10));
  nor2  gate2630(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate2631(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate2632(.a(gate251inter12), .b(gate251inter1), .O(G764));

  xor2  gate1079(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate1080(.a(gate252inter0), .b(s_76), .O(gate252inter1));
  and2  gate1081(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate1082(.a(s_76), .O(gate252inter3));
  inv1  gate1083(.a(s_77), .O(gate252inter4));
  nand2 gate1084(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate1085(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate1086(.a(G709), .O(gate252inter7));
  inv1  gate1087(.a(G745), .O(gate252inter8));
  nand2 gate1088(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate1089(.a(s_77), .b(gate252inter3), .O(gate252inter10));
  nor2  gate1090(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate1091(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate1092(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate715(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate716(.a(gate255inter0), .b(s_24), .O(gate255inter1));
  and2  gate717(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate718(.a(s_24), .O(gate255inter3));
  inv1  gate719(.a(s_25), .O(gate255inter4));
  nand2 gate720(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate721(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate722(.a(G263), .O(gate255inter7));
  inv1  gate723(.a(G751), .O(gate255inter8));
  nand2 gate724(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate725(.a(s_25), .b(gate255inter3), .O(gate255inter10));
  nor2  gate726(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate727(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate728(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate2941(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate2942(.a(gate257inter0), .b(s_342), .O(gate257inter1));
  and2  gate2943(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate2944(.a(s_342), .O(gate257inter3));
  inv1  gate2945(.a(s_343), .O(gate257inter4));
  nand2 gate2946(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate2947(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate2948(.a(G754), .O(gate257inter7));
  inv1  gate2949(.a(G755), .O(gate257inter8));
  nand2 gate2950(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate2951(.a(s_343), .b(gate257inter3), .O(gate257inter10));
  nor2  gate2952(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate2953(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate2954(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );

  xor2  gate1107(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate1108(.a(gate259inter0), .b(s_80), .O(gate259inter1));
  and2  gate1109(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate1110(.a(s_80), .O(gate259inter3));
  inv1  gate1111(.a(s_81), .O(gate259inter4));
  nand2 gate1112(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate1113(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate1114(.a(G758), .O(gate259inter7));
  inv1  gate1115(.a(G759), .O(gate259inter8));
  nand2 gate1116(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate1117(.a(s_81), .b(gate259inter3), .O(gate259inter10));
  nor2  gate1118(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate1119(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate1120(.a(gate259inter12), .b(gate259inter1), .O(G776));

  xor2  gate1023(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate1024(.a(gate260inter0), .b(s_68), .O(gate260inter1));
  and2  gate1025(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate1026(.a(s_68), .O(gate260inter3));
  inv1  gate1027(.a(s_69), .O(gate260inter4));
  nand2 gate1028(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate1029(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate1030(.a(G760), .O(gate260inter7));
  inv1  gate1031(.a(G761), .O(gate260inter8));
  nand2 gate1032(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate1033(.a(s_69), .b(gate260inter3), .O(gate260inter10));
  nor2  gate1034(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate1035(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate1036(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate2577(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate2578(.a(gate263inter0), .b(s_290), .O(gate263inter1));
  and2  gate2579(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate2580(.a(s_290), .O(gate263inter3));
  inv1  gate2581(.a(s_291), .O(gate263inter4));
  nand2 gate2582(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate2583(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate2584(.a(G766), .O(gate263inter7));
  inv1  gate2585(.a(G767), .O(gate263inter8));
  nand2 gate2586(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate2587(.a(s_291), .b(gate263inter3), .O(gate263inter10));
  nor2  gate2588(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate2589(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate2590(.a(gate263inter12), .b(gate263inter1), .O(G788));

  xor2  gate1373(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate1374(.a(gate264inter0), .b(s_118), .O(gate264inter1));
  and2  gate1375(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate1376(.a(s_118), .O(gate264inter3));
  inv1  gate1377(.a(s_119), .O(gate264inter4));
  nand2 gate1378(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate1379(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate1380(.a(G768), .O(gate264inter7));
  inv1  gate1381(.a(G769), .O(gate264inter8));
  nand2 gate1382(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate1383(.a(s_119), .b(gate264inter3), .O(gate264inter10));
  nor2  gate1384(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate1385(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate1386(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate2031(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate2032(.a(gate266inter0), .b(s_212), .O(gate266inter1));
  and2  gate2033(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate2034(.a(s_212), .O(gate266inter3));
  inv1  gate2035(.a(s_213), .O(gate266inter4));
  nand2 gate2036(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate2037(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate2038(.a(G645), .O(gate266inter7));
  inv1  gate2039(.a(G773), .O(gate266inter8));
  nand2 gate2040(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate2041(.a(s_213), .b(gate266inter3), .O(gate266inter10));
  nor2  gate2042(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate2043(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate2044(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate1709(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate1710(.a(gate268inter0), .b(s_166), .O(gate268inter1));
  and2  gate1711(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate1712(.a(s_166), .O(gate268inter3));
  inv1  gate1713(.a(s_167), .O(gate268inter4));
  nand2 gate1714(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1715(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1716(.a(G651), .O(gate268inter7));
  inv1  gate1717(.a(G779), .O(gate268inter8));
  nand2 gate1718(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1719(.a(s_167), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1720(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1721(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1722(.a(gate268inter12), .b(gate268inter1), .O(G803));

  xor2  gate3025(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate3026(.a(gate269inter0), .b(s_354), .O(gate269inter1));
  and2  gate3027(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate3028(.a(s_354), .O(gate269inter3));
  inv1  gate3029(.a(s_355), .O(gate269inter4));
  nand2 gate3030(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate3031(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate3032(.a(G654), .O(gate269inter7));
  inv1  gate3033(.a(G782), .O(gate269inter8));
  nand2 gate3034(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate3035(.a(s_355), .b(gate269inter3), .O(gate269inter10));
  nor2  gate3036(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate3037(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate3038(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate1135(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate1136(.a(gate271inter0), .b(s_84), .O(gate271inter1));
  and2  gate1137(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate1138(.a(s_84), .O(gate271inter3));
  inv1  gate1139(.a(s_85), .O(gate271inter4));
  nand2 gate1140(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate1141(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate1142(.a(G660), .O(gate271inter7));
  inv1  gate1143(.a(G788), .O(gate271inter8));
  nand2 gate1144(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate1145(.a(s_85), .b(gate271inter3), .O(gate271inter10));
  nor2  gate1146(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate1147(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate1148(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate771(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate772(.a(gate274inter0), .b(s_32), .O(gate274inter1));
  and2  gate773(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate774(.a(s_32), .O(gate274inter3));
  inv1  gate775(.a(s_33), .O(gate274inter4));
  nand2 gate776(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate777(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate778(.a(G770), .O(gate274inter7));
  inv1  gate779(.a(G794), .O(gate274inter8));
  nand2 gate780(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate781(.a(s_33), .b(gate274inter3), .O(gate274inter10));
  nor2  gate782(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate783(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate784(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate2535(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate2536(.a(gate278inter0), .b(s_284), .O(gate278inter1));
  and2  gate2537(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate2538(.a(s_284), .O(gate278inter3));
  inv1  gate2539(.a(s_285), .O(gate278inter4));
  nand2 gate2540(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate2541(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate2542(.a(G776), .O(gate278inter7));
  inv1  gate2543(.a(G800), .O(gate278inter8));
  nand2 gate2544(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate2545(.a(s_285), .b(gate278inter3), .O(gate278inter10));
  nor2  gate2546(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate2547(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate2548(.a(gate278inter12), .b(gate278inter1), .O(G823));

  xor2  gate911(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate912(.a(gate279inter0), .b(s_52), .O(gate279inter1));
  and2  gate913(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate914(.a(s_52), .O(gate279inter3));
  inv1  gate915(.a(s_53), .O(gate279inter4));
  nand2 gate916(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate917(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate918(.a(G651), .O(gate279inter7));
  inv1  gate919(.a(G803), .O(gate279inter8));
  nand2 gate920(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate921(.a(s_53), .b(gate279inter3), .O(gate279inter10));
  nor2  gate922(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate923(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate924(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate1471(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate1472(.a(gate283inter0), .b(s_132), .O(gate283inter1));
  and2  gate1473(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate1474(.a(s_132), .O(gate283inter3));
  inv1  gate1475(.a(s_133), .O(gate283inter4));
  nand2 gate1476(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate1477(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate1478(.a(G657), .O(gate283inter7));
  inv1  gate1479(.a(G809), .O(gate283inter8));
  nand2 gate1480(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate1481(.a(s_133), .b(gate283inter3), .O(gate283inter10));
  nor2  gate1482(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate1483(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate1484(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate1009(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate1010(.a(gate285inter0), .b(s_66), .O(gate285inter1));
  and2  gate1011(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate1012(.a(s_66), .O(gate285inter3));
  inv1  gate1013(.a(s_67), .O(gate285inter4));
  nand2 gate1014(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate1015(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate1016(.a(G660), .O(gate285inter7));
  inv1  gate1017(.a(G812), .O(gate285inter8));
  nand2 gate1018(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate1019(.a(s_67), .b(gate285inter3), .O(gate285inter10));
  nor2  gate1020(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate1021(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate1022(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate1247(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate1248(.a(gate287inter0), .b(s_100), .O(gate287inter1));
  and2  gate1249(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate1250(.a(s_100), .O(gate287inter3));
  inv1  gate1251(.a(s_101), .O(gate287inter4));
  nand2 gate1252(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate1253(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate1254(.a(G663), .O(gate287inter7));
  inv1  gate1255(.a(G815), .O(gate287inter8));
  nand2 gate1256(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate1257(.a(s_101), .b(gate287inter3), .O(gate287inter10));
  nor2  gate1258(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate1259(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate1260(.a(gate287inter12), .b(gate287inter1), .O(G832));

  xor2  gate1121(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate1122(.a(gate288inter0), .b(s_82), .O(gate288inter1));
  and2  gate1123(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate1124(.a(s_82), .O(gate288inter3));
  inv1  gate1125(.a(s_83), .O(gate288inter4));
  nand2 gate1126(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate1127(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate1128(.a(G791), .O(gate288inter7));
  inv1  gate1129(.a(G815), .O(gate288inter8));
  nand2 gate1130(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate1131(.a(s_83), .b(gate288inter3), .O(gate288inter10));
  nor2  gate1132(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate1133(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate1134(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate1625(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate1626(.a(gate294inter0), .b(s_154), .O(gate294inter1));
  and2  gate1627(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate1628(.a(s_154), .O(gate294inter3));
  inv1  gate1629(.a(s_155), .O(gate294inter4));
  nand2 gate1630(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate1631(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate1632(.a(G832), .O(gate294inter7));
  inv1  gate1633(.a(G833), .O(gate294inter8));
  nand2 gate1634(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate1635(.a(s_155), .b(gate294inter3), .O(gate294inter10));
  nor2  gate1636(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate1637(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate1638(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate1289(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate1290(.a(gate388inter0), .b(s_106), .O(gate388inter1));
  and2  gate1291(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate1292(.a(s_106), .O(gate388inter3));
  inv1  gate1293(.a(s_107), .O(gate388inter4));
  nand2 gate1294(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate1295(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate1296(.a(G2), .O(gate388inter7));
  inv1  gate1297(.a(G1039), .O(gate388inter8));
  nand2 gate1298(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate1299(.a(s_107), .b(gate388inter3), .O(gate388inter10));
  nor2  gate1300(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate1301(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate1302(.a(gate388inter12), .b(gate388inter1), .O(G1135));
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate2493(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate2494(.a(gate390inter0), .b(s_278), .O(gate390inter1));
  and2  gate2495(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate2496(.a(s_278), .O(gate390inter3));
  inv1  gate2497(.a(s_279), .O(gate390inter4));
  nand2 gate2498(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate2499(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate2500(.a(G4), .O(gate390inter7));
  inv1  gate2501(.a(G1045), .O(gate390inter8));
  nand2 gate2502(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate2503(.a(s_279), .b(gate390inter3), .O(gate390inter10));
  nor2  gate2504(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate2505(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate2506(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate1639(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate1640(.a(gate393inter0), .b(s_156), .O(gate393inter1));
  and2  gate1641(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate1642(.a(s_156), .O(gate393inter3));
  inv1  gate1643(.a(s_157), .O(gate393inter4));
  nand2 gate1644(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate1645(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate1646(.a(G7), .O(gate393inter7));
  inv1  gate1647(.a(G1054), .O(gate393inter8));
  nand2 gate1648(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate1649(.a(s_157), .b(gate393inter3), .O(gate393inter10));
  nor2  gate1650(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate1651(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate1652(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate2157(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate2158(.a(gate397inter0), .b(s_230), .O(gate397inter1));
  and2  gate2159(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate2160(.a(s_230), .O(gate397inter3));
  inv1  gate2161(.a(s_231), .O(gate397inter4));
  nand2 gate2162(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate2163(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate2164(.a(G11), .O(gate397inter7));
  inv1  gate2165(.a(G1066), .O(gate397inter8));
  nand2 gate2166(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate2167(.a(s_231), .b(gate397inter3), .O(gate397inter10));
  nor2  gate2168(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate2169(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate2170(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate897(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate898(.a(gate399inter0), .b(s_50), .O(gate399inter1));
  and2  gate899(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate900(.a(s_50), .O(gate399inter3));
  inv1  gate901(.a(s_51), .O(gate399inter4));
  nand2 gate902(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate903(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate904(.a(G13), .O(gate399inter7));
  inv1  gate905(.a(G1072), .O(gate399inter8));
  nand2 gate906(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate907(.a(s_51), .b(gate399inter3), .O(gate399inter10));
  nor2  gate908(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate909(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate910(.a(gate399inter12), .b(gate399inter1), .O(G1168));

  xor2  gate1387(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate1388(.a(gate400inter0), .b(s_120), .O(gate400inter1));
  and2  gate1389(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate1390(.a(s_120), .O(gate400inter3));
  inv1  gate1391(.a(s_121), .O(gate400inter4));
  nand2 gate1392(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate1393(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate1394(.a(G14), .O(gate400inter7));
  inv1  gate1395(.a(G1075), .O(gate400inter8));
  nand2 gate1396(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate1397(.a(s_121), .b(gate400inter3), .O(gate400inter10));
  nor2  gate1398(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate1399(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate1400(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate2423(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate2424(.a(gate402inter0), .b(s_268), .O(gate402inter1));
  and2  gate2425(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate2426(.a(s_268), .O(gate402inter3));
  inv1  gate2427(.a(s_269), .O(gate402inter4));
  nand2 gate2428(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate2429(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate2430(.a(G16), .O(gate402inter7));
  inv1  gate2431(.a(G1081), .O(gate402inter8));
  nand2 gate2432(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate2433(.a(s_269), .b(gate402inter3), .O(gate402inter10));
  nor2  gate2434(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate2435(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate2436(.a(gate402inter12), .b(gate402inter1), .O(G1177));
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );

  xor2  gate1681(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate1682(.a(gate404inter0), .b(s_162), .O(gate404inter1));
  and2  gate1683(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate1684(.a(s_162), .O(gate404inter3));
  inv1  gate1685(.a(s_163), .O(gate404inter4));
  nand2 gate1686(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate1687(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate1688(.a(G18), .O(gate404inter7));
  inv1  gate1689(.a(G1087), .O(gate404inter8));
  nand2 gate1690(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate1691(.a(s_163), .b(gate404inter3), .O(gate404inter10));
  nor2  gate1692(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate1693(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate1694(.a(gate404inter12), .b(gate404inter1), .O(G1183));
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate2381(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate2382(.a(gate406inter0), .b(s_262), .O(gate406inter1));
  and2  gate2383(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate2384(.a(s_262), .O(gate406inter3));
  inv1  gate2385(.a(s_263), .O(gate406inter4));
  nand2 gate2386(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate2387(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate2388(.a(G20), .O(gate406inter7));
  inv1  gate2389(.a(G1093), .O(gate406inter8));
  nand2 gate2390(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate2391(.a(s_263), .b(gate406inter3), .O(gate406inter10));
  nor2  gate2392(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate2393(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate2394(.a(gate406inter12), .b(gate406inter1), .O(G1189));

  xor2  gate1751(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate1752(.a(gate407inter0), .b(s_172), .O(gate407inter1));
  and2  gate1753(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate1754(.a(s_172), .O(gate407inter3));
  inv1  gate1755(.a(s_173), .O(gate407inter4));
  nand2 gate1756(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate1757(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate1758(.a(G21), .O(gate407inter7));
  inv1  gate1759(.a(G1096), .O(gate407inter8));
  nand2 gate1760(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate1761(.a(s_173), .b(gate407inter3), .O(gate407inter10));
  nor2  gate1762(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate1763(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate1764(.a(gate407inter12), .b(gate407inter1), .O(G1192));

  xor2  gate1947(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate1948(.a(gate408inter0), .b(s_200), .O(gate408inter1));
  and2  gate1949(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate1950(.a(s_200), .O(gate408inter3));
  inv1  gate1951(.a(s_201), .O(gate408inter4));
  nand2 gate1952(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate1953(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate1954(.a(G22), .O(gate408inter7));
  inv1  gate1955(.a(G1099), .O(gate408inter8));
  nand2 gate1956(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate1957(.a(s_201), .b(gate408inter3), .O(gate408inter10));
  nor2  gate1958(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate1959(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate1960(.a(gate408inter12), .b(gate408inter1), .O(G1195));
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate799(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate800(.a(gate410inter0), .b(s_36), .O(gate410inter1));
  and2  gate801(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate802(.a(s_36), .O(gate410inter3));
  inv1  gate803(.a(s_37), .O(gate410inter4));
  nand2 gate804(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate805(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate806(.a(G24), .O(gate410inter7));
  inv1  gate807(.a(G1105), .O(gate410inter8));
  nand2 gate808(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate809(.a(s_37), .b(gate410inter3), .O(gate410inter10));
  nor2  gate810(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate811(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate812(.a(gate410inter12), .b(gate410inter1), .O(G1201));

  xor2  gate2283(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate2284(.a(gate411inter0), .b(s_248), .O(gate411inter1));
  and2  gate2285(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate2286(.a(s_248), .O(gate411inter3));
  inv1  gate2287(.a(s_249), .O(gate411inter4));
  nand2 gate2288(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate2289(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate2290(.a(G25), .O(gate411inter7));
  inv1  gate2291(.a(G1108), .O(gate411inter8));
  nand2 gate2292(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate2293(.a(s_249), .b(gate411inter3), .O(gate411inter10));
  nor2  gate2294(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate2295(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate2296(.a(gate411inter12), .b(gate411inter1), .O(G1204));

  xor2  gate1611(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate1612(.a(gate412inter0), .b(s_152), .O(gate412inter1));
  and2  gate1613(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate1614(.a(s_152), .O(gate412inter3));
  inv1  gate1615(.a(s_153), .O(gate412inter4));
  nand2 gate1616(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate1617(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate1618(.a(G26), .O(gate412inter7));
  inv1  gate1619(.a(G1111), .O(gate412inter8));
  nand2 gate1620(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate1621(.a(s_153), .b(gate412inter3), .O(gate412inter10));
  nor2  gate1622(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate1623(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate1624(.a(gate412inter12), .b(gate412inter1), .O(G1207));

  xor2  gate1765(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate1766(.a(gate413inter0), .b(s_174), .O(gate413inter1));
  and2  gate1767(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate1768(.a(s_174), .O(gate413inter3));
  inv1  gate1769(.a(s_175), .O(gate413inter4));
  nand2 gate1770(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1771(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1772(.a(G27), .O(gate413inter7));
  inv1  gate1773(.a(G1114), .O(gate413inter8));
  nand2 gate1774(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1775(.a(s_175), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1776(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1777(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1778(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate841(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate842(.a(gate415inter0), .b(s_42), .O(gate415inter1));
  and2  gate843(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate844(.a(s_42), .O(gate415inter3));
  inv1  gate845(.a(s_43), .O(gate415inter4));
  nand2 gate846(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate847(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate848(.a(G29), .O(gate415inter7));
  inv1  gate849(.a(G1120), .O(gate415inter8));
  nand2 gate850(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate851(.a(s_43), .b(gate415inter3), .O(gate415inter10));
  nor2  gate852(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate853(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate854(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate3067(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate3068(.a(gate417inter0), .b(s_360), .O(gate417inter1));
  and2  gate3069(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate3070(.a(s_360), .O(gate417inter3));
  inv1  gate3071(.a(s_361), .O(gate417inter4));
  nand2 gate3072(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate3073(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate3074(.a(G31), .O(gate417inter7));
  inv1  gate3075(.a(G1126), .O(gate417inter8));
  nand2 gate3076(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate3077(.a(s_361), .b(gate417inter3), .O(gate417inter10));
  nor2  gate3078(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate3079(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate3080(.a(gate417inter12), .b(gate417inter1), .O(G1222));

  xor2  gate1303(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate1304(.a(gate418inter0), .b(s_108), .O(gate418inter1));
  and2  gate1305(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate1306(.a(s_108), .O(gate418inter3));
  inv1  gate1307(.a(s_109), .O(gate418inter4));
  nand2 gate1308(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate1309(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate1310(.a(G32), .O(gate418inter7));
  inv1  gate1311(.a(G1129), .O(gate418inter8));
  nand2 gate1312(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate1313(.a(s_109), .b(gate418inter3), .O(gate418inter10));
  nor2  gate1314(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate1315(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate1316(.a(gate418inter12), .b(gate418inter1), .O(G1225));

  xor2  gate1905(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate1906(.a(gate419inter0), .b(s_194), .O(gate419inter1));
  and2  gate1907(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate1908(.a(s_194), .O(gate419inter3));
  inv1  gate1909(.a(s_195), .O(gate419inter4));
  nand2 gate1910(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate1911(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate1912(.a(G1), .O(gate419inter7));
  inv1  gate1913(.a(G1132), .O(gate419inter8));
  nand2 gate1914(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate1915(.a(s_195), .b(gate419inter3), .O(gate419inter10));
  nor2  gate1916(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate1917(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate1918(.a(gate419inter12), .b(gate419inter1), .O(G1228));
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate1835(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate1836(.a(gate422inter0), .b(s_184), .O(gate422inter1));
  and2  gate1837(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate1838(.a(s_184), .O(gate422inter3));
  inv1  gate1839(.a(s_185), .O(gate422inter4));
  nand2 gate1840(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate1841(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate1842(.a(G1039), .O(gate422inter7));
  inv1  gate1843(.a(G1135), .O(gate422inter8));
  nand2 gate1844(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate1845(.a(s_185), .b(gate422inter3), .O(gate422inter10));
  nor2  gate1846(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate1847(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate1848(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );

  xor2  gate2857(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate2858(.a(gate424inter0), .b(s_330), .O(gate424inter1));
  and2  gate2859(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate2860(.a(s_330), .O(gate424inter3));
  inv1  gate2861(.a(s_331), .O(gate424inter4));
  nand2 gate2862(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate2863(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate2864(.a(G1042), .O(gate424inter7));
  inv1  gate2865(.a(G1138), .O(gate424inter8));
  nand2 gate2866(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate2867(.a(s_331), .b(gate424inter3), .O(gate424inter10));
  nor2  gate2868(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate2869(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate2870(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );

  xor2  gate729(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate730(.a(gate426inter0), .b(s_26), .O(gate426inter1));
  and2  gate731(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate732(.a(s_26), .O(gate426inter3));
  inv1  gate733(.a(s_27), .O(gate426inter4));
  nand2 gate734(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate735(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate736(.a(G1045), .O(gate426inter7));
  inv1  gate737(.a(G1141), .O(gate426inter8));
  nand2 gate738(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate739(.a(s_27), .b(gate426inter3), .O(gate426inter10));
  nor2  gate740(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate741(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate742(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );

  xor2  gate2465(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate2466(.a(gate429inter0), .b(s_274), .O(gate429inter1));
  and2  gate2467(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate2468(.a(s_274), .O(gate429inter3));
  inv1  gate2469(.a(s_275), .O(gate429inter4));
  nand2 gate2470(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate2471(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate2472(.a(G6), .O(gate429inter7));
  inv1  gate2473(.a(G1147), .O(gate429inter8));
  nand2 gate2474(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate2475(.a(s_275), .b(gate429inter3), .O(gate429inter10));
  nor2  gate2476(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate2477(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate2478(.a(gate429inter12), .b(gate429inter1), .O(G1238));

  xor2  gate1863(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate1864(.a(gate430inter0), .b(s_188), .O(gate430inter1));
  and2  gate1865(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate1866(.a(s_188), .O(gate430inter3));
  inv1  gate1867(.a(s_189), .O(gate430inter4));
  nand2 gate1868(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate1869(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate1870(.a(G1051), .O(gate430inter7));
  inv1  gate1871(.a(G1147), .O(gate430inter8));
  nand2 gate1872(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate1873(.a(s_189), .b(gate430inter3), .O(gate430inter10));
  nor2  gate1874(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate1875(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate1876(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate2759(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate2760(.a(gate432inter0), .b(s_316), .O(gate432inter1));
  and2  gate2761(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate2762(.a(s_316), .O(gate432inter3));
  inv1  gate2763(.a(s_317), .O(gate432inter4));
  nand2 gate2764(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate2765(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate2766(.a(G1054), .O(gate432inter7));
  inv1  gate2767(.a(G1150), .O(gate432inter8));
  nand2 gate2768(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate2769(.a(s_317), .b(gate432inter3), .O(gate432inter10));
  nor2  gate2770(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate2771(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate2772(.a(gate432inter12), .b(gate432inter1), .O(G1241));

  xor2  gate2521(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate2522(.a(gate433inter0), .b(s_282), .O(gate433inter1));
  and2  gate2523(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate2524(.a(s_282), .O(gate433inter3));
  inv1  gate2525(.a(s_283), .O(gate433inter4));
  nand2 gate2526(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate2527(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate2528(.a(G8), .O(gate433inter7));
  inv1  gate2529(.a(G1153), .O(gate433inter8));
  nand2 gate2530(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate2531(.a(s_283), .b(gate433inter3), .O(gate433inter10));
  nor2  gate2532(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate2533(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate2534(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate2213(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate2214(.a(gate435inter0), .b(s_238), .O(gate435inter1));
  and2  gate2215(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate2216(.a(s_238), .O(gate435inter3));
  inv1  gate2217(.a(s_239), .O(gate435inter4));
  nand2 gate2218(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate2219(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate2220(.a(G9), .O(gate435inter7));
  inv1  gate2221(.a(G1156), .O(gate435inter8));
  nand2 gate2222(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate2223(.a(s_239), .b(gate435inter3), .O(gate435inter10));
  nor2  gate2224(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate2225(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate2226(.a(gate435inter12), .b(gate435inter1), .O(G1244));

  xor2  gate813(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate814(.a(gate436inter0), .b(s_38), .O(gate436inter1));
  and2  gate815(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate816(.a(s_38), .O(gate436inter3));
  inv1  gate817(.a(s_39), .O(gate436inter4));
  nand2 gate818(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate819(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate820(.a(G1060), .O(gate436inter7));
  inv1  gate821(.a(G1156), .O(gate436inter8));
  nand2 gate822(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate823(.a(s_39), .b(gate436inter3), .O(gate436inter10));
  nor2  gate824(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate825(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate826(.a(gate436inter12), .b(gate436inter1), .O(G1245));

  xor2  gate1499(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate1500(.a(gate437inter0), .b(s_136), .O(gate437inter1));
  and2  gate1501(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate1502(.a(s_136), .O(gate437inter3));
  inv1  gate1503(.a(s_137), .O(gate437inter4));
  nand2 gate1504(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate1505(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate1506(.a(G10), .O(gate437inter7));
  inv1  gate1507(.a(G1159), .O(gate437inter8));
  nand2 gate1508(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate1509(.a(s_137), .b(gate437inter3), .O(gate437inter10));
  nor2  gate1510(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate1511(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate1512(.a(gate437inter12), .b(gate437inter1), .O(G1246));

  xor2  gate2479(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate2480(.a(gate438inter0), .b(s_276), .O(gate438inter1));
  and2  gate2481(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate2482(.a(s_276), .O(gate438inter3));
  inv1  gate2483(.a(s_277), .O(gate438inter4));
  nand2 gate2484(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate2485(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate2486(.a(G1063), .O(gate438inter7));
  inv1  gate2487(.a(G1159), .O(gate438inter8));
  nand2 gate2488(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate2489(.a(s_277), .b(gate438inter3), .O(gate438inter10));
  nor2  gate2490(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate2491(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate2492(.a(gate438inter12), .b(gate438inter1), .O(G1247));

  xor2  gate1933(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate1934(.a(gate439inter0), .b(s_198), .O(gate439inter1));
  and2  gate1935(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate1936(.a(s_198), .O(gate439inter3));
  inv1  gate1937(.a(s_199), .O(gate439inter4));
  nand2 gate1938(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate1939(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate1940(.a(G11), .O(gate439inter7));
  inv1  gate1941(.a(G1162), .O(gate439inter8));
  nand2 gate1942(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate1943(.a(s_199), .b(gate439inter3), .O(gate439inter10));
  nor2  gate1944(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate1945(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate1946(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate1065(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate1066(.a(gate442inter0), .b(s_74), .O(gate442inter1));
  and2  gate1067(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate1068(.a(s_74), .O(gate442inter3));
  inv1  gate1069(.a(s_75), .O(gate442inter4));
  nand2 gate1070(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate1071(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate1072(.a(G1069), .O(gate442inter7));
  inv1  gate1073(.a(G1165), .O(gate442inter8));
  nand2 gate1074(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate1075(.a(s_75), .b(gate442inter3), .O(gate442inter10));
  nor2  gate1076(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate1077(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate1078(.a(gate442inter12), .b(gate442inter1), .O(G1251));

  xor2  gate953(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate954(.a(gate443inter0), .b(s_58), .O(gate443inter1));
  and2  gate955(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate956(.a(s_58), .O(gate443inter3));
  inv1  gate957(.a(s_59), .O(gate443inter4));
  nand2 gate958(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate959(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate960(.a(G13), .O(gate443inter7));
  inv1  gate961(.a(G1168), .O(gate443inter8));
  nand2 gate962(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate963(.a(s_59), .b(gate443inter3), .O(gate443inter10));
  nor2  gate964(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate965(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate966(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );

  xor2  gate2563(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate2564(.a(gate447inter0), .b(s_288), .O(gate447inter1));
  and2  gate2565(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate2566(.a(s_288), .O(gate447inter3));
  inv1  gate2567(.a(s_289), .O(gate447inter4));
  nand2 gate2568(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate2569(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate2570(.a(G15), .O(gate447inter7));
  inv1  gate2571(.a(G1174), .O(gate447inter8));
  nand2 gate2572(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate2573(.a(s_289), .b(gate447inter3), .O(gate447inter10));
  nor2  gate2574(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate2575(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate2576(.a(gate447inter12), .b(gate447inter1), .O(G1256));
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );

  xor2  gate855(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate856(.a(gate450inter0), .b(s_44), .O(gate450inter1));
  and2  gate857(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate858(.a(s_44), .O(gate450inter3));
  inv1  gate859(.a(s_45), .O(gate450inter4));
  nand2 gate860(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate861(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate862(.a(G1081), .O(gate450inter7));
  inv1  gate863(.a(G1177), .O(gate450inter8));
  nand2 gate864(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate865(.a(s_45), .b(gate450inter3), .O(gate450inter10));
  nor2  gate866(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate867(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate868(.a(gate450inter12), .b(gate450inter1), .O(G1259));
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate1163(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate1164(.a(gate456inter0), .b(s_88), .O(gate456inter1));
  and2  gate1165(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate1166(.a(s_88), .O(gate456inter3));
  inv1  gate1167(.a(s_89), .O(gate456inter4));
  nand2 gate1168(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate1169(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate1170(.a(G1090), .O(gate456inter7));
  inv1  gate1171(.a(G1186), .O(gate456inter8));
  nand2 gate1172(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate1173(.a(s_89), .b(gate456inter3), .O(gate456inter10));
  nor2  gate1174(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate1175(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate1176(.a(gate456inter12), .b(gate456inter1), .O(G1265));

  xor2  gate2913(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate2914(.a(gate457inter0), .b(s_338), .O(gate457inter1));
  and2  gate2915(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate2916(.a(s_338), .O(gate457inter3));
  inv1  gate2917(.a(s_339), .O(gate457inter4));
  nand2 gate2918(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate2919(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate2920(.a(G20), .O(gate457inter7));
  inv1  gate2921(.a(G1189), .O(gate457inter8));
  nand2 gate2922(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate2923(.a(s_339), .b(gate457inter3), .O(gate457inter10));
  nor2  gate2924(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate2925(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate2926(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate617(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate618(.a(gate461inter0), .b(s_10), .O(gate461inter1));
  and2  gate619(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate620(.a(s_10), .O(gate461inter3));
  inv1  gate621(.a(s_11), .O(gate461inter4));
  nand2 gate622(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate623(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate624(.a(G22), .O(gate461inter7));
  inv1  gate625(.a(G1195), .O(gate461inter8));
  nand2 gate626(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate627(.a(s_11), .b(gate461inter3), .O(gate461inter10));
  nor2  gate628(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate629(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate630(.a(gate461inter12), .b(gate461inter1), .O(G1270));
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate1975(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate1976(.a(gate463inter0), .b(s_204), .O(gate463inter1));
  and2  gate1977(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate1978(.a(s_204), .O(gate463inter3));
  inv1  gate1979(.a(s_205), .O(gate463inter4));
  nand2 gate1980(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate1981(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate1982(.a(G23), .O(gate463inter7));
  inv1  gate1983(.a(G1198), .O(gate463inter8));
  nand2 gate1984(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate1985(.a(s_205), .b(gate463inter3), .O(gate463inter10));
  nor2  gate1986(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate1987(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate1988(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate2339(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate2340(.a(gate466inter0), .b(s_256), .O(gate466inter1));
  and2  gate2341(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate2342(.a(s_256), .O(gate466inter3));
  inv1  gate2343(.a(s_257), .O(gate466inter4));
  nand2 gate2344(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate2345(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate2346(.a(G1105), .O(gate466inter7));
  inv1  gate2347(.a(G1201), .O(gate466inter8));
  nand2 gate2348(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate2349(.a(s_257), .b(gate466inter3), .O(gate466inter10));
  nor2  gate2350(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate2351(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate2352(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate2143(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate2144(.a(gate471inter0), .b(s_228), .O(gate471inter1));
  and2  gate2145(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate2146(.a(s_228), .O(gate471inter3));
  inv1  gate2147(.a(s_229), .O(gate471inter4));
  nand2 gate2148(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate2149(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate2150(.a(G27), .O(gate471inter7));
  inv1  gate2151(.a(G1210), .O(gate471inter8));
  nand2 gate2152(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate2153(.a(s_229), .b(gate471inter3), .O(gate471inter10));
  nor2  gate2154(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate2155(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate2156(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate2801(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate2802(.a(gate477inter0), .b(s_322), .O(gate477inter1));
  and2  gate2803(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate2804(.a(s_322), .O(gate477inter3));
  inv1  gate2805(.a(s_323), .O(gate477inter4));
  nand2 gate2806(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate2807(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate2808(.a(G30), .O(gate477inter7));
  inv1  gate2809(.a(G1219), .O(gate477inter8));
  nand2 gate2810(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate2811(.a(s_323), .b(gate477inter3), .O(gate477inter10));
  nor2  gate2812(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate2813(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate2814(.a(gate477inter12), .b(gate477inter1), .O(G1286));

  xor2  gate925(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate926(.a(gate478inter0), .b(s_54), .O(gate478inter1));
  and2  gate927(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate928(.a(s_54), .O(gate478inter3));
  inv1  gate929(.a(s_55), .O(gate478inter4));
  nand2 gate930(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate931(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate932(.a(G1123), .O(gate478inter7));
  inv1  gate933(.a(G1219), .O(gate478inter8));
  nand2 gate934(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate935(.a(s_55), .b(gate478inter3), .O(gate478inter10));
  nor2  gate936(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate937(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate938(.a(gate478inter12), .b(gate478inter1), .O(G1287));

  xor2  gate2773(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate2774(.a(gate479inter0), .b(s_318), .O(gate479inter1));
  and2  gate2775(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate2776(.a(s_318), .O(gate479inter3));
  inv1  gate2777(.a(s_319), .O(gate479inter4));
  nand2 gate2778(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate2779(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate2780(.a(G31), .O(gate479inter7));
  inv1  gate2781(.a(G1222), .O(gate479inter8));
  nand2 gate2782(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate2783(.a(s_319), .b(gate479inter3), .O(gate479inter10));
  nor2  gate2784(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate2785(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate2786(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate3039(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate3040(.a(gate482inter0), .b(s_356), .O(gate482inter1));
  and2  gate3041(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate3042(.a(s_356), .O(gate482inter3));
  inv1  gate3043(.a(s_357), .O(gate482inter4));
  nand2 gate3044(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate3045(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate3046(.a(G1129), .O(gate482inter7));
  inv1  gate3047(.a(G1225), .O(gate482inter8));
  nand2 gate3048(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate3049(.a(s_357), .b(gate482inter3), .O(gate482inter10));
  nor2  gate3050(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate3051(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate3052(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );

  xor2  gate1919(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate1920(.a(gate484inter0), .b(s_196), .O(gate484inter1));
  and2  gate1921(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate1922(.a(s_196), .O(gate484inter3));
  inv1  gate1923(.a(s_197), .O(gate484inter4));
  nand2 gate1924(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate1925(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate1926(.a(G1230), .O(gate484inter7));
  inv1  gate1927(.a(G1231), .O(gate484inter8));
  nand2 gate1928(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate1929(.a(s_197), .b(gate484inter3), .O(gate484inter10));
  nor2  gate1930(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate1931(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate1932(.a(gate484inter12), .b(gate484inter1), .O(G1293));

  xor2  gate2199(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate2200(.a(gate485inter0), .b(s_236), .O(gate485inter1));
  and2  gate2201(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate2202(.a(s_236), .O(gate485inter3));
  inv1  gate2203(.a(s_237), .O(gate485inter4));
  nand2 gate2204(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate2205(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate2206(.a(G1232), .O(gate485inter7));
  inv1  gate2207(.a(G1233), .O(gate485inter8));
  nand2 gate2208(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate2209(.a(s_237), .b(gate485inter3), .O(gate485inter10));
  nor2  gate2210(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate2211(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate2212(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate2297(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate2298(.a(gate487inter0), .b(s_250), .O(gate487inter1));
  and2  gate2299(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate2300(.a(s_250), .O(gate487inter3));
  inv1  gate2301(.a(s_251), .O(gate487inter4));
  nand2 gate2302(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate2303(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate2304(.a(G1236), .O(gate487inter7));
  inv1  gate2305(.a(G1237), .O(gate487inter8));
  nand2 gate2306(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate2307(.a(s_251), .b(gate487inter3), .O(gate487inter10));
  nor2  gate2308(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate2309(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate2310(.a(gate487inter12), .b(gate487inter1), .O(G1296));

  xor2  gate1037(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate1038(.a(gate488inter0), .b(s_70), .O(gate488inter1));
  and2  gate1039(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate1040(.a(s_70), .O(gate488inter3));
  inv1  gate1041(.a(s_71), .O(gate488inter4));
  nand2 gate1042(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate1043(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate1044(.a(G1238), .O(gate488inter7));
  inv1  gate1045(.a(G1239), .O(gate488inter8));
  nand2 gate1046(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate1047(.a(s_71), .b(gate488inter3), .O(gate488inter10));
  nor2  gate1048(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate1049(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate1050(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate1359(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate1360(.a(gate493inter0), .b(s_116), .O(gate493inter1));
  and2  gate1361(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate1362(.a(s_116), .O(gate493inter3));
  inv1  gate1363(.a(s_117), .O(gate493inter4));
  nand2 gate1364(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate1365(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate1366(.a(G1248), .O(gate493inter7));
  inv1  gate1367(.a(G1249), .O(gate493inter8));
  nand2 gate1368(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate1369(.a(s_117), .b(gate493inter3), .O(gate493inter10));
  nor2  gate1370(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate1371(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate1372(.a(gate493inter12), .b(gate493inter1), .O(G1302));

  xor2  gate869(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate870(.a(gate494inter0), .b(s_46), .O(gate494inter1));
  and2  gate871(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate872(.a(s_46), .O(gate494inter3));
  inv1  gate873(.a(s_47), .O(gate494inter4));
  nand2 gate874(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate875(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate876(.a(G1250), .O(gate494inter7));
  inv1  gate877(.a(G1251), .O(gate494inter8));
  nand2 gate878(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate879(.a(s_47), .b(gate494inter3), .O(gate494inter10));
  nor2  gate880(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate881(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate882(.a(gate494inter12), .b(gate494inter1), .O(G1303));

  xor2  gate1191(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate1192(.a(gate495inter0), .b(s_92), .O(gate495inter1));
  and2  gate1193(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate1194(.a(s_92), .O(gate495inter3));
  inv1  gate1195(.a(s_93), .O(gate495inter4));
  nand2 gate1196(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate1197(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate1198(.a(G1252), .O(gate495inter7));
  inv1  gate1199(.a(G1253), .O(gate495inter8));
  nand2 gate1200(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate1201(.a(s_93), .b(gate495inter3), .O(gate495inter10));
  nor2  gate1202(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate1203(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate1204(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate2241(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate2242(.a(gate497inter0), .b(s_242), .O(gate497inter1));
  and2  gate2243(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate2244(.a(s_242), .O(gate497inter3));
  inv1  gate2245(.a(s_243), .O(gate497inter4));
  nand2 gate2246(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate2247(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate2248(.a(G1256), .O(gate497inter7));
  inv1  gate2249(.a(G1257), .O(gate497inter8));
  nand2 gate2250(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate2251(.a(s_243), .b(gate497inter3), .O(gate497inter10));
  nor2  gate2252(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate2253(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate2254(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate2731(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate2732(.a(gate499inter0), .b(s_312), .O(gate499inter1));
  and2  gate2733(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate2734(.a(s_312), .O(gate499inter3));
  inv1  gate2735(.a(s_313), .O(gate499inter4));
  nand2 gate2736(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate2737(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate2738(.a(G1260), .O(gate499inter7));
  inv1  gate2739(.a(G1261), .O(gate499inter8));
  nand2 gate2740(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate2741(.a(s_313), .b(gate499inter3), .O(gate499inter10));
  nor2  gate2742(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate2743(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate2744(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate1177(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate1178(.a(gate502inter0), .b(s_90), .O(gate502inter1));
  and2  gate1179(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate1180(.a(s_90), .O(gate502inter3));
  inv1  gate1181(.a(s_91), .O(gate502inter4));
  nand2 gate1182(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate1183(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate1184(.a(G1266), .O(gate502inter7));
  inv1  gate1185(.a(G1267), .O(gate502inter8));
  nand2 gate1186(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate1187(.a(s_91), .b(gate502inter3), .O(gate502inter10));
  nor2  gate1188(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate1189(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate1190(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate547(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate548(.a(gate509inter0), .b(s_0), .O(gate509inter1));
  and2  gate549(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate550(.a(s_0), .O(gate509inter3));
  inv1  gate551(.a(s_1), .O(gate509inter4));
  nand2 gate552(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate553(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate554(.a(G1280), .O(gate509inter7));
  inv1  gate555(.a(G1281), .O(gate509inter8));
  nand2 gate556(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate557(.a(s_1), .b(gate509inter3), .O(gate509inter10));
  nor2  gate558(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate559(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate560(.a(gate509inter12), .b(gate509inter1), .O(G1318));

  xor2  gate1723(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate1724(.a(gate510inter0), .b(s_168), .O(gate510inter1));
  and2  gate1725(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate1726(.a(s_168), .O(gate510inter3));
  inv1  gate1727(.a(s_169), .O(gate510inter4));
  nand2 gate1728(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate1729(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate1730(.a(G1282), .O(gate510inter7));
  inv1  gate1731(.a(G1283), .O(gate510inter8));
  nand2 gate1732(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate1733(.a(s_169), .b(gate510inter3), .O(gate510inter10));
  nor2  gate1734(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate1735(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate1736(.a(gate510inter12), .b(gate510inter1), .O(G1319));

  xor2  gate1093(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate1094(.a(gate511inter0), .b(s_78), .O(gate511inter1));
  and2  gate1095(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate1096(.a(s_78), .O(gate511inter3));
  inv1  gate1097(.a(s_79), .O(gate511inter4));
  nand2 gate1098(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate1099(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate1100(.a(G1284), .O(gate511inter7));
  inv1  gate1101(.a(G1285), .O(gate511inter8));
  nand2 gate1102(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate1103(.a(s_79), .b(gate511inter3), .O(gate511inter10));
  nor2  gate1104(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate1105(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate1106(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule