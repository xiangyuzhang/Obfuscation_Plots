module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate743(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate744(.a(gate20inter0), .b(s_28), .O(gate20inter1));
  and2  gate745(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate746(.a(s_28), .O(gate20inter3));
  inv1  gate747(.a(s_29), .O(gate20inter4));
  nand2 gate748(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate749(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate750(.a(G23), .O(gate20inter7));
  inv1  gate751(.a(G24), .O(gate20inter8));
  nand2 gate752(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate753(.a(s_29), .b(gate20inter3), .O(gate20inter10));
  nor2  gate754(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate755(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate756(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate1233(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate1234(.a(gate23inter0), .b(s_98), .O(gate23inter1));
  and2  gate1235(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate1236(.a(s_98), .O(gate23inter3));
  inv1  gate1237(.a(s_99), .O(gate23inter4));
  nand2 gate1238(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate1239(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate1240(.a(G29), .O(gate23inter7));
  inv1  gate1241(.a(G30), .O(gate23inter8));
  nand2 gate1242(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate1243(.a(s_99), .b(gate23inter3), .O(gate23inter10));
  nor2  gate1244(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate1245(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate1246(.a(gate23inter12), .b(gate23inter1), .O(G308));

  xor2  gate1961(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate1962(.a(gate24inter0), .b(s_202), .O(gate24inter1));
  and2  gate1963(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate1964(.a(s_202), .O(gate24inter3));
  inv1  gate1965(.a(s_203), .O(gate24inter4));
  nand2 gate1966(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate1967(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate1968(.a(G31), .O(gate24inter7));
  inv1  gate1969(.a(G32), .O(gate24inter8));
  nand2 gate1970(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate1971(.a(s_203), .b(gate24inter3), .O(gate24inter10));
  nor2  gate1972(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate1973(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate1974(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate1569(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate1570(.a(gate27inter0), .b(s_146), .O(gate27inter1));
  and2  gate1571(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate1572(.a(s_146), .O(gate27inter3));
  inv1  gate1573(.a(s_147), .O(gate27inter4));
  nand2 gate1574(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate1575(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate1576(.a(G2), .O(gate27inter7));
  inv1  gate1577(.a(G6), .O(gate27inter8));
  nand2 gate1578(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate1579(.a(s_147), .b(gate27inter3), .O(gate27inter10));
  nor2  gate1580(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate1581(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate1582(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate1135(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate1136(.a(gate33inter0), .b(s_84), .O(gate33inter1));
  and2  gate1137(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate1138(.a(s_84), .O(gate33inter3));
  inv1  gate1139(.a(s_85), .O(gate33inter4));
  nand2 gate1140(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate1141(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate1142(.a(G17), .O(gate33inter7));
  inv1  gate1143(.a(G21), .O(gate33inter8));
  nand2 gate1144(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate1145(.a(s_85), .b(gate33inter3), .O(gate33inter10));
  nor2  gate1146(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate1147(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate1148(.a(gate33inter12), .b(gate33inter1), .O(G338));
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate813(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate814(.a(gate39inter0), .b(s_38), .O(gate39inter1));
  and2  gate815(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate816(.a(s_38), .O(gate39inter3));
  inv1  gate817(.a(s_39), .O(gate39inter4));
  nand2 gate818(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate819(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate820(.a(G20), .O(gate39inter7));
  inv1  gate821(.a(G24), .O(gate39inter8));
  nand2 gate822(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate823(.a(s_39), .b(gate39inter3), .O(gate39inter10));
  nor2  gate824(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate825(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate826(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate785(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate786(.a(gate41inter0), .b(s_34), .O(gate41inter1));
  and2  gate787(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate788(.a(s_34), .O(gate41inter3));
  inv1  gate789(.a(s_35), .O(gate41inter4));
  nand2 gate790(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate791(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate792(.a(G1), .O(gate41inter7));
  inv1  gate793(.a(G266), .O(gate41inter8));
  nand2 gate794(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate795(.a(s_35), .b(gate41inter3), .O(gate41inter10));
  nor2  gate796(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate797(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate798(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate967(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate968(.a(gate51inter0), .b(s_60), .O(gate51inter1));
  and2  gate969(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate970(.a(s_60), .O(gate51inter3));
  inv1  gate971(.a(s_61), .O(gate51inter4));
  nand2 gate972(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate973(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate974(.a(G11), .O(gate51inter7));
  inv1  gate975(.a(G281), .O(gate51inter8));
  nand2 gate976(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate977(.a(s_61), .b(gate51inter3), .O(gate51inter10));
  nor2  gate978(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate979(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate980(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate2031(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate2032(.a(gate54inter0), .b(s_212), .O(gate54inter1));
  and2  gate2033(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate2034(.a(s_212), .O(gate54inter3));
  inv1  gate2035(.a(s_213), .O(gate54inter4));
  nand2 gate2036(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate2037(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate2038(.a(G14), .O(gate54inter7));
  inv1  gate2039(.a(G284), .O(gate54inter8));
  nand2 gate2040(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate2041(.a(s_213), .b(gate54inter3), .O(gate54inter10));
  nor2  gate2042(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate2043(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate2044(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate855(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate856(.a(gate60inter0), .b(s_44), .O(gate60inter1));
  and2  gate857(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate858(.a(s_44), .O(gate60inter3));
  inv1  gate859(.a(s_45), .O(gate60inter4));
  nand2 gate860(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate861(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate862(.a(G20), .O(gate60inter7));
  inv1  gate863(.a(G293), .O(gate60inter8));
  nand2 gate864(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate865(.a(s_45), .b(gate60inter3), .O(gate60inter10));
  nor2  gate866(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate867(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate868(.a(gate60inter12), .b(gate60inter1), .O(G381));

  xor2  gate2381(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate2382(.a(gate61inter0), .b(s_262), .O(gate61inter1));
  and2  gate2383(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate2384(.a(s_262), .O(gate61inter3));
  inv1  gate2385(.a(s_263), .O(gate61inter4));
  nand2 gate2386(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate2387(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate2388(.a(G21), .O(gate61inter7));
  inv1  gate2389(.a(G296), .O(gate61inter8));
  nand2 gate2390(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate2391(.a(s_263), .b(gate61inter3), .O(gate61inter10));
  nor2  gate2392(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate2393(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate2394(.a(gate61inter12), .b(gate61inter1), .O(G382));
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate2241(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate2242(.a(gate65inter0), .b(s_242), .O(gate65inter1));
  and2  gate2243(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate2244(.a(s_242), .O(gate65inter3));
  inv1  gate2245(.a(s_243), .O(gate65inter4));
  nand2 gate2246(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate2247(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate2248(.a(G25), .O(gate65inter7));
  inv1  gate2249(.a(G302), .O(gate65inter8));
  nand2 gate2250(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate2251(.a(s_243), .b(gate65inter3), .O(gate65inter10));
  nor2  gate2252(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate2253(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate2254(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate2353(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate2354(.a(gate70inter0), .b(s_258), .O(gate70inter1));
  and2  gate2355(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate2356(.a(s_258), .O(gate70inter3));
  inv1  gate2357(.a(s_259), .O(gate70inter4));
  nand2 gate2358(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate2359(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate2360(.a(G30), .O(gate70inter7));
  inv1  gate2361(.a(G308), .O(gate70inter8));
  nand2 gate2362(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate2363(.a(s_259), .b(gate70inter3), .O(gate70inter10));
  nor2  gate2364(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate2365(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate2366(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );

  xor2  gate2269(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate2270(.a(gate72inter0), .b(s_246), .O(gate72inter1));
  and2  gate2271(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate2272(.a(s_246), .O(gate72inter3));
  inv1  gate2273(.a(s_247), .O(gate72inter4));
  nand2 gate2274(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate2275(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate2276(.a(G32), .O(gate72inter7));
  inv1  gate2277(.a(G311), .O(gate72inter8));
  nand2 gate2278(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate2279(.a(s_247), .b(gate72inter3), .O(gate72inter10));
  nor2  gate2280(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate2281(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate2282(.a(gate72inter12), .b(gate72inter1), .O(G393));
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate1401(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate1402(.a(gate74inter0), .b(s_122), .O(gate74inter1));
  and2  gate1403(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate1404(.a(s_122), .O(gate74inter3));
  inv1  gate1405(.a(s_123), .O(gate74inter4));
  nand2 gate1406(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate1407(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate1408(.a(G5), .O(gate74inter7));
  inv1  gate1409(.a(G314), .O(gate74inter8));
  nand2 gate1410(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate1411(.a(s_123), .b(gate74inter3), .O(gate74inter10));
  nor2  gate1412(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate1413(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate1414(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate2143(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate2144(.a(gate78inter0), .b(s_228), .O(gate78inter1));
  and2  gate2145(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate2146(.a(s_228), .O(gate78inter3));
  inv1  gate2147(.a(s_229), .O(gate78inter4));
  nand2 gate2148(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate2149(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate2150(.a(G6), .O(gate78inter7));
  inv1  gate2151(.a(G320), .O(gate78inter8));
  nand2 gate2152(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate2153(.a(s_229), .b(gate78inter3), .O(gate78inter10));
  nor2  gate2154(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate2155(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate2156(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate2171(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate2172(.a(gate80inter0), .b(s_232), .O(gate80inter1));
  and2  gate2173(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate2174(.a(s_232), .O(gate80inter3));
  inv1  gate2175(.a(s_233), .O(gate80inter4));
  nand2 gate2176(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate2177(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate2178(.a(G14), .O(gate80inter7));
  inv1  gate2179(.a(G323), .O(gate80inter8));
  nand2 gate2180(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate2181(.a(s_233), .b(gate80inter3), .O(gate80inter10));
  nor2  gate2182(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate2183(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate2184(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );

  xor2  gate1653(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate1654(.a(gate84inter0), .b(s_158), .O(gate84inter1));
  and2  gate1655(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate1656(.a(s_158), .O(gate84inter3));
  inv1  gate1657(.a(s_159), .O(gate84inter4));
  nand2 gate1658(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate1659(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate1660(.a(G15), .O(gate84inter7));
  inv1  gate1661(.a(G329), .O(gate84inter8));
  nand2 gate1662(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate1663(.a(s_159), .b(gate84inter3), .O(gate84inter10));
  nor2  gate1664(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate1665(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate1666(.a(gate84inter12), .b(gate84inter1), .O(G405));
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate1415(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate1416(.a(gate90inter0), .b(s_124), .O(gate90inter1));
  and2  gate1417(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate1418(.a(s_124), .O(gate90inter3));
  inv1  gate1419(.a(s_125), .O(gate90inter4));
  nand2 gate1420(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate1421(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate1422(.a(G21), .O(gate90inter7));
  inv1  gate1423(.a(G338), .O(gate90inter8));
  nand2 gate1424(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate1425(.a(s_125), .b(gate90inter3), .O(gate90inter10));
  nor2  gate1426(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate1427(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate1428(.a(gate90inter12), .b(gate90inter1), .O(G411));
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate2213(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate2214(.a(gate96inter0), .b(s_238), .O(gate96inter1));
  and2  gate2215(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate2216(.a(s_238), .O(gate96inter3));
  inv1  gate2217(.a(s_239), .O(gate96inter4));
  nand2 gate2218(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate2219(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate2220(.a(G30), .O(gate96inter7));
  inv1  gate2221(.a(G347), .O(gate96inter8));
  nand2 gate2222(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate2223(.a(s_239), .b(gate96inter3), .O(gate96inter10));
  nor2  gate2224(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate2225(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate2226(.a(gate96inter12), .b(gate96inter1), .O(G417));
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate2395(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate2396(.a(gate100inter0), .b(s_264), .O(gate100inter1));
  and2  gate2397(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate2398(.a(s_264), .O(gate100inter3));
  inv1  gate2399(.a(s_265), .O(gate100inter4));
  nand2 gate2400(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate2401(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate2402(.a(G31), .O(gate100inter7));
  inv1  gate2403(.a(G353), .O(gate100inter8));
  nand2 gate2404(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate2405(.a(s_265), .b(gate100inter3), .O(gate100inter10));
  nor2  gate2406(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate2407(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate2408(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate2087(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate2088(.a(gate102inter0), .b(s_220), .O(gate102inter1));
  and2  gate2089(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate2090(.a(s_220), .O(gate102inter3));
  inv1  gate2091(.a(s_221), .O(gate102inter4));
  nand2 gate2092(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate2093(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate2094(.a(G24), .O(gate102inter7));
  inv1  gate2095(.a(G356), .O(gate102inter8));
  nand2 gate2096(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate2097(.a(s_221), .b(gate102inter3), .O(gate102inter10));
  nor2  gate2098(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate2099(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate2100(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate1345(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate1346(.a(gate109inter0), .b(s_114), .O(gate109inter1));
  and2  gate1347(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate1348(.a(s_114), .O(gate109inter3));
  inv1  gate1349(.a(s_115), .O(gate109inter4));
  nand2 gate1350(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate1351(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate1352(.a(G370), .O(gate109inter7));
  inv1  gate1353(.a(G371), .O(gate109inter8));
  nand2 gate1354(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate1355(.a(s_115), .b(gate109inter3), .O(gate109inter10));
  nor2  gate1356(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate1357(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate1358(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );

  xor2  gate1765(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate1766(.a(gate113inter0), .b(s_174), .O(gate113inter1));
  and2  gate1767(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate1768(.a(s_174), .O(gate113inter3));
  inv1  gate1769(.a(s_175), .O(gate113inter4));
  nand2 gate1770(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate1771(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate1772(.a(G378), .O(gate113inter7));
  inv1  gate1773(.a(G379), .O(gate113inter8));
  nand2 gate1774(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate1775(.a(s_175), .b(gate113inter3), .O(gate113inter10));
  nor2  gate1776(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate1777(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate1778(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate2199(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate2200(.a(gate115inter0), .b(s_236), .O(gate115inter1));
  and2  gate2201(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate2202(.a(s_236), .O(gate115inter3));
  inv1  gate2203(.a(s_237), .O(gate115inter4));
  nand2 gate2204(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate2205(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate2206(.a(G382), .O(gate115inter7));
  inv1  gate2207(.a(G383), .O(gate115inter8));
  nand2 gate2208(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate2209(.a(s_237), .b(gate115inter3), .O(gate115inter10));
  nor2  gate2210(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate2211(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate2212(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate1835(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate1836(.a(gate119inter0), .b(s_184), .O(gate119inter1));
  and2  gate1837(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate1838(.a(s_184), .O(gate119inter3));
  inv1  gate1839(.a(s_185), .O(gate119inter4));
  nand2 gate1840(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate1841(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate1842(.a(G390), .O(gate119inter7));
  inv1  gate1843(.a(G391), .O(gate119inter8));
  nand2 gate1844(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate1845(.a(s_185), .b(gate119inter3), .O(gate119inter10));
  nor2  gate1846(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate1847(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate1848(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate2409(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate2410(.a(gate124inter0), .b(s_266), .O(gate124inter1));
  and2  gate2411(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate2412(.a(s_266), .O(gate124inter3));
  inv1  gate2413(.a(s_267), .O(gate124inter4));
  nand2 gate2414(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate2415(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate2416(.a(G400), .O(gate124inter7));
  inv1  gate2417(.a(G401), .O(gate124inter8));
  nand2 gate2418(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate2419(.a(s_267), .b(gate124inter3), .O(gate124inter10));
  nor2  gate2420(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate2421(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate2422(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate1849(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate1850(.a(gate126inter0), .b(s_186), .O(gate126inter1));
  and2  gate1851(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate1852(.a(s_186), .O(gate126inter3));
  inv1  gate1853(.a(s_187), .O(gate126inter4));
  nand2 gate1854(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate1855(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate1856(.a(G404), .O(gate126inter7));
  inv1  gate1857(.a(G405), .O(gate126inter8));
  nand2 gate1858(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate1859(.a(s_187), .b(gate126inter3), .O(gate126inter10));
  nor2  gate1860(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate1861(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate1862(.a(gate126inter12), .b(gate126inter1), .O(G489));

  xor2  gate575(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate576(.a(gate127inter0), .b(s_4), .O(gate127inter1));
  and2  gate577(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate578(.a(s_4), .O(gate127inter3));
  inv1  gate579(.a(s_5), .O(gate127inter4));
  nand2 gate580(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate581(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate582(.a(G406), .O(gate127inter7));
  inv1  gate583(.a(G407), .O(gate127inter8));
  nand2 gate584(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate585(.a(s_5), .b(gate127inter3), .O(gate127inter10));
  nor2  gate586(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate587(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate588(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );

  xor2  gate1023(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate1024(.a(gate129inter0), .b(s_68), .O(gate129inter1));
  and2  gate1025(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate1026(.a(s_68), .O(gate129inter3));
  inv1  gate1027(.a(s_69), .O(gate129inter4));
  nand2 gate1028(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate1029(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate1030(.a(G410), .O(gate129inter7));
  inv1  gate1031(.a(G411), .O(gate129inter8));
  nand2 gate1032(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate1033(.a(s_69), .b(gate129inter3), .O(gate129inter10));
  nor2  gate1034(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate1035(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate1036(.a(gate129inter12), .b(gate129inter1), .O(G498));
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate981(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate982(.a(gate131inter0), .b(s_62), .O(gate131inter1));
  and2  gate983(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate984(.a(s_62), .O(gate131inter3));
  inv1  gate985(.a(s_63), .O(gate131inter4));
  nand2 gate986(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate987(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate988(.a(G414), .O(gate131inter7));
  inv1  gate989(.a(G415), .O(gate131inter8));
  nand2 gate990(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate991(.a(s_63), .b(gate131inter3), .O(gate131inter10));
  nor2  gate992(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate993(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate994(.a(gate131inter12), .b(gate131inter1), .O(G504));

  xor2  gate841(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate842(.a(gate132inter0), .b(s_42), .O(gate132inter1));
  and2  gate843(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate844(.a(s_42), .O(gate132inter3));
  inv1  gate845(.a(s_43), .O(gate132inter4));
  nand2 gate846(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate847(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate848(.a(G416), .O(gate132inter7));
  inv1  gate849(.a(G417), .O(gate132inter8));
  nand2 gate850(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate851(.a(s_43), .b(gate132inter3), .O(gate132inter10));
  nor2  gate852(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate853(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate854(.a(gate132inter12), .b(gate132inter1), .O(G507));

  xor2  gate1317(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate1318(.a(gate133inter0), .b(s_110), .O(gate133inter1));
  and2  gate1319(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate1320(.a(s_110), .O(gate133inter3));
  inv1  gate1321(.a(s_111), .O(gate133inter4));
  nand2 gate1322(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate1323(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate1324(.a(G418), .O(gate133inter7));
  inv1  gate1325(.a(G419), .O(gate133inter8));
  nand2 gate1326(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate1327(.a(s_111), .b(gate133inter3), .O(gate133inter10));
  nor2  gate1328(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate1329(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate1330(.a(gate133inter12), .b(gate133inter1), .O(G510));
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate995(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate996(.a(gate137inter0), .b(s_64), .O(gate137inter1));
  and2  gate997(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate998(.a(s_64), .O(gate137inter3));
  inv1  gate999(.a(s_65), .O(gate137inter4));
  nand2 gate1000(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate1001(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate1002(.a(G426), .O(gate137inter7));
  inv1  gate1003(.a(G429), .O(gate137inter8));
  nand2 gate1004(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate1005(.a(s_65), .b(gate137inter3), .O(gate137inter10));
  nor2  gate1006(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate1007(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate1008(.a(gate137inter12), .b(gate137inter1), .O(G522));

  xor2  gate1205(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate1206(.a(gate138inter0), .b(s_94), .O(gate138inter1));
  and2  gate1207(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate1208(.a(s_94), .O(gate138inter3));
  inv1  gate1209(.a(s_95), .O(gate138inter4));
  nand2 gate1210(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate1211(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate1212(.a(G432), .O(gate138inter7));
  inv1  gate1213(.a(G435), .O(gate138inter8));
  nand2 gate1214(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate1215(.a(s_95), .b(gate138inter3), .O(gate138inter10));
  nor2  gate1216(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate1217(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate1218(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );

  xor2  gate1975(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate1976(.a(gate140inter0), .b(s_204), .O(gate140inter1));
  and2  gate1977(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate1978(.a(s_204), .O(gate140inter3));
  inv1  gate1979(.a(s_205), .O(gate140inter4));
  nand2 gate1980(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate1981(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate1982(.a(G444), .O(gate140inter7));
  inv1  gate1983(.a(G447), .O(gate140inter8));
  nand2 gate1984(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate1985(.a(s_205), .b(gate140inter3), .O(gate140inter10));
  nor2  gate1986(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate1987(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate1988(.a(gate140inter12), .b(gate140inter1), .O(G531));
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate2129(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate2130(.a(gate143inter0), .b(s_226), .O(gate143inter1));
  and2  gate2131(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate2132(.a(s_226), .O(gate143inter3));
  inv1  gate2133(.a(s_227), .O(gate143inter4));
  nand2 gate2134(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate2135(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate2136(.a(G462), .O(gate143inter7));
  inv1  gate2137(.a(G465), .O(gate143inter8));
  nand2 gate2138(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate2139(.a(s_227), .b(gate143inter3), .O(gate143inter10));
  nor2  gate2140(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate2141(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate2142(.a(gate143inter12), .b(gate143inter1), .O(G540));

  xor2  gate1009(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate1010(.a(gate144inter0), .b(s_66), .O(gate144inter1));
  and2  gate1011(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate1012(.a(s_66), .O(gate144inter3));
  inv1  gate1013(.a(s_67), .O(gate144inter4));
  nand2 gate1014(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate1015(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate1016(.a(G468), .O(gate144inter7));
  inv1  gate1017(.a(G471), .O(gate144inter8));
  nand2 gate1018(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate1019(.a(s_67), .b(gate144inter3), .O(gate144inter10));
  nor2  gate1020(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate1021(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate1022(.a(gate144inter12), .b(gate144inter1), .O(G543));

  xor2  gate1779(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate1780(.a(gate145inter0), .b(s_176), .O(gate145inter1));
  and2  gate1781(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate1782(.a(s_176), .O(gate145inter3));
  inv1  gate1783(.a(s_177), .O(gate145inter4));
  nand2 gate1784(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate1785(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate1786(.a(G474), .O(gate145inter7));
  inv1  gate1787(.a(G477), .O(gate145inter8));
  nand2 gate1788(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate1789(.a(s_177), .b(gate145inter3), .O(gate145inter10));
  nor2  gate1790(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate1791(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate1792(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate1807(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate1808(.a(gate149inter0), .b(s_180), .O(gate149inter1));
  and2  gate1809(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate1810(.a(s_180), .O(gate149inter3));
  inv1  gate1811(.a(s_181), .O(gate149inter4));
  nand2 gate1812(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate1813(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate1814(.a(G498), .O(gate149inter7));
  inv1  gate1815(.a(G501), .O(gate149inter8));
  nand2 gate1816(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate1817(.a(s_181), .b(gate149inter3), .O(gate149inter10));
  nor2  gate1818(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate1819(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate1820(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );

  xor2  gate2073(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate2074(.a(gate152inter0), .b(s_218), .O(gate152inter1));
  and2  gate2075(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate2076(.a(s_218), .O(gate152inter3));
  inv1  gate2077(.a(s_219), .O(gate152inter4));
  nand2 gate2078(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate2079(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate2080(.a(G516), .O(gate152inter7));
  inv1  gate2081(.a(G519), .O(gate152inter8));
  nand2 gate2082(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate2083(.a(s_219), .b(gate152inter3), .O(gate152inter10));
  nor2  gate2084(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate2085(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate2086(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate1905(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate1906(.a(gate154inter0), .b(s_194), .O(gate154inter1));
  and2  gate1907(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate1908(.a(s_194), .O(gate154inter3));
  inv1  gate1909(.a(s_195), .O(gate154inter4));
  nand2 gate1910(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate1911(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate1912(.a(G429), .O(gate154inter7));
  inv1  gate1913(.a(G522), .O(gate154inter8));
  nand2 gate1914(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate1915(.a(s_195), .b(gate154inter3), .O(gate154inter10));
  nor2  gate1916(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate1917(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate1918(.a(gate154inter12), .b(gate154inter1), .O(G571));

  xor2  gate2367(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate2368(.a(gate155inter0), .b(s_260), .O(gate155inter1));
  and2  gate2369(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate2370(.a(s_260), .O(gate155inter3));
  inv1  gate2371(.a(s_261), .O(gate155inter4));
  nand2 gate2372(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate2373(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate2374(.a(G432), .O(gate155inter7));
  inv1  gate2375(.a(G525), .O(gate155inter8));
  nand2 gate2376(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate2377(.a(s_261), .b(gate155inter3), .O(gate155inter10));
  nor2  gate2378(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate2379(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate2380(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate1667(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate1668(.a(gate159inter0), .b(s_160), .O(gate159inter1));
  and2  gate1669(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate1670(.a(s_160), .O(gate159inter3));
  inv1  gate1671(.a(s_161), .O(gate159inter4));
  nand2 gate1672(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate1673(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate1674(.a(G444), .O(gate159inter7));
  inv1  gate1675(.a(G531), .O(gate159inter8));
  nand2 gate1676(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate1677(.a(s_161), .b(gate159inter3), .O(gate159inter10));
  nor2  gate1678(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate1679(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate1680(.a(gate159inter12), .b(gate159inter1), .O(G576));

  xor2  gate1107(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate1108(.a(gate160inter0), .b(s_80), .O(gate160inter1));
  and2  gate1109(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate1110(.a(s_80), .O(gate160inter3));
  inv1  gate1111(.a(s_81), .O(gate160inter4));
  nand2 gate1112(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate1113(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate1114(.a(G447), .O(gate160inter7));
  inv1  gate1115(.a(G531), .O(gate160inter8));
  nand2 gate1116(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate1117(.a(s_81), .b(gate160inter3), .O(gate160inter10));
  nor2  gate1118(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate1119(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate1120(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate2339(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate2340(.a(gate162inter0), .b(s_256), .O(gate162inter1));
  and2  gate2341(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate2342(.a(s_256), .O(gate162inter3));
  inv1  gate2343(.a(s_257), .O(gate162inter4));
  nand2 gate2344(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate2345(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate2346(.a(G453), .O(gate162inter7));
  inv1  gate2347(.a(G534), .O(gate162inter8));
  nand2 gate2348(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate2349(.a(s_257), .b(gate162inter3), .O(gate162inter10));
  nor2  gate2350(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate2351(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate2352(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );

  xor2  gate1681(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate1682(.a(gate166inter0), .b(s_162), .O(gate166inter1));
  and2  gate1683(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate1684(.a(s_162), .O(gate166inter3));
  inv1  gate1685(.a(s_163), .O(gate166inter4));
  nand2 gate1686(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate1687(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate1688(.a(G465), .O(gate166inter7));
  inv1  gate1689(.a(G540), .O(gate166inter8));
  nand2 gate1690(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate1691(.a(s_163), .b(gate166inter3), .O(gate166inter10));
  nor2  gate1692(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate1693(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate1694(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );

  xor2  gate1751(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate1752(.a(gate169inter0), .b(s_172), .O(gate169inter1));
  and2  gate1753(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate1754(.a(s_172), .O(gate169inter3));
  inv1  gate1755(.a(s_173), .O(gate169inter4));
  nand2 gate1756(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate1757(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate1758(.a(G474), .O(gate169inter7));
  inv1  gate1759(.a(G546), .O(gate169inter8));
  nand2 gate1760(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate1761(.a(s_173), .b(gate169inter3), .O(gate169inter10));
  nor2  gate1762(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate1763(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate1764(.a(gate169inter12), .b(gate169inter1), .O(G586));
nand2 gate170( .a(G477), .b(G546), .O(G587) );

  xor2  gate883(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate884(.a(gate171inter0), .b(s_48), .O(gate171inter1));
  and2  gate885(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate886(.a(s_48), .O(gate171inter3));
  inv1  gate887(.a(s_49), .O(gate171inter4));
  nand2 gate888(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate889(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate890(.a(G480), .O(gate171inter7));
  inv1  gate891(.a(G549), .O(gate171inter8));
  nand2 gate892(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate893(.a(s_49), .b(gate171inter3), .O(gate171inter10));
  nor2  gate894(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate895(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate896(.a(gate171inter12), .b(gate171inter1), .O(G588));
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate1331(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate1332(.a(gate178inter0), .b(s_112), .O(gate178inter1));
  and2  gate1333(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate1334(.a(s_112), .O(gate178inter3));
  inv1  gate1335(.a(s_113), .O(gate178inter4));
  nand2 gate1336(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate1337(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate1338(.a(G501), .O(gate178inter7));
  inv1  gate1339(.a(G558), .O(gate178inter8));
  nand2 gate1340(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate1341(.a(s_113), .b(gate178inter3), .O(gate178inter10));
  nor2  gate1342(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate1343(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate1344(.a(gate178inter12), .b(gate178inter1), .O(G595));
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate2115(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate2116(.a(gate180inter0), .b(s_224), .O(gate180inter1));
  and2  gate2117(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate2118(.a(s_224), .O(gate180inter3));
  inv1  gate2119(.a(s_225), .O(gate180inter4));
  nand2 gate2120(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate2121(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate2122(.a(G507), .O(gate180inter7));
  inv1  gate2123(.a(G561), .O(gate180inter8));
  nand2 gate2124(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate2125(.a(s_225), .b(gate180inter3), .O(gate180inter10));
  nor2  gate2126(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate2127(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate2128(.a(gate180inter12), .b(gate180inter1), .O(G597));
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate589(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate590(.a(gate183inter0), .b(s_6), .O(gate183inter1));
  and2  gate591(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate592(.a(s_6), .O(gate183inter3));
  inv1  gate593(.a(s_7), .O(gate183inter4));
  nand2 gate594(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate595(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate596(.a(G516), .O(gate183inter7));
  inv1  gate597(.a(G567), .O(gate183inter8));
  nand2 gate598(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate599(.a(s_7), .b(gate183inter3), .O(gate183inter10));
  nor2  gate600(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate601(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate602(.a(gate183inter12), .b(gate183inter1), .O(G600));

  xor2  gate1387(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate1388(.a(gate184inter0), .b(s_120), .O(gate184inter1));
  and2  gate1389(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate1390(.a(s_120), .O(gate184inter3));
  inv1  gate1391(.a(s_121), .O(gate184inter4));
  nand2 gate1392(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate1393(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate1394(.a(G519), .O(gate184inter7));
  inv1  gate1395(.a(G567), .O(gate184inter8));
  nand2 gate1396(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate1397(.a(s_121), .b(gate184inter3), .O(gate184inter10));
  nor2  gate1398(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate1399(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate1400(.a(gate184inter12), .b(gate184inter1), .O(G601));

  xor2  gate1793(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate1794(.a(gate185inter0), .b(s_178), .O(gate185inter1));
  and2  gate1795(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate1796(.a(s_178), .O(gate185inter3));
  inv1  gate1797(.a(s_179), .O(gate185inter4));
  nand2 gate1798(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate1799(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate1800(.a(G570), .O(gate185inter7));
  inv1  gate1801(.a(G571), .O(gate185inter8));
  nand2 gate1802(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate1803(.a(s_179), .b(gate185inter3), .O(gate185inter10));
  nor2  gate1804(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate1805(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate1806(.a(gate185inter12), .b(gate185inter1), .O(G602));
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate1177(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate1178(.a(gate193inter0), .b(s_90), .O(gate193inter1));
  and2  gate1179(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate1180(.a(s_90), .O(gate193inter3));
  inv1  gate1181(.a(s_91), .O(gate193inter4));
  nand2 gate1182(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate1183(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate1184(.a(G586), .O(gate193inter7));
  inv1  gate1185(.a(G587), .O(gate193inter8));
  nand2 gate1186(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate1187(.a(s_91), .b(gate193inter3), .O(gate193inter10));
  nor2  gate1188(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate1189(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate1190(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate953(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate954(.a(gate201inter0), .b(s_58), .O(gate201inter1));
  and2  gate955(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate956(.a(s_58), .O(gate201inter3));
  inv1  gate957(.a(s_59), .O(gate201inter4));
  nand2 gate958(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate959(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate960(.a(G602), .O(gate201inter7));
  inv1  gate961(.a(G607), .O(gate201inter8));
  nand2 gate962(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate963(.a(s_59), .b(gate201inter3), .O(gate201inter10));
  nor2  gate964(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate965(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate966(.a(gate201inter12), .b(gate201inter1), .O(G666));

  xor2  gate1527(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate1528(.a(gate202inter0), .b(s_140), .O(gate202inter1));
  and2  gate1529(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate1530(.a(s_140), .O(gate202inter3));
  inv1  gate1531(.a(s_141), .O(gate202inter4));
  nand2 gate1532(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate1533(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate1534(.a(G612), .O(gate202inter7));
  inv1  gate1535(.a(G617), .O(gate202inter8));
  nand2 gate1536(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate1537(.a(s_141), .b(gate202inter3), .O(gate202inter10));
  nor2  gate1538(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate1539(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate1540(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );

  xor2  gate2437(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate2438(.a(gate208inter0), .b(s_270), .O(gate208inter1));
  and2  gate2439(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate2440(.a(s_270), .O(gate208inter3));
  inv1  gate2441(.a(s_271), .O(gate208inter4));
  nand2 gate2442(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate2443(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate2444(.a(G627), .O(gate208inter7));
  inv1  gate2445(.a(G637), .O(gate208inter8));
  nand2 gate2446(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate2447(.a(s_271), .b(gate208inter3), .O(gate208inter10));
  nor2  gate2448(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate2449(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate2450(.a(gate208inter12), .b(gate208inter1), .O(G687));
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate757(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate758(.a(gate213inter0), .b(s_30), .O(gate213inter1));
  and2  gate759(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate760(.a(s_30), .O(gate213inter3));
  inv1  gate761(.a(s_31), .O(gate213inter4));
  nand2 gate762(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate763(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate764(.a(G602), .O(gate213inter7));
  inv1  gate765(.a(G672), .O(gate213inter8));
  nand2 gate766(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate767(.a(s_31), .b(gate213inter3), .O(gate213inter10));
  nor2  gate768(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate769(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate770(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate1219(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate1220(.a(gate215inter0), .b(s_96), .O(gate215inter1));
  and2  gate1221(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate1222(.a(s_96), .O(gate215inter3));
  inv1  gate1223(.a(s_97), .O(gate215inter4));
  nand2 gate1224(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate1225(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate1226(.a(G607), .O(gate215inter7));
  inv1  gate1227(.a(G675), .O(gate215inter8));
  nand2 gate1228(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate1229(.a(s_97), .b(gate215inter3), .O(gate215inter10));
  nor2  gate1230(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate1231(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate1232(.a(gate215inter12), .b(gate215inter1), .O(G696));

  xor2  gate1723(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate1724(.a(gate216inter0), .b(s_168), .O(gate216inter1));
  and2  gate1725(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate1726(.a(s_168), .O(gate216inter3));
  inv1  gate1727(.a(s_169), .O(gate216inter4));
  nand2 gate1728(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate1729(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate1730(.a(G617), .O(gate216inter7));
  inv1  gate1731(.a(G675), .O(gate216inter8));
  nand2 gate1732(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate1733(.a(s_169), .b(gate216inter3), .O(gate216inter10));
  nor2  gate1734(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate1735(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate1736(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate2059(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate2060(.a(gate220inter0), .b(s_216), .O(gate220inter1));
  and2  gate2061(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate2062(.a(s_216), .O(gate220inter3));
  inv1  gate2063(.a(s_217), .O(gate220inter4));
  nand2 gate2064(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate2065(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate2066(.a(G637), .O(gate220inter7));
  inv1  gate2067(.a(G681), .O(gate220inter8));
  nand2 gate2068(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate2069(.a(s_217), .b(gate220inter3), .O(gate220inter10));
  nor2  gate2070(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate2071(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate2072(.a(gate220inter12), .b(gate220inter1), .O(G701));

  xor2  gate617(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate618(.a(gate221inter0), .b(s_10), .O(gate221inter1));
  and2  gate619(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate620(.a(s_10), .O(gate221inter3));
  inv1  gate621(.a(s_11), .O(gate221inter4));
  nand2 gate622(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate623(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate624(.a(G622), .O(gate221inter7));
  inv1  gate625(.a(G684), .O(gate221inter8));
  nand2 gate626(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate627(.a(s_11), .b(gate221inter3), .O(gate221inter10));
  nor2  gate628(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate629(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate630(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate1065(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate1066(.a(gate223inter0), .b(s_74), .O(gate223inter1));
  and2  gate1067(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate1068(.a(s_74), .O(gate223inter3));
  inv1  gate1069(.a(s_75), .O(gate223inter4));
  nand2 gate1070(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate1071(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate1072(.a(G627), .O(gate223inter7));
  inv1  gate1073(.a(G687), .O(gate223inter8));
  nand2 gate1074(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate1075(.a(s_75), .b(gate223inter3), .O(gate223inter10));
  nor2  gate1076(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate1077(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate1078(.a(gate223inter12), .b(gate223inter1), .O(G704));

  xor2  gate1919(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate1920(.a(gate224inter0), .b(s_196), .O(gate224inter1));
  and2  gate1921(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate1922(.a(s_196), .O(gate224inter3));
  inv1  gate1923(.a(s_197), .O(gate224inter4));
  nand2 gate1924(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate1925(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate1926(.a(G637), .O(gate224inter7));
  inv1  gate1927(.a(G687), .O(gate224inter8));
  nand2 gate1928(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate1929(.a(s_197), .b(gate224inter3), .O(gate224inter10));
  nor2  gate1930(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate1931(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate1932(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate1737(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate1738(.a(gate227inter0), .b(s_170), .O(gate227inter1));
  and2  gate1739(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate1740(.a(s_170), .O(gate227inter3));
  inv1  gate1741(.a(s_171), .O(gate227inter4));
  nand2 gate1742(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate1743(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate1744(.a(G694), .O(gate227inter7));
  inv1  gate1745(.a(G695), .O(gate227inter8));
  nand2 gate1746(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate1747(.a(s_171), .b(gate227inter3), .O(gate227inter10));
  nor2  gate1748(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate1749(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate1750(.a(gate227inter12), .b(gate227inter1), .O(G712));
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );

  xor2  gate1191(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate1192(.a(gate238inter0), .b(s_92), .O(gate238inter1));
  and2  gate1193(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate1194(.a(s_92), .O(gate238inter3));
  inv1  gate1195(.a(s_93), .O(gate238inter4));
  nand2 gate1196(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate1197(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate1198(.a(G257), .O(gate238inter7));
  inv1  gate1199(.a(G709), .O(gate238inter8));
  nand2 gate1200(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate1201(.a(s_93), .b(gate238inter3), .O(gate238inter10));
  nor2  gate1202(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate1203(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate1204(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate771(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate772(.a(gate240inter0), .b(s_32), .O(gate240inter1));
  and2  gate773(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate774(.a(s_32), .O(gate240inter3));
  inv1  gate775(.a(s_33), .O(gate240inter4));
  nand2 gate776(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate777(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate778(.a(G263), .O(gate240inter7));
  inv1  gate779(.a(G715), .O(gate240inter8));
  nand2 gate780(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate781(.a(s_33), .b(gate240inter3), .O(gate240inter10));
  nor2  gate782(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate783(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate784(.a(gate240inter12), .b(gate240inter1), .O(G751));

  xor2  gate631(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate632(.a(gate241inter0), .b(s_12), .O(gate241inter1));
  and2  gate633(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate634(.a(s_12), .O(gate241inter3));
  inv1  gate635(.a(s_13), .O(gate241inter4));
  nand2 gate636(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate637(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate638(.a(G242), .O(gate241inter7));
  inv1  gate639(.a(G730), .O(gate241inter8));
  nand2 gate640(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate641(.a(s_13), .b(gate241inter3), .O(gate241inter10));
  nor2  gate642(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate643(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate644(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );

  xor2  gate2157(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate2158(.a(gate246inter0), .b(s_230), .O(gate246inter1));
  and2  gate2159(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate2160(.a(s_230), .O(gate246inter3));
  inv1  gate2161(.a(s_231), .O(gate246inter4));
  nand2 gate2162(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate2163(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate2164(.a(G724), .O(gate246inter7));
  inv1  gate2165(.a(G736), .O(gate246inter8));
  nand2 gate2166(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate2167(.a(s_231), .b(gate246inter3), .O(gate246inter10));
  nor2  gate2168(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate2169(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate2170(.a(gate246inter12), .b(gate246inter1), .O(G759));

  xor2  gate1933(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate1934(.a(gate247inter0), .b(s_198), .O(gate247inter1));
  and2  gate1935(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate1936(.a(s_198), .O(gate247inter3));
  inv1  gate1937(.a(s_199), .O(gate247inter4));
  nand2 gate1938(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate1939(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate1940(.a(G251), .O(gate247inter7));
  inv1  gate1941(.a(G739), .O(gate247inter8));
  nand2 gate1942(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate1943(.a(s_199), .b(gate247inter3), .O(gate247inter10));
  nor2  gate1944(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate1945(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate1946(.a(gate247inter12), .b(gate247inter1), .O(G760));
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );

  xor2  gate2297(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate2298(.a(gate254inter0), .b(s_250), .O(gate254inter1));
  and2  gate2299(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate2300(.a(s_250), .O(gate254inter3));
  inv1  gate2301(.a(s_251), .O(gate254inter4));
  nand2 gate2302(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate2303(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate2304(.a(G712), .O(gate254inter7));
  inv1  gate2305(.a(G748), .O(gate254inter8));
  nand2 gate2306(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate2307(.a(s_251), .b(gate254inter3), .O(gate254inter10));
  nor2  gate2308(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate2309(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate2310(.a(gate254inter12), .b(gate254inter1), .O(G767));
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate1513(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate1514(.a(gate256inter0), .b(s_138), .O(gate256inter1));
  and2  gate1515(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate1516(.a(s_138), .O(gate256inter3));
  inv1  gate1517(.a(s_139), .O(gate256inter4));
  nand2 gate1518(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate1519(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate1520(.a(G715), .O(gate256inter7));
  inv1  gate1521(.a(G751), .O(gate256inter8));
  nand2 gate1522(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate1523(.a(s_139), .b(gate256inter3), .O(gate256inter10));
  nor2  gate1524(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate1525(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate1526(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );

  xor2  gate1611(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate1612(.a(gate259inter0), .b(s_152), .O(gate259inter1));
  and2  gate1613(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate1614(.a(s_152), .O(gate259inter3));
  inv1  gate1615(.a(s_153), .O(gate259inter4));
  nand2 gate1616(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate1617(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate1618(.a(G758), .O(gate259inter7));
  inv1  gate1619(.a(G759), .O(gate259inter8));
  nand2 gate1620(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate1621(.a(s_153), .b(gate259inter3), .O(gate259inter10));
  nor2  gate1622(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate1623(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate1624(.a(gate259inter12), .b(gate259inter1), .O(G776));
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate1891(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate1892(.a(gate261inter0), .b(s_192), .O(gate261inter1));
  and2  gate1893(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate1894(.a(s_192), .O(gate261inter3));
  inv1  gate1895(.a(s_193), .O(gate261inter4));
  nand2 gate1896(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate1897(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate1898(.a(G762), .O(gate261inter7));
  inv1  gate1899(.a(G763), .O(gate261inter8));
  nand2 gate1900(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate1901(.a(s_193), .b(gate261inter3), .O(gate261inter10));
  nor2  gate1902(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate1903(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate1904(.a(gate261inter12), .b(gate261inter1), .O(G782));

  xor2  gate1275(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate1276(.a(gate262inter0), .b(s_104), .O(gate262inter1));
  and2  gate1277(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate1278(.a(s_104), .O(gate262inter3));
  inv1  gate1279(.a(s_105), .O(gate262inter4));
  nand2 gate1280(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate1281(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate1282(.a(G764), .O(gate262inter7));
  inv1  gate1283(.a(G765), .O(gate262inter8));
  nand2 gate1284(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate1285(.a(s_105), .b(gate262inter3), .O(gate262inter10));
  nor2  gate1286(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate1287(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate1288(.a(gate262inter12), .b(gate262inter1), .O(G785));

  xor2  gate1303(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate1304(.a(gate263inter0), .b(s_108), .O(gate263inter1));
  and2  gate1305(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate1306(.a(s_108), .O(gate263inter3));
  inv1  gate1307(.a(s_109), .O(gate263inter4));
  nand2 gate1308(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate1309(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate1310(.a(G766), .O(gate263inter7));
  inv1  gate1311(.a(G767), .O(gate263inter8));
  nand2 gate1312(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate1313(.a(s_109), .b(gate263inter3), .O(gate263inter10));
  nor2  gate1314(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate1315(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate1316(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate1863(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate1864(.a(gate265inter0), .b(s_188), .O(gate265inter1));
  and2  gate1865(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate1866(.a(s_188), .O(gate265inter3));
  inv1  gate1867(.a(s_189), .O(gate265inter4));
  nand2 gate1868(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate1869(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate1870(.a(G642), .O(gate265inter7));
  inv1  gate1871(.a(G770), .O(gate265inter8));
  nand2 gate1872(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate1873(.a(s_189), .b(gate265inter3), .O(gate265inter10));
  nor2  gate1874(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate1875(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate1876(.a(gate265inter12), .b(gate265inter1), .O(G794));
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate2017(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate2018(.a(gate269inter0), .b(s_210), .O(gate269inter1));
  and2  gate2019(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate2020(.a(s_210), .O(gate269inter3));
  inv1  gate2021(.a(s_211), .O(gate269inter4));
  nand2 gate2022(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate2023(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate2024(.a(G654), .O(gate269inter7));
  inv1  gate2025(.a(G782), .O(gate269inter8));
  nand2 gate2026(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate2027(.a(s_211), .b(gate269inter3), .O(gate269inter10));
  nor2  gate2028(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate2029(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate2030(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );

  xor2  gate2101(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate2102(.a(gate275inter0), .b(s_222), .O(gate275inter1));
  and2  gate2103(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate2104(.a(s_222), .O(gate275inter3));
  inv1  gate2105(.a(s_223), .O(gate275inter4));
  nand2 gate2106(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate2107(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate2108(.a(G645), .O(gate275inter7));
  inv1  gate2109(.a(G797), .O(gate275inter8));
  nand2 gate2110(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate2111(.a(s_223), .b(gate275inter3), .O(gate275inter10));
  nor2  gate2112(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate2113(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate2114(.a(gate275inter12), .b(gate275inter1), .O(G820));

  xor2  gate673(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate674(.a(gate276inter0), .b(s_18), .O(gate276inter1));
  and2  gate675(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate676(.a(s_18), .O(gate276inter3));
  inv1  gate677(.a(s_19), .O(gate276inter4));
  nand2 gate678(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate679(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate680(.a(G773), .O(gate276inter7));
  inv1  gate681(.a(G797), .O(gate276inter8));
  nand2 gate682(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate683(.a(s_19), .b(gate276inter3), .O(gate276inter10));
  nor2  gate684(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate685(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate686(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate1037(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate1038(.a(gate278inter0), .b(s_70), .O(gate278inter1));
  and2  gate1039(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate1040(.a(s_70), .O(gate278inter3));
  inv1  gate1041(.a(s_71), .O(gate278inter4));
  nand2 gate1042(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate1043(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate1044(.a(G776), .O(gate278inter7));
  inv1  gate1045(.a(G800), .O(gate278inter8));
  nand2 gate1046(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate1047(.a(s_71), .b(gate278inter3), .O(gate278inter10));
  nor2  gate1048(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate1049(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate1050(.a(gate278inter12), .b(gate278inter1), .O(G823));

  xor2  gate1625(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate1626(.a(gate279inter0), .b(s_154), .O(gate279inter1));
  and2  gate1627(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate1628(.a(s_154), .O(gate279inter3));
  inv1  gate1629(.a(s_155), .O(gate279inter4));
  nand2 gate1630(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate1631(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate1632(.a(G651), .O(gate279inter7));
  inv1  gate1633(.a(G803), .O(gate279inter8));
  nand2 gate1634(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate1635(.a(s_155), .b(gate279inter3), .O(gate279inter10));
  nor2  gate1636(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate1637(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate1638(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate1261(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate1262(.a(gate283inter0), .b(s_102), .O(gate283inter1));
  and2  gate1263(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate1264(.a(s_102), .O(gate283inter3));
  inv1  gate1265(.a(s_103), .O(gate283inter4));
  nand2 gate1266(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate1267(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate1268(.a(G657), .O(gate283inter7));
  inv1  gate1269(.a(G809), .O(gate283inter8));
  nand2 gate1270(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate1271(.a(s_103), .b(gate283inter3), .O(gate283inter10));
  nor2  gate1272(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate1273(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate1274(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate1989(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate1990(.a(gate286inter0), .b(s_206), .O(gate286inter1));
  and2  gate1991(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate1992(.a(s_206), .O(gate286inter3));
  inv1  gate1993(.a(s_207), .O(gate286inter4));
  nand2 gate1994(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate1995(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate1996(.a(G788), .O(gate286inter7));
  inv1  gate1997(.a(G812), .O(gate286inter8));
  nand2 gate1998(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate1999(.a(s_207), .b(gate286inter3), .O(gate286inter10));
  nor2  gate2000(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate2001(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate2002(.a(gate286inter12), .b(gate286inter1), .O(G831));
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate1541(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate1542(.a(gate292inter0), .b(s_142), .O(gate292inter1));
  and2  gate1543(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate1544(.a(s_142), .O(gate292inter3));
  inv1  gate1545(.a(s_143), .O(gate292inter4));
  nand2 gate1546(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate1547(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate1548(.a(G824), .O(gate292inter7));
  inv1  gate1549(.a(G825), .O(gate292inter8));
  nand2 gate1550(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate1551(.a(s_143), .b(gate292inter3), .O(gate292inter10));
  nor2  gate1552(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate1553(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate1554(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate799(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate800(.a(gate295inter0), .b(s_36), .O(gate295inter1));
  and2  gate801(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate802(.a(s_36), .O(gate295inter3));
  inv1  gate803(.a(s_37), .O(gate295inter4));
  nand2 gate804(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate805(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate806(.a(G830), .O(gate295inter7));
  inv1  gate807(.a(G831), .O(gate295inter8));
  nand2 gate808(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate809(.a(s_37), .b(gate295inter3), .O(gate295inter10));
  nor2  gate810(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate811(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate812(.a(gate295inter12), .b(gate295inter1), .O(G912));

  xor2  gate659(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate660(.a(gate296inter0), .b(s_16), .O(gate296inter1));
  and2  gate661(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate662(.a(s_16), .O(gate296inter3));
  inv1  gate663(.a(s_17), .O(gate296inter4));
  nand2 gate664(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate665(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate666(.a(G826), .O(gate296inter7));
  inv1  gate667(.a(G827), .O(gate296inter8));
  nand2 gate668(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate669(.a(s_17), .b(gate296inter3), .O(gate296inter10));
  nor2  gate670(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate671(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate672(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate1947(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate1948(.a(gate387inter0), .b(s_200), .O(gate387inter1));
  and2  gate1949(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate1950(.a(s_200), .O(gate387inter3));
  inv1  gate1951(.a(s_201), .O(gate387inter4));
  nand2 gate1952(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1953(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1954(.a(G1), .O(gate387inter7));
  inv1  gate1955(.a(G1036), .O(gate387inter8));
  nand2 gate1956(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1957(.a(s_201), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1958(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1959(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate1960(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate1051(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate1052(.a(gate389inter0), .b(s_72), .O(gate389inter1));
  and2  gate1053(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate1054(.a(s_72), .O(gate389inter3));
  inv1  gate1055(.a(s_73), .O(gate389inter4));
  nand2 gate1056(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate1057(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate1058(.a(G3), .O(gate389inter7));
  inv1  gate1059(.a(G1042), .O(gate389inter8));
  nand2 gate1060(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate1061(.a(s_73), .b(gate389inter3), .O(gate389inter10));
  nor2  gate1062(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate1063(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate1064(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate1555(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate1556(.a(gate391inter0), .b(s_144), .O(gate391inter1));
  and2  gate1557(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate1558(.a(s_144), .O(gate391inter3));
  inv1  gate1559(.a(s_145), .O(gate391inter4));
  nand2 gate1560(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate1561(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate1562(.a(G5), .O(gate391inter7));
  inv1  gate1563(.a(G1048), .O(gate391inter8));
  nand2 gate1564(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate1565(.a(s_145), .b(gate391inter3), .O(gate391inter10));
  nor2  gate1566(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate1567(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate1568(.a(gate391inter12), .b(gate391inter1), .O(G1144));

  xor2  gate1429(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate1430(.a(gate392inter0), .b(s_126), .O(gate392inter1));
  and2  gate1431(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate1432(.a(s_126), .O(gate392inter3));
  inv1  gate1433(.a(s_127), .O(gate392inter4));
  nand2 gate1434(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate1435(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate1436(.a(G6), .O(gate392inter7));
  inv1  gate1437(.a(G1051), .O(gate392inter8));
  nand2 gate1438(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate1439(.a(s_127), .b(gate392inter3), .O(gate392inter10));
  nor2  gate1440(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate1441(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate1442(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate897(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate898(.a(gate394inter0), .b(s_50), .O(gate394inter1));
  and2  gate899(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate900(.a(s_50), .O(gate394inter3));
  inv1  gate901(.a(s_51), .O(gate394inter4));
  nand2 gate902(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate903(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate904(.a(G8), .O(gate394inter7));
  inv1  gate905(.a(G1057), .O(gate394inter8));
  nand2 gate906(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate907(.a(s_51), .b(gate394inter3), .O(gate394inter10));
  nor2  gate908(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate909(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate910(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );

  xor2  gate1289(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate1290(.a(gate401inter0), .b(s_106), .O(gate401inter1));
  and2  gate1291(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate1292(.a(s_106), .O(gate401inter3));
  inv1  gate1293(.a(s_107), .O(gate401inter4));
  nand2 gate1294(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate1295(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate1296(.a(G15), .O(gate401inter7));
  inv1  gate1297(.a(G1078), .O(gate401inter8));
  nand2 gate1298(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate1299(.a(s_107), .b(gate401inter3), .O(gate401inter10));
  nor2  gate1300(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate1301(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate1302(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate715(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate716(.a(gate403inter0), .b(s_24), .O(gate403inter1));
  and2  gate717(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate718(.a(s_24), .O(gate403inter3));
  inv1  gate719(.a(s_25), .O(gate403inter4));
  nand2 gate720(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate721(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate722(.a(G17), .O(gate403inter7));
  inv1  gate723(.a(G1084), .O(gate403inter8));
  nand2 gate724(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate725(.a(s_25), .b(gate403inter3), .O(gate403inter10));
  nor2  gate726(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate727(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate728(.a(gate403inter12), .b(gate403inter1), .O(G1180));
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );

  xor2  gate1471(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate1472(.a(gate405inter0), .b(s_132), .O(gate405inter1));
  and2  gate1473(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate1474(.a(s_132), .O(gate405inter3));
  inv1  gate1475(.a(s_133), .O(gate405inter4));
  nand2 gate1476(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate1477(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate1478(.a(G19), .O(gate405inter7));
  inv1  gate1479(.a(G1090), .O(gate405inter8));
  nand2 gate1480(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate1481(.a(s_133), .b(gate405inter3), .O(gate405inter10));
  nor2  gate1482(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate1483(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate1484(.a(gate405inter12), .b(gate405inter1), .O(G1186));
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate1093(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate1094(.a(gate411inter0), .b(s_78), .O(gate411inter1));
  and2  gate1095(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate1096(.a(s_78), .O(gate411inter3));
  inv1  gate1097(.a(s_79), .O(gate411inter4));
  nand2 gate1098(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate1099(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate1100(.a(G25), .O(gate411inter7));
  inv1  gate1101(.a(G1108), .O(gate411inter8));
  nand2 gate1102(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate1103(.a(s_79), .b(gate411inter3), .O(gate411inter10));
  nor2  gate1104(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate1105(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate1106(.a(gate411inter12), .b(gate411inter1), .O(G1204));

  xor2  gate1639(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate1640(.a(gate412inter0), .b(s_156), .O(gate412inter1));
  and2  gate1641(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate1642(.a(s_156), .O(gate412inter3));
  inv1  gate1643(.a(s_157), .O(gate412inter4));
  nand2 gate1644(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate1645(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate1646(.a(G26), .O(gate412inter7));
  inv1  gate1647(.a(G1111), .O(gate412inter8));
  nand2 gate1648(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate1649(.a(s_157), .b(gate412inter3), .O(gate412inter10));
  nor2  gate1650(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate1651(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate1652(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate2311(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate2312(.a(gate415inter0), .b(s_252), .O(gate415inter1));
  and2  gate2313(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate2314(.a(s_252), .O(gate415inter3));
  inv1  gate2315(.a(s_253), .O(gate415inter4));
  nand2 gate2316(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate2317(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate2318(.a(G29), .O(gate415inter7));
  inv1  gate2319(.a(G1120), .O(gate415inter8));
  nand2 gate2320(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate2321(.a(s_253), .b(gate415inter3), .O(gate415inter10));
  nor2  gate2322(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate2323(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate2324(.a(gate415inter12), .b(gate415inter1), .O(G1216));

  xor2  gate1709(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate1710(.a(gate416inter0), .b(s_166), .O(gate416inter1));
  and2  gate1711(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate1712(.a(s_166), .O(gate416inter3));
  inv1  gate1713(.a(s_167), .O(gate416inter4));
  nand2 gate1714(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate1715(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate1716(.a(G30), .O(gate416inter7));
  inv1  gate1717(.a(G1123), .O(gate416inter8));
  nand2 gate1718(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate1719(.a(s_167), .b(gate416inter3), .O(gate416inter10));
  nor2  gate1720(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate1721(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate1722(.a(gate416inter12), .b(gate416inter1), .O(G1219));
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate1359(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1360(.a(gate420inter0), .b(s_116), .O(gate420inter1));
  and2  gate1361(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1362(.a(s_116), .O(gate420inter3));
  inv1  gate1363(.a(s_117), .O(gate420inter4));
  nand2 gate1364(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1365(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1366(.a(G1036), .O(gate420inter7));
  inv1  gate1367(.a(G1132), .O(gate420inter8));
  nand2 gate1368(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1369(.a(s_117), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1370(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1371(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1372(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );

  xor2  gate687(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate688(.a(gate424inter0), .b(s_20), .O(gate424inter1));
  and2  gate689(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate690(.a(s_20), .O(gate424inter3));
  inv1  gate691(.a(s_21), .O(gate424inter4));
  nand2 gate692(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate693(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate694(.a(G1042), .O(gate424inter7));
  inv1  gate695(.a(G1138), .O(gate424inter8));
  nand2 gate696(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate697(.a(s_21), .b(gate424inter3), .O(gate424inter10));
  nor2  gate698(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate699(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate700(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate1821(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate1822(.a(gate432inter0), .b(s_182), .O(gate432inter1));
  and2  gate1823(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate1824(.a(s_182), .O(gate432inter3));
  inv1  gate1825(.a(s_183), .O(gate432inter4));
  nand2 gate1826(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate1827(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate1828(.a(G1054), .O(gate432inter7));
  inv1  gate1829(.a(G1150), .O(gate432inter8));
  nand2 gate1830(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate1831(.a(s_183), .b(gate432inter3), .O(gate432inter10));
  nor2  gate1832(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate1833(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate1834(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate827(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate828(.a(gate437inter0), .b(s_40), .O(gate437inter1));
  and2  gate829(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate830(.a(s_40), .O(gate437inter3));
  inv1  gate831(.a(s_41), .O(gate437inter4));
  nand2 gate832(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate833(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate834(.a(G10), .O(gate437inter7));
  inv1  gate835(.a(G1159), .O(gate437inter8));
  nand2 gate836(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate837(.a(s_41), .b(gate437inter3), .O(gate437inter10));
  nor2  gate838(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate839(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate840(.a(gate437inter12), .b(gate437inter1), .O(G1246));
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate1499(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate1500(.a(gate439inter0), .b(s_136), .O(gate439inter1));
  and2  gate1501(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate1502(.a(s_136), .O(gate439inter3));
  inv1  gate1503(.a(s_137), .O(gate439inter4));
  nand2 gate1504(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate1505(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate1506(.a(G11), .O(gate439inter7));
  inv1  gate1507(.a(G1162), .O(gate439inter8));
  nand2 gate1508(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate1509(.a(s_137), .b(gate439inter3), .O(gate439inter10));
  nor2  gate1510(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate1511(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate1512(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate1877(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate1878(.a(gate442inter0), .b(s_190), .O(gate442inter1));
  and2  gate1879(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate1880(.a(s_190), .O(gate442inter3));
  inv1  gate1881(.a(s_191), .O(gate442inter4));
  nand2 gate1882(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate1883(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate1884(.a(G1069), .O(gate442inter7));
  inv1  gate1885(.a(G1165), .O(gate442inter8));
  nand2 gate1886(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate1887(.a(s_191), .b(gate442inter3), .O(gate442inter10));
  nor2  gate1888(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate1889(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate1890(.a(gate442inter12), .b(gate442inter1), .O(G1251));

  xor2  gate1121(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate1122(.a(gate443inter0), .b(s_82), .O(gate443inter1));
  and2  gate1123(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate1124(.a(s_82), .O(gate443inter3));
  inv1  gate1125(.a(s_83), .O(gate443inter4));
  nand2 gate1126(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate1127(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate1128(.a(G13), .O(gate443inter7));
  inv1  gate1129(.a(G1168), .O(gate443inter8));
  nand2 gate1130(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate1131(.a(s_83), .b(gate443inter3), .O(gate443inter10));
  nor2  gate1132(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate1133(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate1134(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate925(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate926(.a(gate445inter0), .b(s_54), .O(gate445inter1));
  and2  gate927(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate928(.a(s_54), .O(gate445inter3));
  inv1  gate929(.a(s_55), .O(gate445inter4));
  nand2 gate930(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate931(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate932(.a(G14), .O(gate445inter7));
  inv1  gate933(.a(G1171), .O(gate445inter8));
  nand2 gate934(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate935(.a(s_55), .b(gate445inter3), .O(gate445inter10));
  nor2  gate936(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate937(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate938(.a(gate445inter12), .b(gate445inter1), .O(G1254));

  xor2  gate1149(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate1150(.a(gate446inter0), .b(s_86), .O(gate446inter1));
  and2  gate1151(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate1152(.a(s_86), .O(gate446inter3));
  inv1  gate1153(.a(s_87), .O(gate446inter4));
  nand2 gate1154(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate1155(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate1156(.a(G1075), .O(gate446inter7));
  inv1  gate1157(.a(G1171), .O(gate446inter8));
  nand2 gate1158(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate1159(.a(s_87), .b(gate446inter3), .O(gate446inter10));
  nor2  gate1160(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate1161(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate1162(.a(gate446inter12), .b(gate446inter1), .O(G1255));
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );

  xor2  gate1163(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate1164(.a(gate449inter0), .b(s_88), .O(gate449inter1));
  and2  gate1165(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate1166(.a(s_88), .O(gate449inter3));
  inv1  gate1167(.a(s_89), .O(gate449inter4));
  nand2 gate1168(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate1169(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate1170(.a(G16), .O(gate449inter7));
  inv1  gate1171(.a(G1177), .O(gate449inter8));
  nand2 gate1172(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate1173(.a(s_89), .b(gate449inter3), .O(gate449inter10));
  nor2  gate1174(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate1175(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate1176(.a(gate449inter12), .b(gate449inter1), .O(G1258));

  xor2  gate2045(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate2046(.a(gate450inter0), .b(s_214), .O(gate450inter1));
  and2  gate2047(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate2048(.a(s_214), .O(gate450inter3));
  inv1  gate2049(.a(s_215), .O(gate450inter4));
  nand2 gate2050(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate2051(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate2052(.a(G1081), .O(gate450inter7));
  inv1  gate2053(.a(G1177), .O(gate450inter8));
  nand2 gate2054(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate2055(.a(s_215), .b(gate450inter3), .O(gate450inter10));
  nor2  gate2056(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate2057(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate2058(.a(gate450inter12), .b(gate450inter1), .O(G1259));
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );

  xor2  gate2325(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate2326(.a(gate455inter0), .b(s_254), .O(gate455inter1));
  and2  gate2327(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate2328(.a(s_254), .O(gate455inter3));
  inv1  gate2329(.a(s_255), .O(gate455inter4));
  nand2 gate2330(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate2331(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate2332(.a(G19), .O(gate455inter7));
  inv1  gate2333(.a(G1186), .O(gate455inter8));
  nand2 gate2334(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate2335(.a(s_255), .b(gate455inter3), .O(gate455inter10));
  nor2  gate2336(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate2337(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate2338(.a(gate455inter12), .b(gate455inter1), .O(G1264));
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate1457(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate1458(.a(gate463inter0), .b(s_130), .O(gate463inter1));
  and2  gate1459(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate1460(.a(s_130), .O(gate463inter3));
  inv1  gate1461(.a(s_131), .O(gate463inter4));
  nand2 gate1462(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate1463(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate1464(.a(G23), .O(gate463inter7));
  inv1  gate1465(.a(G1198), .O(gate463inter8));
  nand2 gate1466(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate1467(.a(s_131), .b(gate463inter3), .O(gate463inter10));
  nor2  gate1468(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate1469(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate1470(.a(gate463inter12), .b(gate463inter1), .O(G1272));

  xor2  gate2227(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate2228(.a(gate464inter0), .b(s_240), .O(gate464inter1));
  and2  gate2229(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate2230(.a(s_240), .O(gate464inter3));
  inv1  gate2231(.a(s_241), .O(gate464inter4));
  nand2 gate2232(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate2233(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate2234(.a(G1102), .O(gate464inter7));
  inv1  gate2235(.a(G1198), .O(gate464inter8));
  nand2 gate2236(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate2237(.a(s_241), .b(gate464inter3), .O(gate464inter10));
  nor2  gate2238(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate2239(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate2240(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );

  xor2  gate2255(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate2256(.a(gate468inter0), .b(s_244), .O(gate468inter1));
  and2  gate2257(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate2258(.a(s_244), .O(gate468inter3));
  inv1  gate2259(.a(s_245), .O(gate468inter4));
  nand2 gate2260(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate2261(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate2262(.a(G1108), .O(gate468inter7));
  inv1  gate2263(.a(G1204), .O(gate468inter8));
  nand2 gate2264(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate2265(.a(s_245), .b(gate468inter3), .O(gate468inter10));
  nor2  gate2266(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate2267(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate2268(.a(gate468inter12), .b(gate468inter1), .O(G1277));

  xor2  gate2423(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate2424(.a(gate469inter0), .b(s_268), .O(gate469inter1));
  and2  gate2425(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate2426(.a(s_268), .O(gate469inter3));
  inv1  gate2427(.a(s_269), .O(gate469inter4));
  nand2 gate2428(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate2429(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate2430(.a(G26), .O(gate469inter7));
  inv1  gate2431(.a(G1207), .O(gate469inter8));
  nand2 gate2432(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate2433(.a(s_269), .b(gate469inter3), .O(gate469inter10));
  nor2  gate2434(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate2435(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate2436(.a(gate469inter12), .b(gate469inter1), .O(G1278));
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate911(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate912(.a(gate471inter0), .b(s_52), .O(gate471inter1));
  and2  gate913(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate914(.a(s_52), .O(gate471inter3));
  inv1  gate915(.a(s_53), .O(gate471inter4));
  nand2 gate916(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate917(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate918(.a(G27), .O(gate471inter7));
  inv1  gate919(.a(G1210), .O(gate471inter8));
  nand2 gate920(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate921(.a(s_53), .b(gate471inter3), .O(gate471inter10));
  nor2  gate922(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate923(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate924(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );

  xor2  gate561(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate562(.a(gate473inter0), .b(s_2), .O(gate473inter1));
  and2  gate563(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate564(.a(s_2), .O(gate473inter3));
  inv1  gate565(.a(s_3), .O(gate473inter4));
  nand2 gate566(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate567(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate568(.a(G28), .O(gate473inter7));
  inv1  gate569(.a(G1213), .O(gate473inter8));
  nand2 gate570(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate571(.a(s_3), .b(gate473inter3), .O(gate473inter10));
  nor2  gate572(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate573(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate574(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate2283(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate2284(.a(gate476inter0), .b(s_248), .O(gate476inter1));
  and2  gate2285(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate2286(.a(s_248), .O(gate476inter3));
  inv1  gate2287(.a(s_249), .O(gate476inter4));
  nand2 gate2288(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate2289(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate2290(.a(G1120), .O(gate476inter7));
  inv1  gate2291(.a(G1216), .O(gate476inter8));
  nand2 gate2292(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate2293(.a(s_249), .b(gate476inter3), .O(gate476inter10));
  nor2  gate2294(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate2295(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate2296(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );

  xor2  gate547(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate548(.a(gate479inter0), .b(s_0), .O(gate479inter1));
  and2  gate549(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate550(.a(s_0), .O(gate479inter3));
  inv1  gate551(.a(s_1), .O(gate479inter4));
  nand2 gate552(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate553(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate554(.a(G31), .O(gate479inter7));
  inv1  gate555(.a(G1222), .O(gate479inter8));
  nand2 gate556(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate557(.a(s_1), .b(gate479inter3), .O(gate479inter10));
  nor2  gate558(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate559(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate560(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate939(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate940(.a(gate481inter0), .b(s_56), .O(gate481inter1));
  and2  gate941(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate942(.a(s_56), .O(gate481inter3));
  inv1  gate943(.a(s_57), .O(gate481inter4));
  nand2 gate944(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate945(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate946(.a(G32), .O(gate481inter7));
  inv1  gate947(.a(G1225), .O(gate481inter8));
  nand2 gate948(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate949(.a(s_57), .b(gate481inter3), .O(gate481inter10));
  nor2  gate950(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate951(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate952(.a(gate481inter12), .b(gate481inter1), .O(G1290));
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate701(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate702(.a(gate490inter0), .b(s_22), .O(gate490inter1));
  and2  gate703(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate704(.a(s_22), .O(gate490inter3));
  inv1  gate705(.a(s_23), .O(gate490inter4));
  nand2 gate706(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate707(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate708(.a(G1242), .O(gate490inter7));
  inv1  gate709(.a(G1243), .O(gate490inter8));
  nand2 gate710(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate711(.a(s_23), .b(gate490inter3), .O(gate490inter10));
  nor2  gate712(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate713(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate714(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate2003(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate2004(.a(gate492inter0), .b(s_208), .O(gate492inter1));
  and2  gate2005(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate2006(.a(s_208), .O(gate492inter3));
  inv1  gate2007(.a(s_209), .O(gate492inter4));
  nand2 gate2008(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate2009(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate2010(.a(G1246), .O(gate492inter7));
  inv1  gate2011(.a(G1247), .O(gate492inter8));
  nand2 gate2012(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate2013(.a(s_209), .b(gate492inter3), .O(gate492inter10));
  nor2  gate2014(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate2015(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate2016(.a(gate492inter12), .b(gate492inter1), .O(G1301));

  xor2  gate1079(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate1080(.a(gate493inter0), .b(s_76), .O(gate493inter1));
  and2  gate1081(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate1082(.a(s_76), .O(gate493inter3));
  inv1  gate1083(.a(s_77), .O(gate493inter4));
  nand2 gate1084(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate1085(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate1086(.a(G1248), .O(gate493inter7));
  inv1  gate1087(.a(G1249), .O(gate493inter8));
  nand2 gate1088(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate1089(.a(s_77), .b(gate493inter3), .O(gate493inter10));
  nor2  gate1090(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate1091(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate1092(.a(gate493inter12), .b(gate493inter1), .O(G1302));
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );

  xor2  gate1443(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate1444(.a(gate495inter0), .b(s_128), .O(gate495inter1));
  and2  gate1445(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate1446(.a(s_128), .O(gate495inter3));
  inv1  gate1447(.a(s_129), .O(gate495inter4));
  nand2 gate1448(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate1449(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate1450(.a(G1252), .O(gate495inter7));
  inv1  gate1451(.a(G1253), .O(gate495inter8));
  nand2 gate1452(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate1453(.a(s_129), .b(gate495inter3), .O(gate495inter10));
  nor2  gate1454(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate1455(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate1456(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );

  xor2  gate1485(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate1486(.a(gate498inter0), .b(s_134), .O(gate498inter1));
  and2  gate1487(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate1488(.a(s_134), .O(gate498inter3));
  inv1  gate1489(.a(s_135), .O(gate498inter4));
  nand2 gate1490(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate1491(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate1492(.a(G1258), .O(gate498inter7));
  inv1  gate1493(.a(G1259), .O(gate498inter8));
  nand2 gate1494(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate1495(.a(s_135), .b(gate498inter3), .O(gate498inter10));
  nor2  gate1496(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate1497(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate1498(.a(gate498inter12), .b(gate498inter1), .O(G1307));
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate1373(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate1374(.a(gate502inter0), .b(s_118), .O(gate502inter1));
  and2  gate1375(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate1376(.a(s_118), .O(gate502inter3));
  inv1  gate1377(.a(s_119), .O(gate502inter4));
  nand2 gate1378(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate1379(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate1380(.a(G1266), .O(gate502inter7));
  inv1  gate1381(.a(G1267), .O(gate502inter8));
  nand2 gate1382(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate1383(.a(s_119), .b(gate502inter3), .O(gate502inter10));
  nor2  gate1384(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate1385(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate1386(.a(gate502inter12), .b(gate502inter1), .O(G1311));

  xor2  gate2185(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate2186(.a(gate503inter0), .b(s_234), .O(gate503inter1));
  and2  gate2187(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate2188(.a(s_234), .O(gate503inter3));
  inv1  gate2189(.a(s_235), .O(gate503inter4));
  nand2 gate2190(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate2191(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate2192(.a(G1268), .O(gate503inter7));
  inv1  gate2193(.a(G1269), .O(gate503inter8));
  nand2 gate2194(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate2195(.a(s_235), .b(gate503inter3), .O(gate503inter10));
  nor2  gate2196(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate2197(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate2198(.a(gate503inter12), .b(gate503inter1), .O(G1312));

  xor2  gate729(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate730(.a(gate504inter0), .b(s_26), .O(gate504inter1));
  and2  gate731(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate732(.a(s_26), .O(gate504inter3));
  inv1  gate733(.a(s_27), .O(gate504inter4));
  nand2 gate734(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate735(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate736(.a(G1270), .O(gate504inter7));
  inv1  gate737(.a(G1271), .O(gate504inter8));
  nand2 gate738(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate739(.a(s_27), .b(gate504inter3), .O(gate504inter10));
  nor2  gate740(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate741(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate742(.a(gate504inter12), .b(gate504inter1), .O(G1313));

  xor2  gate645(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate646(.a(gate505inter0), .b(s_14), .O(gate505inter1));
  and2  gate647(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate648(.a(s_14), .O(gate505inter3));
  inv1  gate649(.a(s_15), .O(gate505inter4));
  nand2 gate650(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate651(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate652(.a(G1272), .O(gate505inter7));
  inv1  gate653(.a(G1273), .O(gate505inter8));
  nand2 gate654(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate655(.a(s_15), .b(gate505inter3), .O(gate505inter10));
  nor2  gate656(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate657(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate658(.a(gate505inter12), .b(gate505inter1), .O(G1314));

  xor2  gate869(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate870(.a(gate506inter0), .b(s_46), .O(gate506inter1));
  and2  gate871(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate872(.a(s_46), .O(gate506inter3));
  inv1  gate873(.a(s_47), .O(gate506inter4));
  nand2 gate874(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate875(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate876(.a(G1274), .O(gate506inter7));
  inv1  gate877(.a(G1275), .O(gate506inter8));
  nand2 gate878(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate879(.a(s_47), .b(gate506inter3), .O(gate506inter10));
  nor2  gate880(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate881(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate882(.a(gate506inter12), .b(gate506inter1), .O(G1315));

  xor2  gate1247(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate1248(.a(gate507inter0), .b(s_100), .O(gate507inter1));
  and2  gate1249(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate1250(.a(s_100), .O(gate507inter3));
  inv1  gate1251(.a(s_101), .O(gate507inter4));
  nand2 gate1252(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate1253(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate1254(.a(G1276), .O(gate507inter7));
  inv1  gate1255(.a(G1277), .O(gate507inter8));
  nand2 gate1256(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate1257(.a(s_101), .b(gate507inter3), .O(gate507inter10));
  nor2  gate1258(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate1259(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate1260(.a(gate507inter12), .b(gate507inter1), .O(G1316));

  xor2  gate1597(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate1598(.a(gate508inter0), .b(s_150), .O(gate508inter1));
  and2  gate1599(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate1600(.a(s_150), .O(gate508inter3));
  inv1  gate1601(.a(s_151), .O(gate508inter4));
  nand2 gate1602(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate1603(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate1604(.a(G1278), .O(gate508inter7));
  inv1  gate1605(.a(G1279), .O(gate508inter8));
  nand2 gate1606(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate1607(.a(s_151), .b(gate508inter3), .O(gate508inter10));
  nor2  gate1608(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate1609(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate1610(.a(gate508inter12), .b(gate508inter1), .O(G1317));

  xor2  gate1695(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate1696(.a(gate509inter0), .b(s_164), .O(gate509inter1));
  and2  gate1697(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate1698(.a(s_164), .O(gate509inter3));
  inv1  gate1699(.a(s_165), .O(gate509inter4));
  nand2 gate1700(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate1701(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate1702(.a(G1280), .O(gate509inter7));
  inv1  gate1703(.a(G1281), .O(gate509inter8));
  nand2 gate1704(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate1705(.a(s_165), .b(gate509inter3), .O(gate509inter10));
  nor2  gate1706(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate1707(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate1708(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate603(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate604(.a(gate511inter0), .b(s_8), .O(gate511inter1));
  and2  gate605(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate606(.a(s_8), .O(gate511inter3));
  inv1  gate607(.a(s_9), .O(gate511inter4));
  nand2 gate608(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate609(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate610(.a(G1284), .O(gate511inter7));
  inv1  gate611(.a(G1285), .O(gate511inter8));
  nand2 gate612(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate613(.a(s_9), .b(gate511inter3), .O(gate511inter10));
  nor2  gate614(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate615(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate616(.a(gate511inter12), .b(gate511inter1), .O(G1320));

  xor2  gate1583(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate1584(.a(gate512inter0), .b(s_148), .O(gate512inter1));
  and2  gate1585(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate1586(.a(s_148), .O(gate512inter3));
  inv1  gate1587(.a(s_149), .O(gate512inter4));
  nand2 gate1588(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate1589(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate1590(.a(G1286), .O(gate512inter7));
  inv1  gate1591(.a(G1287), .O(gate512inter8));
  nand2 gate1592(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate1593(.a(s_149), .b(gate512inter3), .O(gate512inter10));
  nor2  gate1594(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate1595(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate1596(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule