module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate841(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate842(.a(gate28inter0), .b(s_42), .O(gate28inter1));
  and2  gate843(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate844(.a(s_42), .O(gate28inter3));
  inv1  gate845(.a(s_43), .O(gate28inter4));
  nand2 gate846(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate847(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate848(.a(G10), .O(gate28inter7));
  inv1  gate849(.a(G14), .O(gate28inter8));
  nand2 gate850(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate851(.a(s_43), .b(gate28inter3), .O(gate28inter10));
  nor2  gate852(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate853(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate854(.a(gate28inter12), .b(gate28inter1), .O(G323));
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate1429(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1430(.a(gate36inter0), .b(s_126), .O(gate36inter1));
  and2  gate1431(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1432(.a(s_126), .O(gate36inter3));
  inv1  gate1433(.a(s_127), .O(gate36inter4));
  nand2 gate1434(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1435(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1436(.a(G26), .O(gate36inter7));
  inv1  gate1437(.a(G30), .O(gate36inter8));
  nand2 gate1438(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1439(.a(s_127), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1440(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1441(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1442(.a(gate36inter12), .b(gate36inter1), .O(G347));

  xor2  gate1653(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate1654(.a(gate37inter0), .b(s_158), .O(gate37inter1));
  and2  gate1655(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate1656(.a(s_158), .O(gate37inter3));
  inv1  gate1657(.a(s_159), .O(gate37inter4));
  nand2 gate1658(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate1659(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate1660(.a(G19), .O(gate37inter7));
  inv1  gate1661(.a(G23), .O(gate37inter8));
  nand2 gate1662(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate1663(.a(s_159), .b(gate37inter3), .O(gate37inter10));
  nor2  gate1664(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate1665(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate1666(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate1765(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate1766(.a(gate51inter0), .b(s_174), .O(gate51inter1));
  and2  gate1767(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate1768(.a(s_174), .O(gate51inter3));
  inv1  gate1769(.a(s_175), .O(gate51inter4));
  nand2 gate1770(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate1771(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate1772(.a(G11), .O(gate51inter7));
  inv1  gate1773(.a(G281), .O(gate51inter8));
  nand2 gate1774(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate1775(.a(s_175), .b(gate51inter3), .O(gate51inter10));
  nor2  gate1776(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate1777(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate1778(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );

  xor2  gate757(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate758(.a(gate56inter0), .b(s_30), .O(gate56inter1));
  and2  gate759(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate760(.a(s_30), .O(gate56inter3));
  inv1  gate761(.a(s_31), .O(gate56inter4));
  nand2 gate762(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate763(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate764(.a(G16), .O(gate56inter7));
  inv1  gate765(.a(G287), .O(gate56inter8));
  nand2 gate766(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate767(.a(s_31), .b(gate56inter3), .O(gate56inter10));
  nor2  gate768(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate769(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate770(.a(gate56inter12), .b(gate56inter1), .O(G377));

  xor2  gate743(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate744(.a(gate57inter0), .b(s_28), .O(gate57inter1));
  and2  gate745(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate746(.a(s_28), .O(gate57inter3));
  inv1  gate747(.a(s_29), .O(gate57inter4));
  nand2 gate748(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate749(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate750(.a(G17), .O(gate57inter7));
  inv1  gate751(.a(G290), .O(gate57inter8));
  nand2 gate752(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate753(.a(s_29), .b(gate57inter3), .O(gate57inter10));
  nor2  gate754(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate755(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate756(.a(gate57inter12), .b(gate57inter1), .O(G378));

  xor2  gate1023(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate1024(.a(gate58inter0), .b(s_68), .O(gate58inter1));
  and2  gate1025(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate1026(.a(s_68), .O(gate58inter3));
  inv1  gate1027(.a(s_69), .O(gate58inter4));
  nand2 gate1028(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate1029(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate1030(.a(G18), .O(gate58inter7));
  inv1  gate1031(.a(G290), .O(gate58inter8));
  nand2 gate1032(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate1033(.a(s_69), .b(gate58inter3), .O(gate58inter10));
  nor2  gate1034(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate1035(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate1036(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate547(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate548(.a(gate63inter0), .b(s_0), .O(gate63inter1));
  and2  gate549(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate550(.a(s_0), .O(gate63inter3));
  inv1  gate551(.a(s_1), .O(gate63inter4));
  nand2 gate552(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate553(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate554(.a(G23), .O(gate63inter7));
  inv1  gate555(.a(G299), .O(gate63inter8));
  nand2 gate556(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate557(.a(s_1), .b(gate63inter3), .O(gate63inter10));
  nor2  gate558(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate559(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate560(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );

  xor2  gate911(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate912(.a(gate68inter0), .b(s_52), .O(gate68inter1));
  and2  gate913(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate914(.a(s_52), .O(gate68inter3));
  inv1  gate915(.a(s_53), .O(gate68inter4));
  nand2 gate916(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate917(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate918(.a(G28), .O(gate68inter7));
  inv1  gate919(.a(G305), .O(gate68inter8));
  nand2 gate920(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate921(.a(s_53), .b(gate68inter3), .O(gate68inter10));
  nor2  gate922(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate923(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate924(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate1093(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate1094(.a(gate70inter0), .b(s_78), .O(gate70inter1));
  and2  gate1095(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate1096(.a(s_78), .O(gate70inter3));
  inv1  gate1097(.a(s_79), .O(gate70inter4));
  nand2 gate1098(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate1099(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate1100(.a(G30), .O(gate70inter7));
  inv1  gate1101(.a(G308), .O(gate70inter8));
  nand2 gate1102(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate1103(.a(s_79), .b(gate70inter3), .O(gate70inter10));
  nor2  gate1104(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate1105(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate1106(.a(gate70inter12), .b(gate70inter1), .O(G391));

  xor2  gate1247(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate1248(.a(gate71inter0), .b(s_100), .O(gate71inter1));
  and2  gate1249(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate1250(.a(s_100), .O(gate71inter3));
  inv1  gate1251(.a(s_101), .O(gate71inter4));
  nand2 gate1252(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate1253(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate1254(.a(G31), .O(gate71inter7));
  inv1  gate1255(.a(G311), .O(gate71inter8));
  nand2 gate1256(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate1257(.a(s_101), .b(gate71inter3), .O(gate71inter10));
  nor2  gate1258(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate1259(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate1260(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate1219(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate1220(.a(gate85inter0), .b(s_96), .O(gate85inter1));
  and2  gate1221(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate1222(.a(s_96), .O(gate85inter3));
  inv1  gate1223(.a(s_97), .O(gate85inter4));
  nand2 gate1224(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate1225(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate1226(.a(G4), .O(gate85inter7));
  inv1  gate1227(.a(G332), .O(gate85inter8));
  nand2 gate1228(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate1229(.a(s_97), .b(gate85inter3), .O(gate85inter10));
  nor2  gate1230(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate1231(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate1232(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );

  xor2  gate1625(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate1626(.a(gate89inter0), .b(s_154), .O(gate89inter1));
  and2  gate1627(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate1628(.a(s_154), .O(gate89inter3));
  inv1  gate1629(.a(s_155), .O(gate89inter4));
  nand2 gate1630(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate1631(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate1632(.a(G17), .O(gate89inter7));
  inv1  gate1633(.a(G338), .O(gate89inter8));
  nand2 gate1634(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate1635(.a(s_155), .b(gate89inter3), .O(gate89inter10));
  nor2  gate1636(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate1637(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate1638(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );

  xor2  gate1233(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate1234(.a(gate93inter0), .b(s_98), .O(gate93inter1));
  and2  gate1235(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate1236(.a(s_98), .O(gate93inter3));
  inv1  gate1237(.a(s_99), .O(gate93inter4));
  nand2 gate1238(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate1239(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate1240(.a(G18), .O(gate93inter7));
  inv1  gate1241(.a(G344), .O(gate93inter8));
  nand2 gate1242(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate1243(.a(s_99), .b(gate93inter3), .O(gate93inter10));
  nor2  gate1244(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate1245(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate1246(.a(gate93inter12), .b(gate93inter1), .O(G414));
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate1317(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate1318(.a(gate100inter0), .b(s_110), .O(gate100inter1));
  and2  gate1319(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate1320(.a(s_110), .O(gate100inter3));
  inv1  gate1321(.a(s_111), .O(gate100inter4));
  nand2 gate1322(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate1323(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate1324(.a(G31), .O(gate100inter7));
  inv1  gate1325(.a(G353), .O(gate100inter8));
  nand2 gate1326(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate1327(.a(s_111), .b(gate100inter3), .O(gate100inter10));
  nor2  gate1328(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate1329(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate1330(.a(gate100inter12), .b(gate100inter1), .O(G421));

  xor2  gate897(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate898(.a(gate101inter0), .b(s_50), .O(gate101inter1));
  and2  gate899(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate900(.a(s_50), .O(gate101inter3));
  inv1  gate901(.a(s_51), .O(gate101inter4));
  nand2 gate902(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate903(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate904(.a(G20), .O(gate101inter7));
  inv1  gate905(.a(G356), .O(gate101inter8));
  nand2 gate906(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate907(.a(s_51), .b(gate101inter3), .O(gate101inter10));
  nor2  gate908(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate909(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate910(.a(gate101inter12), .b(gate101inter1), .O(G422));

  xor2  gate1079(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate1080(.a(gate102inter0), .b(s_76), .O(gate102inter1));
  and2  gate1081(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate1082(.a(s_76), .O(gate102inter3));
  inv1  gate1083(.a(s_77), .O(gate102inter4));
  nand2 gate1084(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate1085(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate1086(.a(G24), .O(gate102inter7));
  inv1  gate1087(.a(G356), .O(gate102inter8));
  nand2 gate1088(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate1089(.a(s_77), .b(gate102inter3), .O(gate102inter10));
  nor2  gate1090(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate1091(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate1092(.a(gate102inter12), .b(gate102inter1), .O(G423));

  xor2  gate967(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate968(.a(gate103inter0), .b(s_60), .O(gate103inter1));
  and2  gate969(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate970(.a(s_60), .O(gate103inter3));
  inv1  gate971(.a(s_61), .O(gate103inter4));
  nand2 gate972(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate973(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate974(.a(G28), .O(gate103inter7));
  inv1  gate975(.a(G359), .O(gate103inter8));
  nand2 gate976(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate977(.a(s_61), .b(gate103inter3), .O(gate103inter10));
  nor2  gate978(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate979(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate980(.a(gate103inter12), .b(gate103inter1), .O(G424));

  xor2  gate715(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate716(.a(gate104inter0), .b(s_24), .O(gate104inter1));
  and2  gate717(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate718(.a(s_24), .O(gate104inter3));
  inv1  gate719(.a(s_25), .O(gate104inter4));
  nand2 gate720(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate721(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate722(.a(G32), .O(gate104inter7));
  inv1  gate723(.a(G359), .O(gate104inter8));
  nand2 gate724(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate725(.a(s_25), .b(gate104inter3), .O(gate104inter10));
  nor2  gate726(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate727(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate728(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate1345(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate1346(.a(gate108inter0), .b(s_114), .O(gate108inter1));
  and2  gate1347(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate1348(.a(s_114), .O(gate108inter3));
  inv1  gate1349(.a(s_115), .O(gate108inter4));
  nand2 gate1350(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate1351(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate1352(.a(G368), .O(gate108inter7));
  inv1  gate1353(.a(G369), .O(gate108inter8));
  nand2 gate1354(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate1355(.a(s_115), .b(gate108inter3), .O(gate108inter10));
  nor2  gate1356(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate1357(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate1358(.a(gate108inter12), .b(gate108inter1), .O(G435));
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate883(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate884(.a(gate112inter0), .b(s_48), .O(gate112inter1));
  and2  gate885(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate886(.a(s_48), .O(gate112inter3));
  inv1  gate887(.a(s_49), .O(gate112inter4));
  nand2 gate888(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate889(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate890(.a(G376), .O(gate112inter7));
  inv1  gate891(.a(G377), .O(gate112inter8));
  nand2 gate892(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate893(.a(s_49), .b(gate112inter3), .O(gate112inter10));
  nor2  gate894(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate895(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate896(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate659(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate660(.a(gate118inter0), .b(s_16), .O(gate118inter1));
  and2  gate661(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate662(.a(s_16), .O(gate118inter3));
  inv1  gate663(.a(s_17), .O(gate118inter4));
  nand2 gate664(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate665(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate666(.a(G388), .O(gate118inter7));
  inv1  gate667(.a(G389), .O(gate118inter8));
  nand2 gate668(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate669(.a(s_17), .b(gate118inter3), .O(gate118inter10));
  nor2  gate670(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate671(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate672(.a(gate118inter12), .b(gate118inter1), .O(G465));
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate995(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate996(.a(gate121inter0), .b(s_64), .O(gate121inter1));
  and2  gate997(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate998(.a(s_64), .O(gate121inter3));
  inv1  gate999(.a(s_65), .O(gate121inter4));
  nand2 gate1000(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate1001(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate1002(.a(G394), .O(gate121inter7));
  inv1  gate1003(.a(G395), .O(gate121inter8));
  nand2 gate1004(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate1005(.a(s_65), .b(gate121inter3), .O(gate121inter10));
  nor2  gate1006(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate1007(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate1008(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate617(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate618(.a(gate124inter0), .b(s_10), .O(gate124inter1));
  and2  gate619(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate620(.a(s_10), .O(gate124inter3));
  inv1  gate621(.a(s_11), .O(gate124inter4));
  nand2 gate622(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate623(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate624(.a(G400), .O(gate124inter7));
  inv1  gate625(.a(G401), .O(gate124inter8));
  nand2 gate626(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate627(.a(s_11), .b(gate124inter3), .O(gate124inter10));
  nor2  gate628(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate629(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate630(.a(gate124inter12), .b(gate124inter1), .O(G483));

  xor2  gate1191(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate1192(.a(gate125inter0), .b(s_92), .O(gate125inter1));
  and2  gate1193(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate1194(.a(s_92), .O(gate125inter3));
  inv1  gate1195(.a(s_93), .O(gate125inter4));
  nand2 gate1196(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate1197(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate1198(.a(G402), .O(gate125inter7));
  inv1  gate1199(.a(G403), .O(gate125inter8));
  nand2 gate1200(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate1201(.a(s_93), .b(gate125inter3), .O(gate125inter10));
  nor2  gate1202(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate1203(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate1204(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate701(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate702(.a(gate130inter0), .b(s_22), .O(gate130inter1));
  and2  gate703(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate704(.a(s_22), .O(gate130inter3));
  inv1  gate705(.a(s_23), .O(gate130inter4));
  nand2 gate706(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate707(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate708(.a(G412), .O(gate130inter7));
  inv1  gate709(.a(G413), .O(gate130inter8));
  nand2 gate710(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate711(.a(s_23), .b(gate130inter3), .O(gate130inter10));
  nor2  gate712(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate713(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate714(.a(gate130inter12), .b(gate130inter1), .O(G501));
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate645(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate646(.a(gate132inter0), .b(s_14), .O(gate132inter1));
  and2  gate647(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate648(.a(s_14), .O(gate132inter3));
  inv1  gate649(.a(s_15), .O(gate132inter4));
  nand2 gate650(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate651(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate652(.a(G416), .O(gate132inter7));
  inv1  gate653(.a(G417), .O(gate132inter8));
  nand2 gate654(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate655(.a(s_15), .b(gate132inter3), .O(gate132inter10));
  nor2  gate656(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate657(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate658(.a(gate132inter12), .b(gate132inter1), .O(G507));

  xor2  gate589(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate590(.a(gate133inter0), .b(s_6), .O(gate133inter1));
  and2  gate591(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate592(.a(s_6), .O(gate133inter3));
  inv1  gate593(.a(s_7), .O(gate133inter4));
  nand2 gate594(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate595(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate596(.a(G418), .O(gate133inter7));
  inv1  gate597(.a(G419), .O(gate133inter8));
  nand2 gate598(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate599(.a(s_7), .b(gate133inter3), .O(gate133inter10));
  nor2  gate600(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate601(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate602(.a(gate133inter12), .b(gate133inter1), .O(G510));
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );

  xor2  gate1513(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate1514(.a(gate145inter0), .b(s_138), .O(gate145inter1));
  and2  gate1515(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate1516(.a(s_138), .O(gate145inter3));
  inv1  gate1517(.a(s_139), .O(gate145inter4));
  nand2 gate1518(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate1519(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate1520(.a(G474), .O(gate145inter7));
  inv1  gate1521(.a(G477), .O(gate145inter8));
  nand2 gate1522(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate1523(.a(s_139), .b(gate145inter3), .O(gate145inter10));
  nor2  gate1524(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate1525(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate1526(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate981(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate982(.a(gate149inter0), .b(s_62), .O(gate149inter1));
  and2  gate983(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate984(.a(s_62), .O(gate149inter3));
  inv1  gate985(.a(s_63), .O(gate149inter4));
  nand2 gate986(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate987(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate988(.a(G498), .O(gate149inter7));
  inv1  gate989(.a(G501), .O(gate149inter8));
  nand2 gate990(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate991(.a(s_63), .b(gate149inter3), .O(gate149inter10));
  nor2  gate992(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate993(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate994(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );

  xor2  gate1135(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate1136(.a(gate152inter0), .b(s_84), .O(gate152inter1));
  and2  gate1137(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate1138(.a(s_84), .O(gate152inter3));
  inv1  gate1139(.a(s_85), .O(gate152inter4));
  nand2 gate1140(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate1141(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate1142(.a(G516), .O(gate152inter7));
  inv1  gate1143(.a(G519), .O(gate152inter8));
  nand2 gate1144(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate1145(.a(s_85), .b(gate152inter3), .O(gate152inter10));
  nor2  gate1146(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate1147(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate1148(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate1387(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate1388(.a(gate154inter0), .b(s_120), .O(gate154inter1));
  and2  gate1389(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate1390(.a(s_120), .O(gate154inter3));
  inv1  gate1391(.a(s_121), .O(gate154inter4));
  nand2 gate1392(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate1393(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate1394(.a(G429), .O(gate154inter7));
  inv1  gate1395(.a(G522), .O(gate154inter8));
  nand2 gate1396(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate1397(.a(s_121), .b(gate154inter3), .O(gate154inter10));
  nor2  gate1398(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate1399(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate1400(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate1401(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate1402(.a(gate156inter0), .b(s_122), .O(gate156inter1));
  and2  gate1403(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate1404(.a(s_122), .O(gate156inter3));
  inv1  gate1405(.a(s_123), .O(gate156inter4));
  nand2 gate1406(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate1407(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate1408(.a(G435), .O(gate156inter7));
  inv1  gate1409(.a(G525), .O(gate156inter8));
  nand2 gate1410(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate1411(.a(s_123), .b(gate156inter3), .O(gate156inter10));
  nor2  gate1412(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate1413(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate1414(.a(gate156inter12), .b(gate156inter1), .O(G573));

  xor2  gate673(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate674(.a(gate157inter0), .b(s_18), .O(gate157inter1));
  and2  gate675(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate676(.a(s_18), .O(gate157inter3));
  inv1  gate677(.a(s_19), .O(gate157inter4));
  nand2 gate678(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate679(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate680(.a(G438), .O(gate157inter7));
  inv1  gate681(.a(G528), .O(gate157inter8));
  nand2 gate682(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate683(.a(s_19), .b(gate157inter3), .O(gate157inter10));
  nor2  gate684(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate685(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate686(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );

  xor2  gate1177(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate1178(.a(gate163inter0), .b(s_90), .O(gate163inter1));
  and2  gate1179(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate1180(.a(s_90), .O(gate163inter3));
  inv1  gate1181(.a(s_91), .O(gate163inter4));
  nand2 gate1182(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate1183(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate1184(.a(G456), .O(gate163inter7));
  inv1  gate1185(.a(G537), .O(gate163inter8));
  nand2 gate1186(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate1187(.a(s_91), .b(gate163inter3), .O(gate163inter10));
  nor2  gate1188(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate1189(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate1190(.a(gate163inter12), .b(gate163inter1), .O(G580));
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );

  xor2  gate1065(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate1066(.a(gate176inter0), .b(s_74), .O(gate176inter1));
  and2  gate1067(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate1068(.a(s_74), .O(gate176inter3));
  inv1  gate1069(.a(s_75), .O(gate176inter4));
  nand2 gate1070(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate1071(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate1072(.a(G495), .O(gate176inter7));
  inv1  gate1073(.a(G555), .O(gate176inter8));
  nand2 gate1074(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate1075(.a(s_75), .b(gate176inter3), .O(gate176inter10));
  nor2  gate1076(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate1077(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate1078(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate1051(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate1052(.a(gate178inter0), .b(s_72), .O(gate178inter1));
  and2  gate1053(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate1054(.a(s_72), .O(gate178inter3));
  inv1  gate1055(.a(s_73), .O(gate178inter4));
  nand2 gate1056(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate1057(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate1058(.a(G501), .O(gate178inter7));
  inv1  gate1059(.a(G558), .O(gate178inter8));
  nand2 gate1060(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate1061(.a(s_73), .b(gate178inter3), .O(gate178inter10));
  nor2  gate1062(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate1063(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate1064(.a(gate178inter12), .b(gate178inter1), .O(G595));
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );

  xor2  gate1457(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate1458(.a(gate189inter0), .b(s_130), .O(gate189inter1));
  and2  gate1459(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate1460(.a(s_130), .O(gate189inter3));
  inv1  gate1461(.a(s_131), .O(gate189inter4));
  nand2 gate1462(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate1463(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate1464(.a(G578), .O(gate189inter7));
  inv1  gate1465(.a(G579), .O(gate189inter8));
  nand2 gate1466(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate1467(.a(s_131), .b(gate189inter3), .O(gate189inter10));
  nor2  gate1468(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate1469(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate1470(.a(gate189inter12), .b(gate189inter1), .O(G622));
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate561(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate562(.a(gate191inter0), .b(s_2), .O(gate191inter1));
  and2  gate563(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate564(.a(s_2), .O(gate191inter3));
  inv1  gate565(.a(s_3), .O(gate191inter4));
  nand2 gate566(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate567(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate568(.a(G582), .O(gate191inter7));
  inv1  gate569(.a(G583), .O(gate191inter8));
  nand2 gate570(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate571(.a(s_3), .b(gate191inter3), .O(gate191inter10));
  nor2  gate572(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate573(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate574(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate869(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate870(.a(gate200inter0), .b(s_46), .O(gate200inter1));
  and2  gate871(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate872(.a(s_46), .O(gate200inter3));
  inv1  gate873(.a(s_47), .O(gate200inter4));
  nand2 gate874(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate875(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate876(.a(G600), .O(gate200inter7));
  inv1  gate877(.a(G601), .O(gate200inter8));
  nand2 gate878(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate879(.a(s_47), .b(gate200inter3), .O(gate200inter10));
  nor2  gate880(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate881(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate882(.a(gate200inter12), .b(gate200inter1), .O(G663));
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate1793(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate1794(.a(gate211inter0), .b(s_178), .O(gate211inter1));
  and2  gate1795(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate1796(.a(s_178), .O(gate211inter3));
  inv1  gate1797(.a(s_179), .O(gate211inter4));
  nand2 gate1798(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate1799(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate1800(.a(G612), .O(gate211inter7));
  inv1  gate1801(.a(G669), .O(gate211inter8));
  nand2 gate1802(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate1803(.a(s_179), .b(gate211inter3), .O(gate211inter10));
  nor2  gate1804(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate1805(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate1806(.a(gate211inter12), .b(gate211inter1), .O(G692));

  xor2  gate771(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate772(.a(gate212inter0), .b(s_32), .O(gate212inter1));
  and2  gate773(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate774(.a(s_32), .O(gate212inter3));
  inv1  gate775(.a(s_33), .O(gate212inter4));
  nand2 gate776(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate777(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate778(.a(G617), .O(gate212inter7));
  inv1  gate779(.a(G669), .O(gate212inter8));
  nand2 gate780(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate781(.a(s_33), .b(gate212inter3), .O(gate212inter10));
  nor2  gate782(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate783(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate784(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate1751(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate1752(.a(gate214inter0), .b(s_172), .O(gate214inter1));
  and2  gate1753(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate1754(.a(s_172), .O(gate214inter3));
  inv1  gate1755(.a(s_173), .O(gate214inter4));
  nand2 gate1756(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate1757(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate1758(.a(G612), .O(gate214inter7));
  inv1  gate1759(.a(G672), .O(gate214inter8));
  nand2 gate1760(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate1761(.a(s_173), .b(gate214inter3), .O(gate214inter10));
  nor2  gate1762(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate1763(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate1764(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate1779(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate1780(.a(gate220inter0), .b(s_176), .O(gate220inter1));
  and2  gate1781(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate1782(.a(s_176), .O(gate220inter3));
  inv1  gate1783(.a(s_177), .O(gate220inter4));
  nand2 gate1784(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate1785(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate1786(.a(G637), .O(gate220inter7));
  inv1  gate1787(.a(G681), .O(gate220inter8));
  nand2 gate1788(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate1789(.a(s_177), .b(gate220inter3), .O(gate220inter10));
  nor2  gate1790(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate1791(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate1792(.a(gate220inter12), .b(gate220inter1), .O(G701));
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate1583(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate1584(.a(gate223inter0), .b(s_148), .O(gate223inter1));
  and2  gate1585(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate1586(.a(s_148), .O(gate223inter3));
  inv1  gate1587(.a(s_149), .O(gate223inter4));
  nand2 gate1588(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate1589(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate1590(.a(G627), .O(gate223inter7));
  inv1  gate1591(.a(G687), .O(gate223inter8));
  nand2 gate1592(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate1593(.a(s_149), .b(gate223inter3), .O(gate223inter10));
  nor2  gate1594(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate1595(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate1596(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate1485(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate1486(.a(gate226inter0), .b(s_134), .O(gate226inter1));
  and2  gate1487(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate1488(.a(s_134), .O(gate226inter3));
  inv1  gate1489(.a(s_135), .O(gate226inter4));
  nand2 gate1490(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate1491(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate1492(.a(G692), .O(gate226inter7));
  inv1  gate1493(.a(G693), .O(gate226inter8));
  nand2 gate1494(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate1495(.a(s_135), .b(gate226inter3), .O(gate226inter10));
  nor2  gate1496(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate1497(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate1498(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate1163(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate1164(.a(gate231inter0), .b(s_88), .O(gate231inter1));
  and2  gate1165(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate1166(.a(s_88), .O(gate231inter3));
  inv1  gate1167(.a(s_89), .O(gate231inter4));
  nand2 gate1168(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate1169(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate1170(.a(G702), .O(gate231inter7));
  inv1  gate1171(.a(G703), .O(gate231inter8));
  nand2 gate1172(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate1173(.a(s_89), .b(gate231inter3), .O(gate231inter10));
  nor2  gate1174(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate1175(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate1176(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate785(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate786(.a(gate236inter0), .b(s_34), .O(gate236inter1));
  and2  gate787(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate788(.a(s_34), .O(gate236inter3));
  inv1  gate789(.a(s_35), .O(gate236inter4));
  nand2 gate790(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate791(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate792(.a(G251), .O(gate236inter7));
  inv1  gate793(.a(G727), .O(gate236inter8));
  nand2 gate794(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate795(.a(s_35), .b(gate236inter3), .O(gate236inter10));
  nor2  gate796(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate797(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate798(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );

  xor2  gate631(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate632(.a(gate239inter0), .b(s_12), .O(gate239inter1));
  and2  gate633(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate634(.a(s_12), .O(gate239inter3));
  inv1  gate635(.a(s_13), .O(gate239inter4));
  nand2 gate636(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate637(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate638(.a(G260), .O(gate239inter7));
  inv1  gate639(.a(G712), .O(gate239inter8));
  nand2 gate640(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate641(.a(s_13), .b(gate239inter3), .O(gate239inter10));
  nor2  gate642(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate643(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate644(.a(gate239inter12), .b(gate239inter1), .O(G748));
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate1695(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate1696(.a(gate245inter0), .b(s_164), .O(gate245inter1));
  and2  gate1697(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate1698(.a(s_164), .O(gate245inter3));
  inv1  gate1699(.a(s_165), .O(gate245inter4));
  nand2 gate1700(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate1701(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate1702(.a(G248), .O(gate245inter7));
  inv1  gate1703(.a(G736), .O(gate245inter8));
  nand2 gate1704(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate1705(.a(s_165), .b(gate245inter3), .O(gate245inter10));
  nor2  gate1706(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate1707(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate1708(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate1499(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate1500(.a(gate250inter0), .b(s_136), .O(gate250inter1));
  and2  gate1501(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate1502(.a(s_136), .O(gate250inter3));
  inv1  gate1503(.a(s_137), .O(gate250inter4));
  nand2 gate1504(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate1505(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate1506(.a(G706), .O(gate250inter7));
  inv1  gate1507(.a(G742), .O(gate250inter8));
  nand2 gate1508(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate1509(.a(s_137), .b(gate250inter3), .O(gate250inter10));
  nor2  gate1510(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate1511(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate1512(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate1359(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate1360(.a(gate255inter0), .b(s_116), .O(gate255inter1));
  and2  gate1361(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate1362(.a(s_116), .O(gate255inter3));
  inv1  gate1363(.a(s_117), .O(gate255inter4));
  nand2 gate1364(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate1365(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate1366(.a(G263), .O(gate255inter7));
  inv1  gate1367(.a(G751), .O(gate255inter8));
  nand2 gate1368(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate1369(.a(s_117), .b(gate255inter3), .O(gate255inter10));
  nor2  gate1370(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate1371(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate1372(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );

  xor2  gate575(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate576(.a(gate264inter0), .b(s_4), .O(gate264inter1));
  and2  gate577(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate578(.a(s_4), .O(gate264inter3));
  inv1  gate579(.a(s_5), .O(gate264inter4));
  nand2 gate580(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate581(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate582(.a(G768), .O(gate264inter7));
  inv1  gate583(.a(G769), .O(gate264inter8));
  nand2 gate584(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate585(.a(s_5), .b(gate264inter3), .O(gate264inter10));
  nor2  gate586(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate587(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate588(.a(gate264inter12), .b(gate264inter1), .O(G791));

  xor2  gate1443(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate1444(.a(gate265inter0), .b(s_128), .O(gate265inter1));
  and2  gate1445(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate1446(.a(s_128), .O(gate265inter3));
  inv1  gate1447(.a(s_129), .O(gate265inter4));
  nand2 gate1448(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate1449(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate1450(.a(G642), .O(gate265inter7));
  inv1  gate1451(.a(G770), .O(gate265inter8));
  nand2 gate1452(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate1453(.a(s_129), .b(gate265inter3), .O(gate265inter10));
  nor2  gate1454(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate1455(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate1456(.a(gate265inter12), .b(gate265inter1), .O(G794));

  xor2  gate1303(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate1304(.a(gate266inter0), .b(s_108), .O(gate266inter1));
  and2  gate1305(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate1306(.a(s_108), .O(gate266inter3));
  inv1  gate1307(.a(s_109), .O(gate266inter4));
  nand2 gate1308(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate1309(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate1310(.a(G645), .O(gate266inter7));
  inv1  gate1311(.a(G773), .O(gate266inter8));
  nand2 gate1312(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate1313(.a(s_109), .b(gate266inter3), .O(gate266inter10));
  nor2  gate1314(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate1315(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate1316(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate1555(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate1556(.a(gate269inter0), .b(s_144), .O(gate269inter1));
  and2  gate1557(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate1558(.a(s_144), .O(gate269inter3));
  inv1  gate1559(.a(s_145), .O(gate269inter4));
  nand2 gate1560(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate1561(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate1562(.a(G654), .O(gate269inter7));
  inv1  gate1563(.a(G782), .O(gate269inter8));
  nand2 gate1564(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate1565(.a(s_145), .b(gate269inter3), .O(gate269inter10));
  nor2  gate1566(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate1567(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate1568(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );

  xor2  gate1037(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate1038(.a(gate273inter0), .b(s_70), .O(gate273inter1));
  and2  gate1039(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate1040(.a(s_70), .O(gate273inter3));
  inv1  gate1041(.a(s_71), .O(gate273inter4));
  nand2 gate1042(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate1043(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate1044(.a(G642), .O(gate273inter7));
  inv1  gate1045(.a(G794), .O(gate273inter8));
  nand2 gate1046(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate1047(.a(s_71), .b(gate273inter3), .O(gate273inter10));
  nor2  gate1048(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate1049(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate1050(.a(gate273inter12), .b(gate273inter1), .O(G818));
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate1261(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate1262(.a(gate276inter0), .b(s_102), .O(gate276inter1));
  and2  gate1263(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate1264(.a(s_102), .O(gate276inter3));
  inv1  gate1265(.a(s_103), .O(gate276inter4));
  nand2 gate1266(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate1267(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate1268(.a(G773), .O(gate276inter7));
  inv1  gate1269(.a(G797), .O(gate276inter8));
  nand2 gate1270(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate1271(.a(s_103), .b(gate276inter3), .O(gate276inter10));
  nor2  gate1272(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate1273(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate1274(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate799(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate800(.a(gate278inter0), .b(s_36), .O(gate278inter1));
  and2  gate801(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate802(.a(s_36), .O(gate278inter3));
  inv1  gate803(.a(s_37), .O(gate278inter4));
  nand2 gate804(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate805(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate806(.a(G776), .O(gate278inter7));
  inv1  gate807(.a(G800), .O(gate278inter8));
  nand2 gate808(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate809(.a(s_37), .b(gate278inter3), .O(gate278inter10));
  nor2  gate810(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate811(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate812(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate729(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate730(.a(gate286inter0), .b(s_26), .O(gate286inter1));
  and2  gate731(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate732(.a(s_26), .O(gate286inter3));
  inv1  gate733(.a(s_27), .O(gate286inter4));
  nand2 gate734(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate735(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate736(.a(G788), .O(gate286inter7));
  inv1  gate737(.a(G812), .O(gate286inter8));
  nand2 gate738(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate739(.a(s_27), .b(gate286inter3), .O(gate286inter10));
  nor2  gate740(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate741(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate742(.a(gate286inter12), .b(gate286inter1), .O(G831));
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate1205(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate1206(.a(gate291inter0), .b(s_94), .O(gate291inter1));
  and2  gate1207(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate1208(.a(s_94), .O(gate291inter3));
  inv1  gate1209(.a(s_95), .O(gate291inter4));
  nand2 gate1210(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate1211(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate1212(.a(G822), .O(gate291inter7));
  inv1  gate1213(.a(G823), .O(gate291inter8));
  nand2 gate1214(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate1215(.a(s_95), .b(gate291inter3), .O(gate291inter10));
  nor2  gate1216(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate1217(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate1218(.a(gate291inter12), .b(gate291inter1), .O(G860));

  xor2  gate1639(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate1640(.a(gate292inter0), .b(s_156), .O(gate292inter1));
  and2  gate1641(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate1642(.a(s_156), .O(gate292inter3));
  inv1  gate1643(.a(s_157), .O(gate292inter4));
  nand2 gate1644(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate1645(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate1646(.a(G824), .O(gate292inter7));
  inv1  gate1647(.a(G825), .O(gate292inter8));
  nand2 gate1648(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate1649(.a(s_157), .b(gate292inter3), .O(gate292inter10));
  nor2  gate1650(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate1651(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate1652(.a(gate292inter12), .b(gate292inter1), .O(G873));

  xor2  gate1149(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate1150(.a(gate293inter0), .b(s_86), .O(gate293inter1));
  and2  gate1151(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate1152(.a(s_86), .O(gate293inter3));
  inv1  gate1153(.a(s_87), .O(gate293inter4));
  nand2 gate1154(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate1155(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate1156(.a(G828), .O(gate293inter7));
  inv1  gate1157(.a(G829), .O(gate293inter8));
  nand2 gate1158(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate1159(.a(s_87), .b(gate293inter3), .O(gate293inter10));
  nor2  gate1160(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate1161(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate1162(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );

  xor2  gate1275(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate1276(.a(gate392inter0), .b(s_104), .O(gate392inter1));
  and2  gate1277(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate1278(.a(s_104), .O(gate392inter3));
  inv1  gate1279(.a(s_105), .O(gate392inter4));
  nand2 gate1280(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate1281(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate1282(.a(G6), .O(gate392inter7));
  inv1  gate1283(.a(G1051), .O(gate392inter8));
  nand2 gate1284(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate1285(.a(s_105), .b(gate392inter3), .O(gate392inter10));
  nor2  gate1286(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate1287(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate1288(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );

  xor2  gate953(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate954(.a(gate405inter0), .b(s_58), .O(gate405inter1));
  and2  gate955(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate956(.a(s_58), .O(gate405inter3));
  inv1  gate957(.a(s_59), .O(gate405inter4));
  nand2 gate958(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate959(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate960(.a(G19), .O(gate405inter7));
  inv1  gate961(.a(G1090), .O(gate405inter8));
  nand2 gate962(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate963(.a(s_59), .b(gate405inter3), .O(gate405inter10));
  nor2  gate964(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate965(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate966(.a(gate405inter12), .b(gate405inter1), .O(G1186));

  xor2  gate1597(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate1598(.a(gate406inter0), .b(s_150), .O(gate406inter1));
  and2  gate1599(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate1600(.a(s_150), .O(gate406inter3));
  inv1  gate1601(.a(s_151), .O(gate406inter4));
  nand2 gate1602(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate1603(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate1604(.a(G20), .O(gate406inter7));
  inv1  gate1605(.a(G1093), .O(gate406inter8));
  nand2 gate1606(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate1607(.a(s_151), .b(gate406inter3), .O(gate406inter10));
  nor2  gate1608(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate1609(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate1610(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate1807(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate1808(.a(gate411inter0), .b(s_180), .O(gate411inter1));
  and2  gate1809(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate1810(.a(s_180), .O(gate411inter3));
  inv1  gate1811(.a(s_181), .O(gate411inter4));
  nand2 gate1812(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate1813(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate1814(.a(G25), .O(gate411inter7));
  inv1  gate1815(.a(G1108), .O(gate411inter8));
  nand2 gate1816(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate1817(.a(s_181), .b(gate411inter3), .O(gate411inter10));
  nor2  gate1818(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate1819(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate1820(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );

  xor2  gate827(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate828(.a(gate414inter0), .b(s_40), .O(gate414inter1));
  and2  gate829(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate830(.a(s_40), .O(gate414inter3));
  inv1  gate831(.a(s_41), .O(gate414inter4));
  nand2 gate832(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate833(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate834(.a(G28), .O(gate414inter7));
  inv1  gate835(.a(G1117), .O(gate414inter8));
  nand2 gate836(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate837(.a(s_41), .b(gate414inter3), .O(gate414inter10));
  nor2  gate838(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate839(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate840(.a(gate414inter12), .b(gate414inter1), .O(G1213));
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );

  xor2  gate1289(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate1290(.a(gate418inter0), .b(s_106), .O(gate418inter1));
  and2  gate1291(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate1292(.a(s_106), .O(gate418inter3));
  inv1  gate1293(.a(s_107), .O(gate418inter4));
  nand2 gate1294(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate1295(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate1296(.a(G32), .O(gate418inter7));
  inv1  gate1297(.a(G1129), .O(gate418inter8));
  nand2 gate1298(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate1299(.a(s_107), .b(gate418inter3), .O(gate418inter10));
  nor2  gate1300(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate1301(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate1302(.a(gate418inter12), .b(gate418inter1), .O(G1225));

  xor2  gate1681(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate1682(.a(gate419inter0), .b(s_162), .O(gate419inter1));
  and2  gate1683(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate1684(.a(s_162), .O(gate419inter3));
  inv1  gate1685(.a(s_163), .O(gate419inter4));
  nand2 gate1686(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate1687(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate1688(.a(G1), .O(gate419inter7));
  inv1  gate1689(.a(G1132), .O(gate419inter8));
  nand2 gate1690(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate1691(.a(s_163), .b(gate419inter3), .O(gate419inter10));
  nor2  gate1692(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate1693(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate1694(.a(gate419inter12), .b(gate419inter1), .O(G1228));
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate603(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate604(.a(gate422inter0), .b(s_8), .O(gate422inter1));
  and2  gate605(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate606(.a(s_8), .O(gate422inter3));
  inv1  gate607(.a(s_9), .O(gate422inter4));
  nand2 gate608(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate609(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate610(.a(G1039), .O(gate422inter7));
  inv1  gate611(.a(G1135), .O(gate422inter8));
  nand2 gate612(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate613(.a(s_9), .b(gate422inter3), .O(gate422inter10));
  nor2  gate614(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate615(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate616(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate1709(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate1710(.a(gate430inter0), .b(s_166), .O(gate430inter1));
  and2  gate1711(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate1712(.a(s_166), .O(gate430inter3));
  inv1  gate1713(.a(s_167), .O(gate430inter4));
  nand2 gate1714(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate1715(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate1716(.a(G1051), .O(gate430inter7));
  inv1  gate1717(.a(G1147), .O(gate430inter8));
  nand2 gate1718(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate1719(.a(s_167), .b(gate430inter3), .O(gate430inter10));
  nor2  gate1720(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate1721(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate1722(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );

  xor2  gate687(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate688(.a(gate436inter0), .b(s_20), .O(gate436inter1));
  and2  gate689(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate690(.a(s_20), .O(gate436inter3));
  inv1  gate691(.a(s_21), .O(gate436inter4));
  nand2 gate692(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate693(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate694(.a(G1060), .O(gate436inter7));
  inv1  gate695(.a(G1156), .O(gate436inter8));
  nand2 gate696(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate697(.a(s_21), .b(gate436inter3), .O(gate436inter10));
  nor2  gate698(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate699(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate700(.a(gate436inter12), .b(gate436inter1), .O(G1245));
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate1373(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate1374(.a(gate439inter0), .b(s_118), .O(gate439inter1));
  and2  gate1375(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate1376(.a(s_118), .O(gate439inter3));
  inv1  gate1377(.a(s_119), .O(gate439inter4));
  nand2 gate1378(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate1379(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate1380(.a(G11), .O(gate439inter7));
  inv1  gate1381(.a(G1162), .O(gate439inter8));
  nand2 gate1382(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate1383(.a(s_119), .b(gate439inter3), .O(gate439inter10));
  nor2  gate1384(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate1385(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate1386(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate1107(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate1108(.a(gate448inter0), .b(s_80), .O(gate448inter1));
  and2  gate1109(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate1110(.a(s_80), .O(gate448inter3));
  inv1  gate1111(.a(s_81), .O(gate448inter4));
  nand2 gate1112(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate1113(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate1114(.a(G1078), .O(gate448inter7));
  inv1  gate1115(.a(G1174), .O(gate448inter8));
  nand2 gate1116(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate1117(.a(s_81), .b(gate448inter3), .O(gate448inter10));
  nor2  gate1118(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate1119(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate1120(.a(gate448inter12), .b(gate448inter1), .O(G1257));
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );

  xor2  gate939(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate940(.a(gate454inter0), .b(s_56), .O(gate454inter1));
  and2  gate941(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate942(.a(s_56), .O(gate454inter3));
  inv1  gate943(.a(s_57), .O(gate454inter4));
  nand2 gate944(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate945(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate946(.a(G1087), .O(gate454inter7));
  inv1  gate947(.a(G1183), .O(gate454inter8));
  nand2 gate948(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate949(.a(s_57), .b(gate454inter3), .O(gate454inter10));
  nor2  gate950(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate951(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate952(.a(gate454inter12), .b(gate454inter1), .O(G1263));
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate1527(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate1528(.a(gate457inter0), .b(s_140), .O(gate457inter1));
  and2  gate1529(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate1530(.a(s_140), .O(gate457inter3));
  inv1  gate1531(.a(s_141), .O(gate457inter4));
  nand2 gate1532(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate1533(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate1534(.a(G20), .O(gate457inter7));
  inv1  gate1535(.a(G1189), .O(gate457inter8));
  nand2 gate1536(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate1537(.a(s_141), .b(gate457inter3), .O(gate457inter10));
  nor2  gate1538(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate1539(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate1540(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate1611(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate1612(.a(gate460inter0), .b(s_152), .O(gate460inter1));
  and2  gate1613(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate1614(.a(s_152), .O(gate460inter3));
  inv1  gate1615(.a(s_153), .O(gate460inter4));
  nand2 gate1616(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate1617(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate1618(.a(G1096), .O(gate460inter7));
  inv1  gate1619(.a(G1192), .O(gate460inter8));
  nand2 gate1620(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate1621(.a(s_153), .b(gate460inter3), .O(gate460inter10));
  nor2  gate1622(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate1623(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate1624(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate1121(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate1122(.a(gate464inter0), .b(s_82), .O(gate464inter1));
  and2  gate1123(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate1124(.a(s_82), .O(gate464inter3));
  inv1  gate1125(.a(s_83), .O(gate464inter4));
  nand2 gate1126(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate1127(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate1128(.a(G1102), .O(gate464inter7));
  inv1  gate1129(.a(G1198), .O(gate464inter8));
  nand2 gate1130(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate1131(.a(s_83), .b(gate464inter3), .O(gate464inter10));
  nor2  gate1132(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate1133(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate1134(.a(gate464inter12), .b(gate464inter1), .O(G1273));

  xor2  gate1737(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate1738(.a(gate465inter0), .b(s_170), .O(gate465inter1));
  and2  gate1739(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate1740(.a(s_170), .O(gate465inter3));
  inv1  gate1741(.a(s_171), .O(gate465inter4));
  nand2 gate1742(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate1743(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate1744(.a(G24), .O(gate465inter7));
  inv1  gate1745(.a(G1201), .O(gate465inter8));
  nand2 gate1746(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate1747(.a(s_171), .b(gate465inter3), .O(gate465inter10));
  nor2  gate1748(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate1749(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate1750(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate1667(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate1668(.a(gate467inter0), .b(s_160), .O(gate467inter1));
  and2  gate1669(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate1670(.a(s_160), .O(gate467inter3));
  inv1  gate1671(.a(s_161), .O(gate467inter4));
  nand2 gate1672(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate1673(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate1674(.a(G25), .O(gate467inter7));
  inv1  gate1675(.a(G1204), .O(gate467inter8));
  nand2 gate1676(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate1677(.a(s_161), .b(gate467inter3), .O(gate467inter10));
  nor2  gate1678(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate1679(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate1680(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );

  xor2  gate1009(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate1010(.a(gate470inter0), .b(s_66), .O(gate470inter1));
  and2  gate1011(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate1012(.a(s_66), .O(gate470inter3));
  inv1  gate1013(.a(s_67), .O(gate470inter4));
  nand2 gate1014(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate1015(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate1016(.a(G1111), .O(gate470inter7));
  inv1  gate1017(.a(G1207), .O(gate470inter8));
  nand2 gate1018(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate1019(.a(s_67), .b(gate470inter3), .O(gate470inter10));
  nor2  gate1020(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate1021(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate1022(.a(gate470inter12), .b(gate470inter1), .O(G1279));
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );

  xor2  gate1723(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate1724(.a(gate473inter0), .b(s_168), .O(gate473inter1));
  and2  gate1725(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate1726(.a(s_168), .O(gate473inter3));
  inv1  gate1727(.a(s_169), .O(gate473inter4));
  nand2 gate1728(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate1729(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate1730(.a(G28), .O(gate473inter7));
  inv1  gate1731(.a(G1213), .O(gate473inter8));
  nand2 gate1732(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate1733(.a(s_169), .b(gate473inter3), .O(gate473inter10));
  nor2  gate1734(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate1735(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate1736(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate1331(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate1332(.a(gate476inter0), .b(s_112), .O(gate476inter1));
  and2  gate1333(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate1334(.a(s_112), .O(gate476inter3));
  inv1  gate1335(.a(s_113), .O(gate476inter4));
  nand2 gate1336(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate1337(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate1338(.a(G1120), .O(gate476inter7));
  inv1  gate1339(.a(G1216), .O(gate476inter8));
  nand2 gate1340(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate1341(.a(s_113), .b(gate476inter3), .O(gate476inter10));
  nor2  gate1342(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate1343(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate1344(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate1541(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate1542(.a(gate481inter0), .b(s_142), .O(gate481inter1));
  and2  gate1543(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate1544(.a(s_142), .O(gate481inter3));
  inv1  gate1545(.a(s_143), .O(gate481inter4));
  nand2 gate1546(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate1547(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate1548(.a(G32), .O(gate481inter7));
  inv1  gate1549(.a(G1225), .O(gate481inter8));
  nand2 gate1550(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate1551(.a(s_143), .b(gate481inter3), .O(gate481inter10));
  nor2  gate1552(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate1553(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate1554(.a(gate481inter12), .b(gate481inter1), .O(G1290));
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate925(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate926(.a(gate486inter0), .b(s_54), .O(gate486inter1));
  and2  gate927(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate928(.a(s_54), .O(gate486inter3));
  inv1  gate929(.a(s_55), .O(gate486inter4));
  nand2 gate930(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate931(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate932(.a(G1234), .O(gate486inter7));
  inv1  gate933(.a(G1235), .O(gate486inter8));
  nand2 gate934(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate935(.a(s_55), .b(gate486inter3), .O(gate486inter10));
  nor2  gate936(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate937(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate938(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate1569(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate1570(.a(gate489inter0), .b(s_146), .O(gate489inter1));
  and2  gate1571(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate1572(.a(s_146), .O(gate489inter3));
  inv1  gate1573(.a(s_147), .O(gate489inter4));
  nand2 gate1574(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate1575(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate1576(.a(G1240), .O(gate489inter7));
  inv1  gate1577(.a(G1241), .O(gate489inter8));
  nand2 gate1578(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate1579(.a(s_147), .b(gate489inter3), .O(gate489inter10));
  nor2  gate1580(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate1581(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate1582(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate1415(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate1416(.a(gate493inter0), .b(s_124), .O(gate493inter1));
  and2  gate1417(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate1418(.a(s_124), .O(gate493inter3));
  inv1  gate1419(.a(s_125), .O(gate493inter4));
  nand2 gate1420(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate1421(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate1422(.a(G1248), .O(gate493inter7));
  inv1  gate1423(.a(G1249), .O(gate493inter8));
  nand2 gate1424(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate1425(.a(s_125), .b(gate493inter3), .O(gate493inter10));
  nor2  gate1426(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate1427(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate1428(.a(gate493inter12), .b(gate493inter1), .O(G1302));
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate1471(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate1472(.a(gate503inter0), .b(s_132), .O(gate503inter1));
  and2  gate1473(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate1474(.a(s_132), .O(gate503inter3));
  inv1  gate1475(.a(s_133), .O(gate503inter4));
  nand2 gate1476(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate1477(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate1478(.a(G1268), .O(gate503inter7));
  inv1  gate1479(.a(G1269), .O(gate503inter8));
  nand2 gate1480(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate1481(.a(s_133), .b(gate503inter3), .O(gate503inter10));
  nor2  gate1482(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate1483(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate1484(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate855(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate856(.a(gate511inter0), .b(s_44), .O(gate511inter1));
  and2  gate857(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate858(.a(s_44), .O(gate511inter3));
  inv1  gate859(.a(s_45), .O(gate511inter4));
  nand2 gate860(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate861(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate862(.a(G1284), .O(gate511inter7));
  inv1  gate863(.a(G1285), .O(gate511inter8));
  nand2 gate864(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate865(.a(s_45), .b(gate511inter3), .O(gate511inter10));
  nor2  gate866(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate867(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate868(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );

  xor2  gate813(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate814(.a(gate513inter0), .b(s_38), .O(gate513inter1));
  and2  gate815(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate816(.a(s_38), .O(gate513inter3));
  inv1  gate817(.a(s_39), .O(gate513inter4));
  nand2 gate818(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate819(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate820(.a(G1288), .O(gate513inter7));
  inv1  gate821(.a(G1289), .O(gate513inter8));
  nand2 gate822(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate823(.a(s_39), .b(gate513inter3), .O(gate513inter10));
  nor2  gate824(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate825(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate826(.a(gate513inter12), .b(gate513inter1), .O(G1322));
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule