module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281, s_282, s_283, s_284, s_285, s_286, s_287, s_288, s_289, s_290, s_291, s_292, s_293, s_294, s_295, s_296, s_297, s_298, s_299, s_300, s_301, s_302, s_303, s_304, s_305, s_306, s_307, s_308, s_309, s_310, s_311, s_312, s_313, s_314, s_315, s_316, s_317, s_318, s_319, s_320, s_321;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate2703(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate2704(.a(gate9inter0), .b(s_308), .O(gate9inter1));
  and2  gate2705(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate2706(.a(s_308), .O(gate9inter3));
  inv1  gate2707(.a(s_309), .O(gate9inter4));
  nand2 gate2708(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate2709(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate2710(.a(G1), .O(gate9inter7));
  inv1  gate2711(.a(G2), .O(gate9inter8));
  nand2 gate2712(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate2713(.a(s_309), .b(gate9inter3), .O(gate9inter10));
  nor2  gate2714(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate2715(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate2716(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate1877(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate1878(.a(gate16inter0), .b(s_190), .O(gate16inter1));
  and2  gate1879(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate1880(.a(s_190), .O(gate16inter3));
  inv1  gate1881(.a(s_191), .O(gate16inter4));
  nand2 gate1882(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate1883(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate1884(.a(G15), .O(gate16inter7));
  inv1  gate1885(.a(G16), .O(gate16inter8));
  nand2 gate1886(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate1887(.a(s_191), .b(gate16inter3), .O(gate16inter10));
  nor2  gate1888(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate1889(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate1890(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate1303(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate1304(.a(gate18inter0), .b(s_108), .O(gate18inter1));
  and2  gate1305(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate1306(.a(s_108), .O(gate18inter3));
  inv1  gate1307(.a(s_109), .O(gate18inter4));
  nand2 gate1308(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate1309(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate1310(.a(G19), .O(gate18inter7));
  inv1  gate1311(.a(G20), .O(gate18inter8));
  nand2 gate1312(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate1313(.a(s_109), .b(gate18inter3), .O(gate18inter10));
  nor2  gate1314(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate1315(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate1316(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate1499(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate1500(.a(gate20inter0), .b(s_136), .O(gate20inter1));
  and2  gate1501(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate1502(.a(s_136), .O(gate20inter3));
  inv1  gate1503(.a(s_137), .O(gate20inter4));
  nand2 gate1504(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate1505(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate1506(.a(G23), .O(gate20inter7));
  inv1  gate1507(.a(G24), .O(gate20inter8));
  nand2 gate1508(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate1509(.a(s_137), .b(gate20inter3), .O(gate20inter10));
  nor2  gate1510(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate1511(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate1512(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate2479(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate2480(.a(gate23inter0), .b(s_276), .O(gate23inter1));
  and2  gate2481(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate2482(.a(s_276), .O(gate23inter3));
  inv1  gate2483(.a(s_277), .O(gate23inter4));
  nand2 gate2484(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate2485(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate2486(.a(G29), .O(gate23inter7));
  inv1  gate2487(.a(G30), .O(gate23inter8));
  nand2 gate2488(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate2489(.a(s_277), .b(gate23inter3), .O(gate23inter10));
  nor2  gate2490(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate2491(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate2492(.a(gate23inter12), .b(gate23inter1), .O(G308));

  xor2  gate1779(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate1780(.a(gate24inter0), .b(s_176), .O(gate24inter1));
  and2  gate1781(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate1782(.a(s_176), .O(gate24inter3));
  inv1  gate1783(.a(s_177), .O(gate24inter4));
  nand2 gate1784(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate1785(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate1786(.a(G31), .O(gate24inter7));
  inv1  gate1787(.a(G32), .O(gate24inter8));
  nand2 gate1788(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate1789(.a(s_177), .b(gate24inter3), .O(gate24inter10));
  nor2  gate1790(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate1791(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate1792(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate561(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate562(.a(gate26inter0), .b(s_2), .O(gate26inter1));
  and2  gate563(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate564(.a(s_2), .O(gate26inter3));
  inv1  gate565(.a(s_3), .O(gate26inter4));
  nand2 gate566(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate567(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate568(.a(G9), .O(gate26inter7));
  inv1  gate569(.a(G13), .O(gate26inter8));
  nand2 gate570(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate571(.a(s_3), .b(gate26inter3), .O(gate26inter10));
  nor2  gate572(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate573(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate574(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate673(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate674(.a(gate31inter0), .b(s_18), .O(gate31inter1));
  and2  gate675(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate676(.a(s_18), .O(gate31inter3));
  inv1  gate677(.a(s_19), .O(gate31inter4));
  nand2 gate678(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate679(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate680(.a(G4), .O(gate31inter7));
  inv1  gate681(.a(G8), .O(gate31inter8));
  nand2 gate682(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate683(.a(s_19), .b(gate31inter3), .O(gate31inter10));
  nor2  gate684(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate685(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate686(.a(gate31inter12), .b(gate31inter1), .O(G332));

  xor2  gate1457(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate1458(.a(gate32inter0), .b(s_130), .O(gate32inter1));
  and2  gate1459(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate1460(.a(s_130), .O(gate32inter3));
  inv1  gate1461(.a(s_131), .O(gate32inter4));
  nand2 gate1462(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate1463(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate1464(.a(G12), .O(gate32inter7));
  inv1  gate1465(.a(G16), .O(gate32inter8));
  nand2 gate1466(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate1467(.a(s_131), .b(gate32inter3), .O(gate32inter10));
  nor2  gate1468(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate1469(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate1470(.a(gate32inter12), .b(gate32inter1), .O(G335));
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate1653(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate1654(.a(gate34inter0), .b(s_158), .O(gate34inter1));
  and2  gate1655(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate1656(.a(s_158), .O(gate34inter3));
  inv1  gate1657(.a(s_159), .O(gate34inter4));
  nand2 gate1658(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate1659(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate1660(.a(G25), .O(gate34inter7));
  inv1  gate1661(.a(G29), .O(gate34inter8));
  nand2 gate1662(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate1663(.a(s_159), .b(gate34inter3), .O(gate34inter10));
  nor2  gate1664(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate1665(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate1666(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate1317(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1318(.a(gate36inter0), .b(s_110), .O(gate36inter1));
  and2  gate1319(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1320(.a(s_110), .O(gate36inter3));
  inv1  gate1321(.a(s_111), .O(gate36inter4));
  nand2 gate1322(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1323(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1324(.a(G26), .O(gate36inter7));
  inv1  gate1325(.a(G30), .O(gate36inter8));
  nand2 gate1326(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1327(.a(s_111), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1328(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1329(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1330(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate771(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate772(.a(gate38inter0), .b(s_32), .O(gate38inter1));
  and2  gate773(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate774(.a(s_32), .O(gate38inter3));
  inv1  gate775(.a(s_33), .O(gate38inter4));
  nand2 gate776(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate777(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate778(.a(G27), .O(gate38inter7));
  inv1  gate779(.a(G31), .O(gate38inter8));
  nand2 gate780(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate781(.a(s_33), .b(gate38inter3), .O(gate38inter10));
  nor2  gate782(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate783(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate784(.a(gate38inter12), .b(gate38inter1), .O(G353));
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate2199(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate2200(.a(gate41inter0), .b(s_236), .O(gate41inter1));
  and2  gate2201(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate2202(.a(s_236), .O(gate41inter3));
  inv1  gate2203(.a(s_237), .O(gate41inter4));
  nand2 gate2204(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate2205(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate2206(.a(G1), .O(gate41inter7));
  inv1  gate2207(.a(G266), .O(gate41inter8));
  nand2 gate2208(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate2209(.a(s_237), .b(gate41inter3), .O(gate41inter10));
  nor2  gate2210(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate2211(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate2212(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate2241(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate2242(.a(gate46inter0), .b(s_242), .O(gate46inter1));
  and2  gate2243(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate2244(.a(s_242), .O(gate46inter3));
  inv1  gate2245(.a(s_243), .O(gate46inter4));
  nand2 gate2246(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate2247(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate2248(.a(G6), .O(gate46inter7));
  inv1  gate2249(.a(G272), .O(gate46inter8));
  nand2 gate2250(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate2251(.a(s_243), .b(gate46inter3), .O(gate46inter10));
  nor2  gate2252(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate2253(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate2254(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );

  xor2  gate1219(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate1220(.a(gate50inter0), .b(s_96), .O(gate50inter1));
  and2  gate1221(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate1222(.a(s_96), .O(gate50inter3));
  inv1  gate1223(.a(s_97), .O(gate50inter4));
  nand2 gate1224(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate1225(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate1226(.a(G10), .O(gate50inter7));
  inv1  gate1227(.a(G278), .O(gate50inter8));
  nand2 gate1228(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate1229(.a(s_97), .b(gate50inter3), .O(gate50inter10));
  nor2  gate1230(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate1231(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate1232(.a(gate50inter12), .b(gate50inter1), .O(G371));
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );

  xor2  gate1947(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate1948(.a(gate53inter0), .b(s_200), .O(gate53inter1));
  and2  gate1949(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate1950(.a(s_200), .O(gate53inter3));
  inv1  gate1951(.a(s_201), .O(gate53inter4));
  nand2 gate1952(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate1953(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate1954(.a(G13), .O(gate53inter7));
  inv1  gate1955(.a(G284), .O(gate53inter8));
  nand2 gate1956(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate1957(.a(s_201), .b(gate53inter3), .O(gate53inter10));
  nor2  gate1958(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate1959(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate1960(.a(gate53inter12), .b(gate53inter1), .O(G374));

  xor2  gate2661(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate2662(.a(gate54inter0), .b(s_302), .O(gate54inter1));
  and2  gate2663(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate2664(.a(s_302), .O(gate54inter3));
  inv1  gate2665(.a(s_303), .O(gate54inter4));
  nand2 gate2666(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate2667(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate2668(.a(G14), .O(gate54inter7));
  inv1  gate2669(.a(G284), .O(gate54inter8));
  nand2 gate2670(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate2671(.a(s_303), .b(gate54inter3), .O(gate54inter10));
  nor2  gate2672(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate2673(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate2674(.a(gate54inter12), .b(gate54inter1), .O(G375));

  xor2  gate1919(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate1920(.a(gate55inter0), .b(s_196), .O(gate55inter1));
  and2  gate1921(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate1922(.a(s_196), .O(gate55inter3));
  inv1  gate1923(.a(s_197), .O(gate55inter4));
  nand2 gate1924(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate1925(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate1926(.a(G15), .O(gate55inter7));
  inv1  gate1927(.a(G287), .O(gate55inter8));
  nand2 gate1928(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate1929(.a(s_197), .b(gate55inter3), .O(gate55inter10));
  nor2  gate1930(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate1931(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate1932(.a(gate55inter12), .b(gate55inter1), .O(G376));

  xor2  gate1037(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate1038(.a(gate56inter0), .b(s_70), .O(gate56inter1));
  and2  gate1039(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate1040(.a(s_70), .O(gate56inter3));
  inv1  gate1041(.a(s_71), .O(gate56inter4));
  nand2 gate1042(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate1043(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate1044(.a(G16), .O(gate56inter7));
  inv1  gate1045(.a(G287), .O(gate56inter8));
  nand2 gate1046(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate1047(.a(s_71), .b(gate56inter3), .O(gate56inter10));
  nor2  gate1048(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate1049(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate1050(.a(gate56inter12), .b(gate56inter1), .O(G377));

  xor2  gate1121(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate1122(.a(gate57inter0), .b(s_82), .O(gate57inter1));
  and2  gate1123(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate1124(.a(s_82), .O(gate57inter3));
  inv1  gate1125(.a(s_83), .O(gate57inter4));
  nand2 gate1126(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate1127(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate1128(.a(G17), .O(gate57inter7));
  inv1  gate1129(.a(G290), .O(gate57inter8));
  nand2 gate1130(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate1131(.a(s_83), .b(gate57inter3), .O(gate57inter10));
  nor2  gate1132(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate1133(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate1134(.a(gate57inter12), .b(gate57inter1), .O(G378));
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate1737(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate1738(.a(gate59inter0), .b(s_170), .O(gate59inter1));
  and2  gate1739(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate1740(.a(s_170), .O(gate59inter3));
  inv1  gate1741(.a(s_171), .O(gate59inter4));
  nand2 gate1742(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate1743(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate1744(.a(G19), .O(gate59inter7));
  inv1  gate1745(.a(G293), .O(gate59inter8));
  nand2 gate1746(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate1747(.a(s_171), .b(gate59inter3), .O(gate59inter10));
  nor2  gate1748(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate1749(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate1750(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );

  xor2  gate2115(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate2116(.a(gate61inter0), .b(s_224), .O(gate61inter1));
  and2  gate2117(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate2118(.a(s_224), .O(gate61inter3));
  inv1  gate2119(.a(s_225), .O(gate61inter4));
  nand2 gate2120(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate2121(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate2122(.a(G21), .O(gate61inter7));
  inv1  gate2123(.a(G296), .O(gate61inter8));
  nand2 gate2124(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate2125(.a(s_225), .b(gate61inter3), .O(gate61inter10));
  nor2  gate2126(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate2127(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate2128(.a(gate61inter12), .b(gate61inter1), .O(G382));
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );

  xor2  gate2171(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate2172(.a(gate64inter0), .b(s_232), .O(gate64inter1));
  and2  gate2173(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate2174(.a(s_232), .O(gate64inter3));
  inv1  gate2175(.a(s_233), .O(gate64inter4));
  nand2 gate2176(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate2177(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate2178(.a(G24), .O(gate64inter7));
  inv1  gate2179(.a(G299), .O(gate64inter8));
  nand2 gate2180(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate2181(.a(s_233), .b(gate64inter3), .O(gate64inter10));
  nor2  gate2182(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate2183(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate2184(.a(gate64inter12), .b(gate64inter1), .O(G385));

  xor2  gate1583(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate1584(.a(gate65inter0), .b(s_148), .O(gate65inter1));
  and2  gate1585(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate1586(.a(s_148), .O(gate65inter3));
  inv1  gate1587(.a(s_149), .O(gate65inter4));
  nand2 gate1588(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate1589(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate1590(.a(G25), .O(gate65inter7));
  inv1  gate1591(.a(G302), .O(gate65inter8));
  nand2 gate1592(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate1593(.a(s_149), .b(gate65inter3), .O(gate65inter10));
  nor2  gate1594(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate1595(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate1596(.a(gate65inter12), .b(gate65inter1), .O(G386));

  xor2  gate1191(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate1192(.a(gate66inter0), .b(s_92), .O(gate66inter1));
  and2  gate1193(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate1194(.a(s_92), .O(gate66inter3));
  inv1  gate1195(.a(s_93), .O(gate66inter4));
  nand2 gate1196(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate1197(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate1198(.a(G26), .O(gate66inter7));
  inv1  gate1199(.a(G302), .O(gate66inter8));
  nand2 gate1200(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate1201(.a(s_93), .b(gate66inter3), .O(gate66inter10));
  nor2  gate1202(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate1203(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate1204(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );

  xor2  gate2367(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate2368(.a(gate68inter0), .b(s_260), .O(gate68inter1));
  and2  gate2369(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate2370(.a(s_260), .O(gate68inter3));
  inv1  gate2371(.a(s_261), .O(gate68inter4));
  nand2 gate2372(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate2373(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate2374(.a(G28), .O(gate68inter7));
  inv1  gate2375(.a(G305), .O(gate68inter8));
  nand2 gate2376(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate2377(.a(s_261), .b(gate68inter3), .O(gate68inter10));
  nor2  gate2378(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate2379(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate2380(.a(gate68inter12), .b(gate68inter1), .O(G389));

  xor2  gate1807(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate1808(.a(gate69inter0), .b(s_180), .O(gate69inter1));
  and2  gate1809(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate1810(.a(s_180), .O(gate69inter3));
  inv1  gate1811(.a(s_181), .O(gate69inter4));
  nand2 gate1812(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate1813(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate1814(.a(G29), .O(gate69inter7));
  inv1  gate1815(.a(G308), .O(gate69inter8));
  nand2 gate1816(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate1817(.a(s_181), .b(gate69inter3), .O(gate69inter10));
  nor2  gate1818(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate1819(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate1820(.a(gate69inter12), .b(gate69inter1), .O(G390));
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate981(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate982(.a(gate71inter0), .b(s_62), .O(gate71inter1));
  and2  gate983(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate984(.a(s_62), .O(gate71inter3));
  inv1  gate985(.a(s_63), .O(gate71inter4));
  nand2 gate986(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate987(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate988(.a(G31), .O(gate71inter7));
  inv1  gate989(.a(G311), .O(gate71inter8));
  nand2 gate990(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate991(.a(s_63), .b(gate71inter3), .O(gate71inter10));
  nor2  gate992(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate993(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate994(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate1667(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate1668(.a(gate75inter0), .b(s_160), .O(gate75inter1));
  and2  gate1669(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate1670(.a(s_160), .O(gate75inter3));
  inv1  gate1671(.a(s_161), .O(gate75inter4));
  nand2 gate1672(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate1673(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate1674(.a(G9), .O(gate75inter7));
  inv1  gate1675(.a(G317), .O(gate75inter8));
  nand2 gate1676(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate1677(.a(s_161), .b(gate75inter3), .O(gate75inter10));
  nor2  gate1678(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate1679(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate1680(.a(gate75inter12), .b(gate75inter1), .O(G396));

  xor2  gate2759(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate2760(.a(gate76inter0), .b(s_316), .O(gate76inter1));
  and2  gate2761(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate2762(.a(s_316), .O(gate76inter3));
  inv1  gate2763(.a(s_317), .O(gate76inter4));
  nand2 gate2764(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate2765(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate2766(.a(G13), .O(gate76inter7));
  inv1  gate2767(.a(G317), .O(gate76inter8));
  nand2 gate2768(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate2769(.a(s_317), .b(gate76inter3), .O(gate76inter10));
  nor2  gate2770(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate2771(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate2772(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate911(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate912(.a(gate78inter0), .b(s_52), .O(gate78inter1));
  and2  gate913(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate914(.a(s_52), .O(gate78inter3));
  inv1  gate915(.a(s_53), .O(gate78inter4));
  nand2 gate916(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate917(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate918(.a(G6), .O(gate78inter7));
  inv1  gate919(.a(G320), .O(gate78inter8));
  nand2 gate920(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate921(.a(s_53), .b(gate78inter3), .O(gate78inter10));
  nor2  gate922(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate923(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate924(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate1331(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate1332(.a(gate82inter0), .b(s_112), .O(gate82inter1));
  and2  gate1333(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate1334(.a(s_112), .O(gate82inter3));
  inv1  gate1335(.a(s_113), .O(gate82inter4));
  nand2 gate1336(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate1337(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate1338(.a(G7), .O(gate82inter7));
  inv1  gate1339(.a(G326), .O(gate82inter8));
  nand2 gate1340(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate1341(.a(s_113), .b(gate82inter3), .O(gate82inter10));
  nor2  gate1342(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate1343(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate1344(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );

  xor2  gate2185(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate2186(.a(gate84inter0), .b(s_234), .O(gate84inter1));
  and2  gate2187(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate2188(.a(s_234), .O(gate84inter3));
  inv1  gate2189(.a(s_235), .O(gate84inter4));
  nand2 gate2190(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate2191(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate2192(.a(G15), .O(gate84inter7));
  inv1  gate2193(.a(G329), .O(gate84inter8));
  nand2 gate2194(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate2195(.a(s_235), .b(gate84inter3), .O(gate84inter10));
  nor2  gate2196(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate2197(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate2198(.a(gate84inter12), .b(gate84inter1), .O(G405));
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate2045(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate2046(.a(gate86inter0), .b(s_214), .O(gate86inter1));
  and2  gate2047(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate2048(.a(s_214), .O(gate86inter3));
  inv1  gate2049(.a(s_215), .O(gate86inter4));
  nand2 gate2050(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate2051(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate2052(.a(G8), .O(gate86inter7));
  inv1  gate2053(.a(G332), .O(gate86inter8));
  nand2 gate2054(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate2055(.a(s_215), .b(gate86inter3), .O(gate86inter10));
  nor2  gate2056(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate2057(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate2058(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate659(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate660(.a(gate88inter0), .b(s_16), .O(gate88inter1));
  and2  gate661(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate662(.a(s_16), .O(gate88inter3));
  inv1  gate663(.a(s_17), .O(gate88inter4));
  nand2 gate664(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate665(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate666(.a(G16), .O(gate88inter7));
  inv1  gate667(.a(G335), .O(gate88inter8));
  nand2 gate668(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate669(.a(s_17), .b(gate88inter3), .O(gate88inter10));
  nor2  gate670(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate671(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate672(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate1149(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate1150(.a(gate98inter0), .b(s_86), .O(gate98inter1));
  and2  gate1151(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate1152(.a(s_86), .O(gate98inter3));
  inv1  gate1153(.a(s_87), .O(gate98inter4));
  nand2 gate1154(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1155(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1156(.a(G23), .O(gate98inter7));
  inv1  gate1157(.a(G350), .O(gate98inter8));
  nand2 gate1158(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1159(.a(s_87), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1160(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1161(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1162(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate939(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate940(.a(gate100inter0), .b(s_56), .O(gate100inter1));
  and2  gate941(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate942(.a(s_56), .O(gate100inter3));
  inv1  gate943(.a(s_57), .O(gate100inter4));
  nand2 gate944(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate945(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate946(.a(G31), .O(gate100inter7));
  inv1  gate947(.a(G353), .O(gate100inter8));
  nand2 gate948(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate949(.a(s_57), .b(gate100inter3), .O(gate100inter10));
  nor2  gate950(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate951(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate952(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate2143(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate2144(.a(gate102inter0), .b(s_228), .O(gate102inter1));
  and2  gate2145(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate2146(.a(s_228), .O(gate102inter3));
  inv1  gate2147(.a(s_229), .O(gate102inter4));
  nand2 gate2148(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate2149(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate2150(.a(G24), .O(gate102inter7));
  inv1  gate2151(.a(G356), .O(gate102inter8));
  nand2 gate2152(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate2153(.a(s_229), .b(gate102inter3), .O(gate102inter10));
  nor2  gate2154(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate2155(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate2156(.a(gate102inter12), .b(gate102inter1), .O(G423));

  xor2  gate1275(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate1276(.a(gate103inter0), .b(s_104), .O(gate103inter1));
  and2  gate1277(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate1278(.a(s_104), .O(gate103inter3));
  inv1  gate1279(.a(s_105), .O(gate103inter4));
  nand2 gate1280(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate1281(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate1282(.a(G28), .O(gate103inter7));
  inv1  gate1283(.a(G359), .O(gate103inter8));
  nand2 gate1284(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate1285(.a(s_105), .b(gate103inter3), .O(gate103inter10));
  nor2  gate1286(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate1287(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate1288(.a(gate103inter12), .b(gate103inter1), .O(G424));

  xor2  gate1597(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate1598(.a(gate104inter0), .b(s_150), .O(gate104inter1));
  and2  gate1599(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate1600(.a(s_150), .O(gate104inter3));
  inv1  gate1601(.a(s_151), .O(gate104inter4));
  nand2 gate1602(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate1603(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate1604(.a(G32), .O(gate104inter7));
  inv1  gate1605(.a(G359), .O(gate104inter8));
  nand2 gate1606(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate1607(.a(s_151), .b(gate104inter3), .O(gate104inter10));
  nor2  gate1608(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate1609(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate1610(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate925(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate926(.a(gate106inter0), .b(s_54), .O(gate106inter1));
  and2  gate927(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate928(.a(s_54), .O(gate106inter3));
  inv1  gate929(.a(s_55), .O(gate106inter4));
  nand2 gate930(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate931(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate932(.a(G364), .O(gate106inter7));
  inv1  gate933(.a(G365), .O(gate106inter8));
  nand2 gate934(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate935(.a(s_55), .b(gate106inter3), .O(gate106inter10));
  nor2  gate936(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate937(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate938(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate1849(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate1850(.a(gate109inter0), .b(s_186), .O(gate109inter1));
  and2  gate1851(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate1852(.a(s_186), .O(gate109inter3));
  inv1  gate1853(.a(s_187), .O(gate109inter4));
  nand2 gate1854(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate1855(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate1856(.a(G370), .O(gate109inter7));
  inv1  gate1857(.a(G371), .O(gate109inter8));
  nand2 gate1858(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate1859(.a(s_187), .b(gate109inter3), .O(gate109inter10));
  nor2  gate1860(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate1861(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate1862(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );

  xor2  gate1345(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate1346(.a(gate111inter0), .b(s_114), .O(gate111inter1));
  and2  gate1347(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate1348(.a(s_114), .O(gate111inter3));
  inv1  gate1349(.a(s_115), .O(gate111inter4));
  nand2 gate1350(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate1351(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate1352(.a(G374), .O(gate111inter7));
  inv1  gate1353(.a(G375), .O(gate111inter8));
  nand2 gate1354(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate1355(.a(s_115), .b(gate111inter3), .O(gate111inter10));
  nor2  gate1356(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate1357(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate1358(.a(gate111inter12), .b(gate111inter1), .O(G444));
nand2 gate112( .a(G376), .b(G377), .O(G447) );

  xor2  gate1821(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate1822(.a(gate113inter0), .b(s_182), .O(gate113inter1));
  and2  gate1823(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate1824(.a(s_182), .O(gate113inter3));
  inv1  gate1825(.a(s_183), .O(gate113inter4));
  nand2 gate1826(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate1827(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate1828(.a(G378), .O(gate113inter7));
  inv1  gate1829(.a(G379), .O(gate113inter8));
  nand2 gate1830(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate1831(.a(s_183), .b(gate113inter3), .O(gate113inter10));
  nor2  gate1832(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate1833(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate1834(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate1247(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate1248(.a(gate115inter0), .b(s_100), .O(gate115inter1));
  and2  gate1249(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate1250(.a(s_100), .O(gate115inter3));
  inv1  gate1251(.a(s_101), .O(gate115inter4));
  nand2 gate1252(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate1253(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate1254(.a(G382), .O(gate115inter7));
  inv1  gate1255(.a(G383), .O(gate115inter8));
  nand2 gate1256(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate1257(.a(s_101), .b(gate115inter3), .O(gate115inter10));
  nor2  gate1258(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate1259(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate1260(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate2353(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate2354(.a(gate119inter0), .b(s_258), .O(gate119inter1));
  and2  gate2355(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate2356(.a(s_258), .O(gate119inter3));
  inv1  gate2357(.a(s_259), .O(gate119inter4));
  nand2 gate2358(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate2359(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate2360(.a(G390), .O(gate119inter7));
  inv1  gate2361(.a(G391), .O(gate119inter8));
  nand2 gate2362(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate2363(.a(s_259), .b(gate119inter3), .O(gate119inter10));
  nor2  gate2364(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate2365(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate2366(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate1905(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate1906(.a(gate121inter0), .b(s_194), .O(gate121inter1));
  and2  gate1907(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate1908(.a(s_194), .O(gate121inter3));
  inv1  gate1909(.a(s_195), .O(gate121inter4));
  nand2 gate1910(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate1911(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate1912(.a(G394), .O(gate121inter7));
  inv1  gate1913(.a(G395), .O(gate121inter8));
  nand2 gate1914(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate1915(.a(s_195), .b(gate121inter3), .O(gate121inter10));
  nor2  gate1916(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate1917(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate1918(.a(gate121inter12), .b(gate121inter1), .O(G474));

  xor2  gate1289(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate1290(.a(gate122inter0), .b(s_106), .O(gate122inter1));
  and2  gate1291(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate1292(.a(s_106), .O(gate122inter3));
  inv1  gate1293(.a(s_107), .O(gate122inter4));
  nand2 gate1294(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate1295(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate1296(.a(G396), .O(gate122inter7));
  inv1  gate1297(.a(G397), .O(gate122inter8));
  nand2 gate1298(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate1299(.a(s_107), .b(gate122inter3), .O(gate122inter10));
  nor2  gate1300(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate1301(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate1302(.a(gate122inter12), .b(gate122inter1), .O(G477));
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate1093(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate1094(.a(gate126inter0), .b(s_78), .O(gate126inter1));
  and2  gate1095(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate1096(.a(s_78), .O(gate126inter3));
  inv1  gate1097(.a(s_79), .O(gate126inter4));
  nand2 gate1098(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate1099(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate1100(.a(G404), .O(gate126inter7));
  inv1  gate1101(.a(G405), .O(gate126inter8));
  nand2 gate1102(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate1103(.a(s_79), .b(gate126inter3), .O(gate126inter10));
  nor2  gate1104(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate1105(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate1106(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate2521(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate2522(.a(gate128inter0), .b(s_282), .O(gate128inter1));
  and2  gate2523(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate2524(.a(s_282), .O(gate128inter3));
  inv1  gate2525(.a(s_283), .O(gate128inter4));
  nand2 gate2526(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate2527(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate2528(.a(G408), .O(gate128inter7));
  inv1  gate2529(.a(G409), .O(gate128inter8));
  nand2 gate2530(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate2531(.a(s_283), .b(gate128inter3), .O(gate128inter10));
  nor2  gate2532(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate2533(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate2534(.a(gate128inter12), .b(gate128inter1), .O(G495));

  xor2  gate1933(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate1934(.a(gate129inter0), .b(s_198), .O(gate129inter1));
  and2  gate1935(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate1936(.a(s_198), .O(gate129inter3));
  inv1  gate1937(.a(s_199), .O(gate129inter4));
  nand2 gate1938(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate1939(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate1940(.a(G410), .O(gate129inter7));
  inv1  gate1941(.a(G411), .O(gate129inter8));
  nand2 gate1942(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate1943(.a(s_199), .b(gate129inter3), .O(gate129inter10));
  nor2  gate1944(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate1945(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate1946(.a(gate129inter12), .b(gate129inter1), .O(G498));
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate1555(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate1556(.a(gate132inter0), .b(s_144), .O(gate132inter1));
  and2  gate1557(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate1558(.a(s_144), .O(gate132inter3));
  inv1  gate1559(.a(s_145), .O(gate132inter4));
  nand2 gate1560(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate1561(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate1562(.a(G416), .O(gate132inter7));
  inv1  gate1563(.a(G417), .O(gate132inter8));
  nand2 gate1564(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate1565(.a(s_145), .b(gate132inter3), .O(gate132inter10));
  nor2  gate1566(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate1567(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate1568(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate2731(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate2732(.a(gate136inter0), .b(s_312), .O(gate136inter1));
  and2  gate2733(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate2734(.a(s_312), .O(gate136inter3));
  inv1  gate2735(.a(s_313), .O(gate136inter4));
  nand2 gate2736(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate2737(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate2738(.a(G424), .O(gate136inter7));
  inv1  gate2739(.a(G425), .O(gate136inter8));
  nand2 gate2740(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate2741(.a(s_313), .b(gate136inter3), .O(gate136inter10));
  nor2  gate2742(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate2743(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate2744(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate1023(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate1024(.a(gate141inter0), .b(s_68), .O(gate141inter1));
  and2  gate1025(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate1026(.a(s_68), .O(gate141inter3));
  inv1  gate1027(.a(s_69), .O(gate141inter4));
  nand2 gate1028(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate1029(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate1030(.a(G450), .O(gate141inter7));
  inv1  gate1031(.a(G453), .O(gate141inter8));
  nand2 gate1032(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate1033(.a(s_69), .b(gate141inter3), .O(gate141inter10));
  nor2  gate1034(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate1035(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate1036(.a(gate141inter12), .b(gate141inter1), .O(G534));

  xor2  gate2535(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate2536(.a(gate142inter0), .b(s_284), .O(gate142inter1));
  and2  gate2537(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate2538(.a(s_284), .O(gate142inter3));
  inv1  gate2539(.a(s_285), .O(gate142inter4));
  nand2 gate2540(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate2541(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate2542(.a(G456), .O(gate142inter7));
  inv1  gate2543(.a(G459), .O(gate142inter8));
  nand2 gate2544(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate2545(.a(s_285), .b(gate142inter3), .O(gate142inter10));
  nor2  gate2546(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate2547(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate2548(.a(gate142inter12), .b(gate142inter1), .O(G537));
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate2213(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate2214(.a(gate144inter0), .b(s_238), .O(gate144inter1));
  and2  gate2215(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate2216(.a(s_238), .O(gate144inter3));
  inv1  gate2217(.a(s_239), .O(gate144inter4));
  nand2 gate2218(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate2219(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate2220(.a(G468), .O(gate144inter7));
  inv1  gate2221(.a(G471), .O(gate144inter8));
  nand2 gate2222(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate2223(.a(s_239), .b(gate144inter3), .O(gate144inter10));
  nor2  gate2224(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate2225(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate2226(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate2689(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate2690(.a(gate151inter0), .b(s_306), .O(gate151inter1));
  and2  gate2691(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate2692(.a(s_306), .O(gate151inter3));
  inv1  gate2693(.a(s_307), .O(gate151inter4));
  nand2 gate2694(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate2695(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate2696(.a(G510), .O(gate151inter7));
  inv1  gate2697(.a(G513), .O(gate151inter8));
  nand2 gate2698(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate2699(.a(s_307), .b(gate151inter3), .O(gate151inter10));
  nor2  gate2700(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate2701(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate2702(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate897(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate898(.a(gate153inter0), .b(s_50), .O(gate153inter1));
  and2  gate899(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate900(.a(s_50), .O(gate153inter3));
  inv1  gate901(.a(s_51), .O(gate153inter4));
  nand2 gate902(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate903(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate904(.a(G426), .O(gate153inter7));
  inv1  gate905(.a(G522), .O(gate153inter8));
  nand2 gate906(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate907(.a(s_51), .b(gate153inter3), .O(gate153inter10));
  nor2  gate908(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate909(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate910(.a(gate153inter12), .b(gate153inter1), .O(G570));

  xor2  gate687(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate688(.a(gate154inter0), .b(s_20), .O(gate154inter1));
  and2  gate689(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate690(.a(s_20), .O(gate154inter3));
  inv1  gate691(.a(s_21), .O(gate154inter4));
  nand2 gate692(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate693(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate694(.a(G429), .O(gate154inter7));
  inv1  gate695(.a(G522), .O(gate154inter8));
  nand2 gate696(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate697(.a(s_21), .b(gate154inter3), .O(gate154inter10));
  nor2  gate698(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate699(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate700(.a(gate154inter12), .b(gate154inter1), .O(G571));

  xor2  gate2101(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate2102(.a(gate155inter0), .b(s_222), .O(gate155inter1));
  and2  gate2103(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate2104(.a(s_222), .O(gate155inter3));
  inv1  gate2105(.a(s_223), .O(gate155inter4));
  nand2 gate2106(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate2107(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate2108(.a(G432), .O(gate155inter7));
  inv1  gate2109(.a(G525), .O(gate155inter8));
  nand2 gate2110(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate2111(.a(s_223), .b(gate155inter3), .O(gate155inter10));
  nor2  gate2112(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate2113(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate2114(.a(gate155inter12), .b(gate155inter1), .O(G572));

  xor2  gate1709(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate1710(.a(gate156inter0), .b(s_166), .O(gate156inter1));
  and2  gate1711(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate1712(.a(s_166), .O(gate156inter3));
  inv1  gate1713(.a(s_167), .O(gate156inter4));
  nand2 gate1714(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate1715(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate1716(.a(G435), .O(gate156inter7));
  inv1  gate1717(.a(G525), .O(gate156inter8));
  nand2 gate1718(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate1719(.a(s_167), .b(gate156inter3), .O(gate156inter10));
  nor2  gate1720(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate1721(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate1722(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate645(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate646(.a(gate158inter0), .b(s_14), .O(gate158inter1));
  and2  gate647(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate648(.a(s_14), .O(gate158inter3));
  inv1  gate649(.a(s_15), .O(gate158inter4));
  nand2 gate650(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate651(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate652(.a(G441), .O(gate158inter7));
  inv1  gate653(.a(G528), .O(gate158inter8));
  nand2 gate654(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate655(.a(s_15), .b(gate158inter3), .O(gate158inter10));
  nor2  gate656(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate657(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate658(.a(gate158inter12), .b(gate158inter1), .O(G575));

  xor2  gate1793(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate1794(.a(gate159inter0), .b(s_178), .O(gate159inter1));
  and2  gate1795(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate1796(.a(s_178), .O(gate159inter3));
  inv1  gate1797(.a(s_179), .O(gate159inter4));
  nand2 gate1798(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate1799(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate1800(.a(G444), .O(gate159inter7));
  inv1  gate1801(.a(G531), .O(gate159inter8));
  nand2 gate1802(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate1803(.a(s_179), .b(gate159inter3), .O(gate159inter10));
  nor2  gate1804(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate1805(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate1806(.a(gate159inter12), .b(gate159inter1), .O(G576));

  xor2  gate2507(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate2508(.a(gate160inter0), .b(s_280), .O(gate160inter1));
  and2  gate2509(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate2510(.a(s_280), .O(gate160inter3));
  inv1  gate2511(.a(s_281), .O(gate160inter4));
  nand2 gate2512(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate2513(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate2514(.a(G447), .O(gate160inter7));
  inv1  gate2515(.a(G531), .O(gate160inter8));
  nand2 gate2516(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate2517(.a(s_281), .b(gate160inter3), .O(gate160inter10));
  nor2  gate2518(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate2519(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate2520(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate2577(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate2578(.a(gate162inter0), .b(s_290), .O(gate162inter1));
  and2  gate2579(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate2580(.a(s_290), .O(gate162inter3));
  inv1  gate2581(.a(s_291), .O(gate162inter4));
  nand2 gate2582(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate2583(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate2584(.a(G453), .O(gate162inter7));
  inv1  gate2585(.a(G534), .O(gate162inter8));
  nand2 gate2586(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate2587(.a(s_291), .b(gate162inter3), .O(gate162inter10));
  nor2  gate2588(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate2589(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate2590(.a(gate162inter12), .b(gate162inter1), .O(G579));

  xor2  gate757(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate758(.a(gate163inter0), .b(s_30), .O(gate163inter1));
  and2  gate759(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate760(.a(s_30), .O(gate163inter3));
  inv1  gate761(.a(s_31), .O(gate163inter4));
  nand2 gate762(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate763(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate764(.a(G456), .O(gate163inter7));
  inv1  gate765(.a(G537), .O(gate163inter8));
  nand2 gate766(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate767(.a(s_31), .b(gate163inter3), .O(gate163inter10));
  nor2  gate768(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate769(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate770(.a(gate163inter12), .b(gate163inter1), .O(G580));

  xor2  gate2549(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate2550(.a(gate164inter0), .b(s_286), .O(gate164inter1));
  and2  gate2551(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate2552(.a(s_286), .O(gate164inter3));
  inv1  gate2553(.a(s_287), .O(gate164inter4));
  nand2 gate2554(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate2555(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate2556(.a(G459), .O(gate164inter7));
  inv1  gate2557(.a(G537), .O(gate164inter8));
  nand2 gate2558(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate2559(.a(s_287), .b(gate164inter3), .O(gate164inter10));
  nor2  gate2560(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate2561(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate2562(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );

  xor2  gate1205(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate1206(.a(gate167inter0), .b(s_94), .O(gate167inter1));
  and2  gate1207(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate1208(.a(s_94), .O(gate167inter3));
  inv1  gate1209(.a(s_95), .O(gate167inter4));
  nand2 gate1210(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate1211(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate1212(.a(G468), .O(gate167inter7));
  inv1  gate1213(.a(G543), .O(gate167inter8));
  nand2 gate1214(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate1215(.a(s_95), .b(gate167inter3), .O(gate167inter10));
  nor2  gate1216(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate1217(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate1218(.a(gate167inter12), .b(gate167inter1), .O(G584));
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate1765(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate1766(.a(gate170inter0), .b(s_174), .O(gate170inter1));
  and2  gate1767(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate1768(.a(s_174), .O(gate170inter3));
  inv1  gate1769(.a(s_175), .O(gate170inter4));
  nand2 gate1770(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate1771(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate1772(.a(G477), .O(gate170inter7));
  inv1  gate1773(.a(G546), .O(gate170inter8));
  nand2 gate1774(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate1775(.a(s_175), .b(gate170inter3), .O(gate170inter10));
  nor2  gate1776(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate1777(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate1778(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate1863(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate1864(.a(gate172inter0), .b(s_188), .O(gate172inter1));
  and2  gate1865(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate1866(.a(s_188), .O(gate172inter3));
  inv1  gate1867(.a(s_189), .O(gate172inter4));
  nand2 gate1868(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate1869(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate1870(.a(G483), .O(gate172inter7));
  inv1  gate1871(.a(G549), .O(gate172inter8));
  nand2 gate1872(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate1873(.a(s_189), .b(gate172inter3), .O(gate172inter10));
  nor2  gate1874(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate1875(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate1876(.a(gate172inter12), .b(gate172inter1), .O(G589));

  xor2  gate603(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate604(.a(gate173inter0), .b(s_8), .O(gate173inter1));
  and2  gate605(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate606(.a(s_8), .O(gate173inter3));
  inv1  gate607(.a(s_9), .O(gate173inter4));
  nand2 gate608(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate609(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate610(.a(G486), .O(gate173inter7));
  inv1  gate611(.a(G552), .O(gate173inter8));
  nand2 gate612(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate613(.a(s_9), .b(gate173inter3), .O(gate173inter10));
  nor2  gate614(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate615(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate616(.a(gate173inter12), .b(gate173inter1), .O(G590));

  xor2  gate1485(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate1486(.a(gate174inter0), .b(s_134), .O(gate174inter1));
  and2  gate1487(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate1488(.a(s_134), .O(gate174inter3));
  inv1  gate1489(.a(s_135), .O(gate174inter4));
  nand2 gate1490(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate1491(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate1492(.a(G489), .O(gate174inter7));
  inv1  gate1493(.a(G552), .O(gate174inter8));
  nand2 gate1494(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate1495(.a(s_135), .b(gate174inter3), .O(gate174inter10));
  nor2  gate1496(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate1497(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate1498(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate1723(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate1724(.a(gate178inter0), .b(s_168), .O(gate178inter1));
  and2  gate1725(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate1726(.a(s_168), .O(gate178inter3));
  inv1  gate1727(.a(s_169), .O(gate178inter4));
  nand2 gate1728(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate1729(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate1730(.a(G501), .O(gate178inter7));
  inv1  gate1731(.a(G558), .O(gate178inter8));
  nand2 gate1732(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate1733(.a(s_169), .b(gate178inter3), .O(gate178inter10));
  nor2  gate1734(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate1735(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate1736(.a(gate178inter12), .b(gate178inter1), .O(G595));
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate715(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate716(.a(gate181inter0), .b(s_24), .O(gate181inter1));
  and2  gate717(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate718(.a(s_24), .O(gate181inter3));
  inv1  gate719(.a(s_25), .O(gate181inter4));
  nand2 gate720(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate721(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate722(.a(G510), .O(gate181inter7));
  inv1  gate723(.a(G564), .O(gate181inter8));
  nand2 gate724(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate725(.a(s_25), .b(gate181inter3), .O(gate181inter10));
  nor2  gate726(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate727(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate728(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate2087(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate2088(.a(gate183inter0), .b(s_220), .O(gate183inter1));
  and2  gate2089(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate2090(.a(s_220), .O(gate183inter3));
  inv1  gate2091(.a(s_221), .O(gate183inter4));
  nand2 gate2092(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate2093(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate2094(.a(G516), .O(gate183inter7));
  inv1  gate2095(.a(G567), .O(gate183inter8));
  nand2 gate2096(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate2097(.a(s_221), .b(gate183inter3), .O(gate183inter10));
  nor2  gate2098(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate2099(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate2100(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate1177(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1178(.a(gate186inter0), .b(s_90), .O(gate186inter1));
  and2  gate1179(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1180(.a(s_90), .O(gate186inter3));
  inv1  gate1181(.a(s_91), .O(gate186inter4));
  nand2 gate1182(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1183(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1184(.a(G572), .O(gate186inter7));
  inv1  gate1185(.a(G573), .O(gate186inter8));
  nand2 gate1186(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1187(.a(s_91), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1188(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1189(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1190(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate1611(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate1612(.a(gate190inter0), .b(s_152), .O(gate190inter1));
  and2  gate1613(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate1614(.a(s_152), .O(gate190inter3));
  inv1  gate1615(.a(s_153), .O(gate190inter4));
  nand2 gate1616(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate1617(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate1618(.a(G580), .O(gate190inter7));
  inv1  gate1619(.a(G581), .O(gate190inter8));
  nand2 gate1620(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate1621(.a(s_153), .b(gate190inter3), .O(gate190inter10));
  nor2  gate1622(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate1623(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate1624(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate2423(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate2424(.a(gate193inter0), .b(s_268), .O(gate193inter1));
  and2  gate2425(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate2426(.a(s_268), .O(gate193inter3));
  inv1  gate2427(.a(s_269), .O(gate193inter4));
  nand2 gate2428(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate2429(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate2430(.a(G586), .O(gate193inter7));
  inv1  gate2431(.a(G587), .O(gate193inter8));
  nand2 gate2432(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate2433(.a(s_269), .b(gate193inter3), .O(gate193inter10));
  nor2  gate2434(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate2435(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate2436(.a(gate193inter12), .b(gate193inter1), .O(G642));

  xor2  gate1163(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate1164(.a(gate194inter0), .b(s_88), .O(gate194inter1));
  and2  gate1165(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate1166(.a(s_88), .O(gate194inter3));
  inv1  gate1167(.a(s_89), .O(gate194inter4));
  nand2 gate1168(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate1169(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate1170(.a(G588), .O(gate194inter7));
  inv1  gate1171(.a(G589), .O(gate194inter8));
  nand2 gate1172(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate1173(.a(s_89), .b(gate194inter3), .O(gate194inter10));
  nor2  gate1174(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate1175(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate1176(.a(gate194inter12), .b(gate194inter1), .O(G645));
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate1639(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate1640(.a(gate196inter0), .b(s_156), .O(gate196inter1));
  and2  gate1641(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate1642(.a(s_156), .O(gate196inter3));
  inv1  gate1643(.a(s_157), .O(gate196inter4));
  nand2 gate1644(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate1645(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate1646(.a(G592), .O(gate196inter7));
  inv1  gate1647(.a(G593), .O(gate196inter8));
  nand2 gate1648(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate1649(.a(s_157), .b(gate196inter3), .O(gate196inter10));
  nor2  gate1650(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate1651(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate1652(.a(gate196inter12), .b(gate196inter1), .O(G651));

  xor2  gate2129(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate2130(.a(gate197inter0), .b(s_226), .O(gate197inter1));
  and2  gate2131(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate2132(.a(s_226), .O(gate197inter3));
  inv1  gate2133(.a(s_227), .O(gate197inter4));
  nand2 gate2134(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate2135(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate2136(.a(G594), .O(gate197inter7));
  inv1  gate2137(.a(G595), .O(gate197inter8));
  nand2 gate2138(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate2139(.a(s_227), .b(gate197inter3), .O(gate197inter10));
  nor2  gate2140(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate2141(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate2142(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );

  xor2  gate1443(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate1444(.a(gate199inter0), .b(s_128), .O(gate199inter1));
  and2  gate1445(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate1446(.a(s_128), .O(gate199inter3));
  inv1  gate1447(.a(s_129), .O(gate199inter4));
  nand2 gate1448(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate1449(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate1450(.a(G598), .O(gate199inter7));
  inv1  gate1451(.a(G599), .O(gate199inter8));
  nand2 gate1452(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate1453(.a(s_129), .b(gate199inter3), .O(gate199inter10));
  nor2  gate1454(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate1455(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate1456(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate2633(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate2634(.a(gate203inter0), .b(s_298), .O(gate203inter1));
  and2  gate2635(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate2636(.a(s_298), .O(gate203inter3));
  inv1  gate2637(.a(s_299), .O(gate203inter4));
  nand2 gate2638(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate2639(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate2640(.a(G602), .O(gate203inter7));
  inv1  gate2641(.a(G612), .O(gate203inter8));
  nand2 gate2642(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate2643(.a(s_299), .b(gate203inter3), .O(gate203inter10));
  nor2  gate2644(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate2645(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate2646(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate1695(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate1696(.a(gate205inter0), .b(s_164), .O(gate205inter1));
  and2  gate1697(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate1698(.a(s_164), .O(gate205inter3));
  inv1  gate1699(.a(s_165), .O(gate205inter4));
  nand2 gate1700(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate1701(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate1702(.a(G622), .O(gate205inter7));
  inv1  gate1703(.a(G627), .O(gate205inter8));
  nand2 gate1704(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate1705(.a(s_165), .b(gate205inter3), .O(gate205inter10));
  nor2  gate1706(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate1707(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate1708(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );

  xor2  gate2675(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate2676(.a(gate208inter0), .b(s_304), .O(gate208inter1));
  and2  gate2677(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate2678(.a(s_304), .O(gate208inter3));
  inv1  gate2679(.a(s_305), .O(gate208inter4));
  nand2 gate2680(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate2681(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate2682(.a(G627), .O(gate208inter7));
  inv1  gate2683(.a(G637), .O(gate208inter8));
  nand2 gate2684(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate2685(.a(s_305), .b(gate208inter3), .O(gate208inter10));
  nor2  gate2686(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate2687(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate2688(.a(gate208inter12), .b(gate208inter1), .O(G687));
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate813(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate814(.a(gate213inter0), .b(s_38), .O(gate213inter1));
  and2  gate815(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate816(.a(s_38), .O(gate213inter3));
  inv1  gate817(.a(s_39), .O(gate213inter4));
  nand2 gate818(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate819(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate820(.a(G602), .O(gate213inter7));
  inv1  gate821(.a(G672), .O(gate213inter8));
  nand2 gate822(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate823(.a(s_39), .b(gate213inter3), .O(gate213inter10));
  nor2  gate824(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate825(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate826(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate953(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate954(.a(gate219inter0), .b(s_58), .O(gate219inter1));
  and2  gate955(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate956(.a(s_58), .O(gate219inter3));
  inv1  gate957(.a(s_59), .O(gate219inter4));
  nand2 gate958(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate959(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate960(.a(G632), .O(gate219inter7));
  inv1  gate961(.a(G681), .O(gate219inter8));
  nand2 gate962(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate963(.a(s_59), .b(gate219inter3), .O(gate219inter10));
  nor2  gate964(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate965(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate966(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate1009(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate1010(.a(gate226inter0), .b(s_66), .O(gate226inter1));
  and2  gate1011(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate1012(.a(s_66), .O(gate226inter3));
  inv1  gate1013(.a(s_67), .O(gate226inter4));
  nand2 gate1014(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate1015(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate1016(.a(G692), .O(gate226inter7));
  inv1  gate1017(.a(G693), .O(gate226inter8));
  nand2 gate1018(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate1019(.a(s_67), .b(gate226inter3), .O(gate226inter10));
  nor2  gate1020(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate1021(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate1022(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate2451(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate2452(.a(gate233inter0), .b(s_272), .O(gate233inter1));
  and2  gate2453(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate2454(.a(s_272), .O(gate233inter3));
  inv1  gate2455(.a(s_273), .O(gate233inter4));
  nand2 gate2456(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate2457(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate2458(.a(G242), .O(gate233inter7));
  inv1  gate2459(.a(G718), .O(gate233inter8));
  nand2 gate2460(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate2461(.a(s_273), .b(gate233inter3), .O(gate233inter10));
  nor2  gate2462(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate2463(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate2464(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );

  xor2  gate1989(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate1990(.a(gate235inter0), .b(s_206), .O(gate235inter1));
  and2  gate1991(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate1992(.a(s_206), .O(gate235inter3));
  inv1  gate1993(.a(s_207), .O(gate235inter4));
  nand2 gate1994(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate1995(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate1996(.a(G248), .O(gate235inter7));
  inv1  gate1997(.a(G724), .O(gate235inter8));
  nand2 gate1998(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate1999(.a(s_207), .b(gate235inter3), .O(gate235inter10));
  nor2  gate2000(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate2001(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate2002(.a(gate235inter12), .b(gate235inter1), .O(G736));

  xor2  gate2157(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate2158(.a(gate236inter0), .b(s_230), .O(gate236inter1));
  and2  gate2159(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate2160(.a(s_230), .O(gate236inter3));
  inv1  gate2161(.a(s_231), .O(gate236inter4));
  nand2 gate2162(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate2163(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate2164(.a(G251), .O(gate236inter7));
  inv1  gate2165(.a(G727), .O(gate236inter8));
  nand2 gate2166(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate2167(.a(s_231), .b(gate236inter3), .O(gate236inter10));
  nor2  gate2168(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate2169(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate2170(.a(gate236inter12), .b(gate236inter1), .O(G739));

  xor2  gate2465(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate2466(.a(gate237inter0), .b(s_274), .O(gate237inter1));
  and2  gate2467(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate2468(.a(s_274), .O(gate237inter3));
  inv1  gate2469(.a(s_275), .O(gate237inter4));
  nand2 gate2470(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate2471(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate2472(.a(G254), .O(gate237inter7));
  inv1  gate2473(.a(G706), .O(gate237inter8));
  nand2 gate2474(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate2475(.a(s_275), .b(gate237inter3), .O(gate237inter10));
  nor2  gate2476(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate2477(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate2478(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate2773(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate2774(.a(gate240inter0), .b(s_318), .O(gate240inter1));
  and2  gate2775(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate2776(.a(s_318), .O(gate240inter3));
  inv1  gate2777(.a(s_319), .O(gate240inter4));
  nand2 gate2778(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate2779(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate2780(.a(G263), .O(gate240inter7));
  inv1  gate2781(.a(G715), .O(gate240inter8));
  nand2 gate2782(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate2783(.a(s_319), .b(gate240inter3), .O(gate240inter10));
  nor2  gate2784(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate2785(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate2786(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate1513(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate1514(.a(gate249inter0), .b(s_138), .O(gate249inter1));
  and2  gate1515(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate1516(.a(s_138), .O(gate249inter3));
  inv1  gate1517(.a(s_139), .O(gate249inter4));
  nand2 gate1518(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate1519(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate1520(.a(G254), .O(gate249inter7));
  inv1  gate1521(.a(G742), .O(gate249inter8));
  nand2 gate1522(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate1523(.a(s_139), .b(gate249inter3), .O(gate249inter10));
  nor2  gate1524(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate1525(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate1526(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );

  xor2  gate1387(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate1388(.a(gate251inter0), .b(s_120), .O(gate251inter1));
  and2  gate1389(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate1390(.a(s_120), .O(gate251inter3));
  inv1  gate1391(.a(s_121), .O(gate251inter4));
  nand2 gate1392(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate1393(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate1394(.a(G257), .O(gate251inter7));
  inv1  gate1395(.a(G745), .O(gate251inter8));
  nand2 gate1396(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate1397(.a(s_121), .b(gate251inter3), .O(gate251inter10));
  nor2  gate1398(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate1399(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate1400(.a(gate251inter12), .b(gate251inter1), .O(G764));
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate2437(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate2438(.a(gate253inter0), .b(s_270), .O(gate253inter1));
  and2  gate2439(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate2440(.a(s_270), .O(gate253inter3));
  inv1  gate2441(.a(s_271), .O(gate253inter4));
  nand2 gate2442(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate2443(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate2444(.a(G260), .O(gate253inter7));
  inv1  gate2445(.a(G748), .O(gate253inter8));
  nand2 gate2446(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate2447(.a(s_271), .b(gate253inter3), .O(gate253inter10));
  nor2  gate2448(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate2449(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate2450(.a(gate253inter12), .b(gate253inter1), .O(G766));

  xor2  gate1569(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate1570(.a(gate254inter0), .b(s_146), .O(gate254inter1));
  and2  gate1571(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate1572(.a(s_146), .O(gate254inter3));
  inv1  gate1573(.a(s_147), .O(gate254inter4));
  nand2 gate1574(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate1575(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate1576(.a(G712), .O(gate254inter7));
  inv1  gate1577(.a(G748), .O(gate254inter8));
  nand2 gate1578(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate1579(.a(s_147), .b(gate254inter3), .O(gate254inter10));
  nor2  gate1580(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate1581(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate1582(.a(gate254inter12), .b(gate254inter1), .O(G767));

  xor2  gate1261(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate1262(.a(gate255inter0), .b(s_102), .O(gate255inter1));
  and2  gate1263(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate1264(.a(s_102), .O(gate255inter3));
  inv1  gate1265(.a(s_103), .O(gate255inter4));
  nand2 gate1266(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate1267(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate1268(.a(G263), .O(gate255inter7));
  inv1  gate1269(.a(G751), .O(gate255inter8));
  nand2 gate1270(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate1271(.a(s_103), .b(gate255inter3), .O(gate255inter10));
  nor2  gate1272(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate1273(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate1274(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate2059(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate2060(.a(gate262inter0), .b(s_216), .O(gate262inter1));
  and2  gate2061(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate2062(.a(s_216), .O(gate262inter3));
  inv1  gate2063(.a(s_217), .O(gate262inter4));
  nand2 gate2064(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate2065(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate2066(.a(G764), .O(gate262inter7));
  inv1  gate2067(.a(G765), .O(gate262inter8));
  nand2 gate2068(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate2069(.a(s_217), .b(gate262inter3), .O(gate262inter10));
  nor2  gate2070(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate2071(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate2072(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );

  xor2  gate2787(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate2788(.a(gate264inter0), .b(s_320), .O(gate264inter1));
  and2  gate2789(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate2790(.a(s_320), .O(gate264inter3));
  inv1  gate2791(.a(s_321), .O(gate264inter4));
  nand2 gate2792(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate2793(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate2794(.a(G768), .O(gate264inter7));
  inv1  gate2795(.a(G769), .O(gate264inter8));
  nand2 gate2796(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate2797(.a(s_321), .b(gate264inter3), .O(gate264inter10));
  nor2  gate2798(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate2799(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate2800(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate785(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate786(.a(gate270inter0), .b(s_34), .O(gate270inter1));
  and2  gate787(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate788(.a(s_34), .O(gate270inter3));
  inv1  gate789(.a(s_35), .O(gate270inter4));
  nand2 gate790(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate791(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate792(.a(G657), .O(gate270inter7));
  inv1  gate793(.a(G785), .O(gate270inter8));
  nand2 gate794(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate795(.a(s_35), .b(gate270inter3), .O(gate270inter10));
  nor2  gate796(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate797(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate798(.a(gate270inter12), .b(gate270inter1), .O(G809));
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );

  xor2  gate1233(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate1234(.a(gate273inter0), .b(s_98), .O(gate273inter1));
  and2  gate1235(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate1236(.a(s_98), .O(gate273inter3));
  inv1  gate1237(.a(s_99), .O(gate273inter4));
  nand2 gate1238(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate1239(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate1240(.a(G642), .O(gate273inter7));
  inv1  gate1241(.a(G794), .O(gate273inter8));
  nand2 gate1242(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate1243(.a(s_99), .b(gate273inter3), .O(gate273inter10));
  nor2  gate1244(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate1245(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate1246(.a(gate273inter12), .b(gate273inter1), .O(G818));

  xor2  gate2717(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate2718(.a(gate274inter0), .b(s_310), .O(gate274inter1));
  and2  gate2719(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate2720(.a(s_310), .O(gate274inter3));
  inv1  gate2721(.a(s_311), .O(gate274inter4));
  nand2 gate2722(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate2723(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate2724(.a(G770), .O(gate274inter7));
  inv1  gate2725(.a(G794), .O(gate274inter8));
  nand2 gate2726(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate2727(.a(s_311), .b(gate274inter3), .O(gate274inter10));
  nor2  gate2728(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate2729(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate2730(.a(gate274inter12), .b(gate274inter1), .O(G819));

  xor2  gate1051(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate1052(.a(gate275inter0), .b(s_72), .O(gate275inter1));
  and2  gate1053(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate1054(.a(s_72), .O(gate275inter3));
  inv1  gate1055(.a(s_73), .O(gate275inter4));
  nand2 gate1056(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate1057(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate1058(.a(G645), .O(gate275inter7));
  inv1  gate1059(.a(G797), .O(gate275inter8));
  nand2 gate1060(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate1061(.a(s_73), .b(gate275inter3), .O(gate275inter10));
  nor2  gate1062(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate1063(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate1064(.a(gate275inter12), .b(gate275inter1), .O(G820));

  xor2  gate2619(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate2620(.a(gate276inter0), .b(s_296), .O(gate276inter1));
  and2  gate2621(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate2622(.a(s_296), .O(gate276inter3));
  inv1  gate2623(.a(s_297), .O(gate276inter4));
  nand2 gate2624(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate2625(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate2626(.a(G773), .O(gate276inter7));
  inv1  gate2627(.a(G797), .O(gate276inter8));
  nand2 gate2628(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate2629(.a(s_297), .b(gate276inter3), .O(gate276inter10));
  nor2  gate2630(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate2631(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate2632(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate1401(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate1402(.a(gate278inter0), .b(s_122), .O(gate278inter1));
  and2  gate1403(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate1404(.a(s_122), .O(gate278inter3));
  inv1  gate1405(.a(s_123), .O(gate278inter4));
  nand2 gate1406(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate1407(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate1408(.a(G776), .O(gate278inter7));
  inv1  gate1409(.a(G800), .O(gate278inter8));
  nand2 gate1410(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate1411(.a(s_123), .b(gate278inter3), .O(gate278inter10));
  nor2  gate1412(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate1413(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate1414(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate2031(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate2032(.a(gate285inter0), .b(s_212), .O(gate285inter1));
  and2  gate2033(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate2034(.a(s_212), .O(gate285inter3));
  inv1  gate2035(.a(s_213), .O(gate285inter4));
  nand2 gate2036(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate2037(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate2038(.a(G660), .O(gate285inter7));
  inv1  gate2039(.a(G812), .O(gate285inter8));
  nand2 gate2040(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate2041(.a(s_213), .b(gate285inter3), .O(gate285inter10));
  nor2  gate2042(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate2043(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate2044(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate2563(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate2564(.a(gate287inter0), .b(s_288), .O(gate287inter1));
  and2  gate2565(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate2566(.a(s_288), .O(gate287inter3));
  inv1  gate2567(.a(s_289), .O(gate287inter4));
  nand2 gate2568(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate2569(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate2570(.a(G663), .O(gate287inter7));
  inv1  gate2571(.a(G815), .O(gate287inter8));
  nand2 gate2572(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate2573(.a(s_289), .b(gate287inter3), .O(gate287inter10));
  nor2  gate2574(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate2575(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate2576(.a(gate287inter12), .b(gate287inter1), .O(G832));

  xor2  gate855(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate856(.a(gate288inter0), .b(s_44), .O(gate288inter1));
  and2  gate857(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate858(.a(s_44), .O(gate288inter3));
  inv1  gate859(.a(s_45), .O(gate288inter4));
  nand2 gate860(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate861(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate862(.a(G791), .O(gate288inter7));
  inv1  gate863(.a(G815), .O(gate288inter8));
  nand2 gate864(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate865(.a(s_45), .b(gate288inter3), .O(gate288inter10));
  nor2  gate866(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate867(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate868(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate2269(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate2270(.a(gate290inter0), .b(s_246), .O(gate290inter1));
  and2  gate2271(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate2272(.a(s_246), .O(gate290inter3));
  inv1  gate2273(.a(s_247), .O(gate290inter4));
  nand2 gate2274(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate2275(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate2276(.a(G820), .O(gate290inter7));
  inv1  gate2277(.a(G821), .O(gate290inter8));
  nand2 gate2278(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate2279(.a(s_247), .b(gate290inter3), .O(gate290inter10));
  nor2  gate2280(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate2281(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate2282(.a(gate290inter12), .b(gate290inter1), .O(G847));

  xor2  gate617(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate618(.a(gate291inter0), .b(s_10), .O(gate291inter1));
  and2  gate619(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate620(.a(s_10), .O(gate291inter3));
  inv1  gate621(.a(s_11), .O(gate291inter4));
  nand2 gate622(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate623(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate624(.a(G822), .O(gate291inter7));
  inv1  gate625(.a(G823), .O(gate291inter8));
  nand2 gate626(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate627(.a(s_11), .b(gate291inter3), .O(gate291inter10));
  nor2  gate628(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate629(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate630(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate1107(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate1108(.a(gate293inter0), .b(s_80), .O(gate293inter1));
  and2  gate1109(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate1110(.a(s_80), .O(gate293inter3));
  inv1  gate1111(.a(s_81), .O(gate293inter4));
  nand2 gate1112(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate1113(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate1114(.a(G828), .O(gate293inter7));
  inv1  gate1115(.a(G829), .O(gate293inter8));
  nand2 gate1116(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate1117(.a(s_81), .b(gate293inter3), .O(gate293inter10));
  nor2  gate1118(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate1119(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate1120(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate2297(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate2298(.a(gate387inter0), .b(s_250), .O(gate387inter1));
  and2  gate2299(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate2300(.a(s_250), .O(gate387inter3));
  inv1  gate2301(.a(s_251), .O(gate387inter4));
  nand2 gate2302(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate2303(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate2304(.a(G1), .O(gate387inter7));
  inv1  gate2305(.a(G1036), .O(gate387inter8));
  nand2 gate2306(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate2307(.a(s_251), .b(gate387inter3), .O(gate387inter10));
  nor2  gate2308(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate2309(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate2310(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate2325(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate2326(.a(gate389inter0), .b(s_254), .O(gate389inter1));
  and2  gate2327(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate2328(.a(s_254), .O(gate389inter3));
  inv1  gate2329(.a(s_255), .O(gate389inter4));
  nand2 gate2330(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate2331(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate2332(.a(G3), .O(gate389inter7));
  inv1  gate2333(.a(G1042), .O(gate389inter8));
  nand2 gate2334(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate2335(.a(s_255), .b(gate389inter3), .O(gate389inter10));
  nor2  gate2336(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate2337(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate2338(.a(gate389inter12), .b(gate389inter1), .O(G1138));

  xor2  gate1527(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate1528(.a(gate390inter0), .b(s_140), .O(gate390inter1));
  and2  gate1529(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate1530(.a(s_140), .O(gate390inter3));
  inv1  gate1531(.a(s_141), .O(gate390inter4));
  nand2 gate1532(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate1533(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate1534(.a(G4), .O(gate390inter7));
  inv1  gate1535(.a(G1045), .O(gate390inter8));
  nand2 gate1536(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate1537(.a(s_141), .b(gate390inter3), .O(gate390inter10));
  nor2  gate1538(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate1539(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate1540(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );

  xor2  gate2255(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate2256(.a(gate392inter0), .b(s_244), .O(gate392inter1));
  and2  gate2257(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate2258(.a(s_244), .O(gate392inter3));
  inv1  gate2259(.a(s_245), .O(gate392inter4));
  nand2 gate2260(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate2261(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate2262(.a(G6), .O(gate392inter7));
  inv1  gate2263(.a(G1051), .O(gate392inter8));
  nand2 gate2264(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate2265(.a(s_245), .b(gate392inter3), .O(gate392inter10));
  nor2  gate2266(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate2267(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate2268(.a(gate392inter12), .b(gate392inter1), .O(G1147));

  xor2  gate1079(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate1080(.a(gate393inter0), .b(s_76), .O(gate393inter1));
  and2  gate1081(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate1082(.a(s_76), .O(gate393inter3));
  inv1  gate1083(.a(s_77), .O(gate393inter4));
  nand2 gate1084(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate1085(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate1086(.a(G7), .O(gate393inter7));
  inv1  gate1087(.a(G1054), .O(gate393inter8));
  nand2 gate1088(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate1089(.a(s_77), .b(gate393inter3), .O(gate393inter10));
  nor2  gate1090(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate1091(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate1092(.a(gate393inter12), .b(gate393inter1), .O(G1150));

  xor2  gate841(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate842(.a(gate394inter0), .b(s_42), .O(gate394inter1));
  and2  gate843(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate844(.a(s_42), .O(gate394inter3));
  inv1  gate845(.a(s_43), .O(gate394inter4));
  nand2 gate846(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate847(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate848(.a(G8), .O(gate394inter7));
  inv1  gate849(.a(G1057), .O(gate394inter8));
  nand2 gate850(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate851(.a(s_43), .b(gate394inter3), .O(gate394inter10));
  nor2  gate852(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate853(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate854(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate1065(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate1066(.a(gate397inter0), .b(s_74), .O(gate397inter1));
  and2  gate1067(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate1068(.a(s_74), .O(gate397inter3));
  inv1  gate1069(.a(s_75), .O(gate397inter4));
  nand2 gate1070(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate1071(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate1072(.a(G11), .O(gate397inter7));
  inv1  gate1073(.a(G1066), .O(gate397inter8));
  nand2 gate1074(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate1075(.a(s_75), .b(gate397inter3), .O(gate397inter10));
  nor2  gate1076(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate1077(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate1078(.a(gate397inter12), .b(gate397inter1), .O(G1162));

  xor2  gate1751(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate1752(.a(gate398inter0), .b(s_172), .O(gate398inter1));
  and2  gate1753(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate1754(.a(s_172), .O(gate398inter3));
  inv1  gate1755(.a(s_173), .O(gate398inter4));
  nand2 gate1756(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate1757(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate1758(.a(G12), .O(gate398inter7));
  inv1  gate1759(.a(G1069), .O(gate398inter8));
  nand2 gate1760(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate1761(.a(s_173), .b(gate398inter3), .O(gate398inter10));
  nor2  gate1762(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate1763(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate1764(.a(gate398inter12), .b(gate398inter1), .O(G1165));

  xor2  gate1471(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate1472(.a(gate399inter0), .b(s_132), .O(gate399inter1));
  and2  gate1473(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate1474(.a(s_132), .O(gate399inter3));
  inv1  gate1475(.a(s_133), .O(gate399inter4));
  nand2 gate1476(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate1477(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate1478(.a(G13), .O(gate399inter7));
  inv1  gate1479(.a(G1072), .O(gate399inter8));
  nand2 gate1480(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate1481(.a(s_133), .b(gate399inter3), .O(gate399inter10));
  nor2  gate1482(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate1483(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate1484(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );

  xor2  gate631(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate632(.a(gate401inter0), .b(s_12), .O(gate401inter1));
  and2  gate633(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate634(.a(s_12), .O(gate401inter3));
  inv1  gate635(.a(s_13), .O(gate401inter4));
  nand2 gate636(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate637(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate638(.a(G15), .O(gate401inter7));
  inv1  gate639(.a(G1078), .O(gate401inter8));
  nand2 gate640(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate641(.a(s_13), .b(gate401inter3), .O(gate401inter10));
  nor2  gate642(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate643(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate644(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );

  xor2  gate2745(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate2746(.a(gate405inter0), .b(s_314), .O(gate405inter1));
  and2  gate2747(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate2748(.a(s_314), .O(gate405inter3));
  inv1  gate2749(.a(s_315), .O(gate405inter4));
  nand2 gate2750(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate2751(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate2752(.a(G19), .O(gate405inter7));
  inv1  gate2753(.a(G1090), .O(gate405inter8));
  nand2 gate2754(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate2755(.a(s_315), .b(gate405inter3), .O(gate405inter10));
  nor2  gate2756(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate2757(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate2758(.a(gate405inter12), .b(gate405inter1), .O(G1186));
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate1975(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate1976(.a(gate407inter0), .b(s_204), .O(gate407inter1));
  and2  gate1977(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate1978(.a(s_204), .O(gate407inter3));
  inv1  gate1979(.a(s_205), .O(gate407inter4));
  nand2 gate1980(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate1981(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate1982(.a(G21), .O(gate407inter7));
  inv1  gate1983(.a(G1096), .O(gate407inter8));
  nand2 gate1984(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate1985(.a(s_205), .b(gate407inter3), .O(gate407inter10));
  nor2  gate1986(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate1987(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate1988(.a(gate407inter12), .b(gate407inter1), .O(G1192));

  xor2  gate1835(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate1836(.a(gate408inter0), .b(s_184), .O(gate408inter1));
  and2  gate1837(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate1838(.a(s_184), .O(gate408inter3));
  inv1  gate1839(.a(s_185), .O(gate408inter4));
  nand2 gate1840(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate1841(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate1842(.a(G22), .O(gate408inter7));
  inv1  gate1843(.a(G1099), .O(gate408inter8));
  nand2 gate1844(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate1845(.a(s_185), .b(gate408inter3), .O(gate408inter10));
  nor2  gate1846(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate1847(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate1848(.a(gate408inter12), .b(gate408inter1), .O(G1195));

  xor2  gate2073(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate2074(.a(gate409inter0), .b(s_218), .O(gate409inter1));
  and2  gate2075(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate2076(.a(s_218), .O(gate409inter3));
  inv1  gate2077(.a(s_219), .O(gate409inter4));
  nand2 gate2078(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate2079(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate2080(.a(G23), .O(gate409inter7));
  inv1  gate2081(.a(G1102), .O(gate409inter8));
  nand2 gate2082(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate2083(.a(s_219), .b(gate409inter3), .O(gate409inter10));
  nor2  gate2084(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate2085(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate2086(.a(gate409inter12), .b(gate409inter1), .O(G1198));

  xor2  gate2395(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate2396(.a(gate410inter0), .b(s_264), .O(gate410inter1));
  and2  gate2397(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate2398(.a(s_264), .O(gate410inter3));
  inv1  gate2399(.a(s_265), .O(gate410inter4));
  nand2 gate2400(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate2401(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate2402(.a(G24), .O(gate410inter7));
  inv1  gate2403(.a(G1105), .O(gate410inter8));
  nand2 gate2404(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate2405(.a(s_265), .b(gate410inter3), .O(gate410inter10));
  nor2  gate2406(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate2407(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate2408(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate2381(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate2382(.a(gate415inter0), .b(s_262), .O(gate415inter1));
  and2  gate2383(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate2384(.a(s_262), .O(gate415inter3));
  inv1  gate2385(.a(s_263), .O(gate415inter4));
  nand2 gate2386(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate2387(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate2388(.a(G29), .O(gate415inter7));
  inv1  gate2389(.a(G1120), .O(gate415inter8));
  nand2 gate2390(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate2391(.a(s_263), .b(gate415inter3), .O(gate415inter10));
  nor2  gate2392(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate2393(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate2394(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate2605(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate2606(.a(gate421inter0), .b(s_294), .O(gate421inter1));
  and2  gate2607(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate2608(.a(s_294), .O(gate421inter3));
  inv1  gate2609(.a(s_295), .O(gate421inter4));
  nand2 gate2610(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate2611(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate2612(.a(G2), .O(gate421inter7));
  inv1  gate2613(.a(G1135), .O(gate421inter8));
  nand2 gate2614(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate2615(.a(s_295), .b(gate421inter3), .O(gate421inter10));
  nor2  gate2616(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate2617(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate2618(.a(gate421inter12), .b(gate421inter1), .O(G1230));
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );

  xor2  gate2017(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate2018(.a(gate424inter0), .b(s_210), .O(gate424inter1));
  and2  gate2019(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate2020(.a(s_210), .O(gate424inter3));
  inv1  gate2021(.a(s_211), .O(gate424inter4));
  nand2 gate2022(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate2023(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate2024(.a(G1042), .O(gate424inter7));
  inv1  gate2025(.a(G1138), .O(gate424inter8));
  nand2 gate2026(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate2027(.a(s_211), .b(gate424inter3), .O(gate424inter10));
  nor2  gate2028(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate2029(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate2030(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate2409(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate2410(.a(gate431inter0), .b(s_266), .O(gate431inter1));
  and2  gate2411(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate2412(.a(s_266), .O(gate431inter3));
  inv1  gate2413(.a(s_267), .O(gate431inter4));
  nand2 gate2414(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate2415(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate2416(.a(G7), .O(gate431inter7));
  inv1  gate2417(.a(G1150), .O(gate431inter8));
  nand2 gate2418(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate2419(.a(s_267), .b(gate431inter3), .O(gate431inter10));
  nor2  gate2420(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate2421(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate2422(.a(gate431inter12), .b(gate431inter1), .O(G1240));

  xor2  gate2003(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate2004(.a(gate432inter0), .b(s_208), .O(gate432inter1));
  and2  gate2005(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate2006(.a(s_208), .O(gate432inter3));
  inv1  gate2007(.a(s_209), .O(gate432inter4));
  nand2 gate2008(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate2009(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate2010(.a(G1054), .O(gate432inter7));
  inv1  gate2011(.a(G1150), .O(gate432inter8));
  nand2 gate2012(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate2013(.a(s_209), .b(gate432inter3), .O(gate432inter10));
  nor2  gate2014(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate2015(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate2016(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate1429(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate1430(.a(gate434inter0), .b(s_126), .O(gate434inter1));
  and2  gate1431(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate1432(.a(s_126), .O(gate434inter3));
  inv1  gate1433(.a(s_127), .O(gate434inter4));
  nand2 gate1434(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate1435(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate1436(.a(G1057), .O(gate434inter7));
  inv1  gate1437(.a(G1153), .O(gate434inter8));
  nand2 gate1438(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate1439(.a(s_127), .b(gate434inter3), .O(gate434inter10));
  nor2  gate1440(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate1441(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate1442(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );

  xor2  gate2339(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate2340(.a(gate436inter0), .b(s_256), .O(gate436inter1));
  and2  gate2341(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate2342(.a(s_256), .O(gate436inter3));
  inv1  gate2343(.a(s_257), .O(gate436inter4));
  nand2 gate2344(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate2345(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate2346(.a(G1060), .O(gate436inter7));
  inv1  gate2347(.a(G1156), .O(gate436inter8));
  nand2 gate2348(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate2349(.a(s_257), .b(gate436inter3), .O(gate436inter10));
  nor2  gate2350(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate2351(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate2352(.a(gate436inter12), .b(gate436inter1), .O(G1245));
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate1681(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate1682(.a(gate439inter0), .b(s_162), .O(gate439inter1));
  and2  gate1683(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate1684(.a(s_162), .O(gate439inter3));
  inv1  gate1685(.a(s_163), .O(gate439inter4));
  nand2 gate1686(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate1687(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate1688(.a(G11), .O(gate439inter7));
  inv1  gate1689(.a(G1162), .O(gate439inter8));
  nand2 gate1690(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate1691(.a(s_163), .b(gate439inter3), .O(gate439inter10));
  nor2  gate1692(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate1693(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate1694(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate799(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate800(.a(gate441inter0), .b(s_36), .O(gate441inter1));
  and2  gate801(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate802(.a(s_36), .O(gate441inter3));
  inv1  gate803(.a(s_37), .O(gate441inter4));
  nand2 gate804(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate805(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate806(.a(G12), .O(gate441inter7));
  inv1  gate807(.a(G1165), .O(gate441inter8));
  nand2 gate808(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate809(.a(s_37), .b(gate441inter3), .O(gate441inter10));
  nor2  gate810(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate811(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate812(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate729(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate730(.a(gate444inter0), .b(s_26), .O(gate444inter1));
  and2  gate731(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate732(.a(s_26), .O(gate444inter3));
  inv1  gate733(.a(s_27), .O(gate444inter4));
  nand2 gate734(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate735(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate736(.a(G1072), .O(gate444inter7));
  inv1  gate737(.a(G1168), .O(gate444inter8));
  nand2 gate738(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate739(.a(s_27), .b(gate444inter3), .O(gate444inter10));
  nor2  gate740(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate741(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate742(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );

  xor2  gate2227(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate2228(.a(gate451inter0), .b(s_240), .O(gate451inter1));
  and2  gate2229(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate2230(.a(s_240), .O(gate451inter3));
  inv1  gate2231(.a(s_241), .O(gate451inter4));
  nand2 gate2232(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate2233(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate2234(.a(G17), .O(gate451inter7));
  inv1  gate2235(.a(G1180), .O(gate451inter8));
  nand2 gate2236(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate2237(.a(s_241), .b(gate451inter3), .O(gate451inter10));
  nor2  gate2238(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate2239(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate2240(.a(gate451inter12), .b(gate451inter1), .O(G1260));
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );

  xor2  gate2283(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate2284(.a(gate455inter0), .b(s_248), .O(gate455inter1));
  and2  gate2285(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate2286(.a(s_248), .O(gate455inter3));
  inv1  gate2287(.a(s_249), .O(gate455inter4));
  nand2 gate2288(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate2289(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate2290(.a(G19), .O(gate455inter7));
  inv1  gate2291(.a(G1186), .O(gate455inter8));
  nand2 gate2292(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate2293(.a(s_249), .b(gate455inter3), .O(gate455inter10));
  nor2  gate2294(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate2295(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate2296(.a(gate455inter12), .b(gate455inter1), .O(G1264));

  xor2  gate2647(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate2648(.a(gate456inter0), .b(s_300), .O(gate456inter1));
  and2  gate2649(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate2650(.a(s_300), .O(gate456inter3));
  inv1  gate2651(.a(s_301), .O(gate456inter4));
  nand2 gate2652(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate2653(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate2654(.a(G1090), .O(gate456inter7));
  inv1  gate2655(.a(G1186), .O(gate456inter8));
  nand2 gate2656(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate2657(.a(s_301), .b(gate456inter3), .O(gate456inter10));
  nor2  gate2658(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate2659(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate2660(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );

  xor2  gate827(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate828(.a(gate458inter0), .b(s_40), .O(gate458inter1));
  and2  gate829(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate830(.a(s_40), .O(gate458inter3));
  inv1  gate831(.a(s_41), .O(gate458inter4));
  nand2 gate832(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate833(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate834(.a(G1093), .O(gate458inter7));
  inv1  gate835(.a(G1189), .O(gate458inter8));
  nand2 gate836(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate837(.a(s_41), .b(gate458inter3), .O(gate458inter10));
  nor2  gate838(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate839(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate840(.a(gate458inter12), .b(gate458inter1), .O(G1267));
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate883(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate884(.a(gate460inter0), .b(s_48), .O(gate460inter1));
  and2  gate885(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate886(.a(s_48), .O(gate460inter3));
  inv1  gate887(.a(s_49), .O(gate460inter4));
  nand2 gate888(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate889(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate890(.a(G1096), .O(gate460inter7));
  inv1  gate891(.a(G1192), .O(gate460inter8));
  nand2 gate892(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate893(.a(s_49), .b(gate460inter3), .O(gate460inter10));
  nor2  gate894(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate895(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate896(.a(gate460inter12), .b(gate460inter1), .O(G1269));

  xor2  gate2493(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate2494(.a(gate461inter0), .b(s_278), .O(gate461inter1));
  and2  gate2495(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate2496(.a(s_278), .O(gate461inter3));
  inv1  gate2497(.a(s_279), .O(gate461inter4));
  nand2 gate2498(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate2499(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate2500(.a(G22), .O(gate461inter7));
  inv1  gate2501(.a(G1195), .O(gate461inter8));
  nand2 gate2502(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate2503(.a(s_279), .b(gate461inter3), .O(gate461inter10));
  nor2  gate2504(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate2505(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate2506(.a(gate461inter12), .b(gate461inter1), .O(G1270));
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate1359(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate1360(.a(gate463inter0), .b(s_116), .O(gate463inter1));
  and2  gate1361(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate1362(.a(s_116), .O(gate463inter3));
  inv1  gate1363(.a(s_117), .O(gate463inter4));
  nand2 gate1364(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate1365(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate1366(.a(G23), .O(gate463inter7));
  inv1  gate1367(.a(G1198), .O(gate463inter8));
  nand2 gate1368(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate1369(.a(s_117), .b(gate463inter3), .O(gate463inter10));
  nor2  gate1370(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate1371(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate1372(.a(gate463inter12), .b(gate463inter1), .O(G1272));

  xor2  gate1135(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate1136(.a(gate464inter0), .b(s_84), .O(gate464inter1));
  and2  gate1137(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate1138(.a(s_84), .O(gate464inter3));
  inv1  gate1139(.a(s_85), .O(gate464inter4));
  nand2 gate1140(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate1141(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate1142(.a(G1102), .O(gate464inter7));
  inv1  gate1143(.a(G1198), .O(gate464inter8));
  nand2 gate1144(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate1145(.a(s_85), .b(gate464inter3), .O(gate464inter10));
  nor2  gate1146(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate1147(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate1148(.a(gate464inter12), .b(gate464inter1), .O(G1273));

  xor2  gate1541(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate1542(.a(gate465inter0), .b(s_142), .O(gate465inter1));
  and2  gate1543(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate1544(.a(s_142), .O(gate465inter3));
  inv1  gate1545(.a(s_143), .O(gate465inter4));
  nand2 gate1546(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate1547(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate1548(.a(G24), .O(gate465inter7));
  inv1  gate1549(.a(G1201), .O(gate465inter8));
  nand2 gate1550(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate1551(.a(s_143), .b(gate465inter3), .O(gate465inter10));
  nor2  gate1552(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate1553(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate1554(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );

  xor2  gate869(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate870(.a(gate468inter0), .b(s_46), .O(gate468inter1));
  and2  gate871(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate872(.a(s_46), .O(gate468inter3));
  inv1  gate873(.a(s_47), .O(gate468inter4));
  nand2 gate874(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate875(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate876(.a(G1108), .O(gate468inter7));
  inv1  gate877(.a(G1204), .O(gate468inter8));
  nand2 gate878(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate879(.a(s_47), .b(gate468inter3), .O(gate468inter10));
  nor2  gate880(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate881(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate882(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate743(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate744(.a(gate474inter0), .b(s_28), .O(gate474inter1));
  and2  gate745(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate746(.a(s_28), .O(gate474inter3));
  inv1  gate747(.a(s_29), .O(gate474inter4));
  nand2 gate748(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate749(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate750(.a(G1117), .O(gate474inter7));
  inv1  gate751(.a(G1213), .O(gate474inter8));
  nand2 gate752(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate753(.a(s_29), .b(gate474inter3), .O(gate474inter10));
  nor2  gate754(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate755(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate756(.a(gate474inter12), .b(gate474inter1), .O(G1283));
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate995(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate996(.a(gate476inter0), .b(s_64), .O(gate476inter1));
  and2  gate997(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate998(.a(s_64), .O(gate476inter3));
  inv1  gate999(.a(s_65), .O(gate476inter4));
  nand2 gate1000(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate1001(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate1002(.a(G1120), .O(gate476inter7));
  inv1  gate1003(.a(G1216), .O(gate476inter8));
  nand2 gate1004(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate1005(.a(s_65), .b(gate476inter3), .O(gate476inter10));
  nor2  gate1006(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate1007(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate1008(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate1961(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate1962(.a(gate480inter0), .b(s_202), .O(gate480inter1));
  and2  gate1963(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate1964(.a(s_202), .O(gate480inter3));
  inv1  gate1965(.a(s_203), .O(gate480inter4));
  nand2 gate1966(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate1967(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate1968(.a(G1126), .O(gate480inter7));
  inv1  gate1969(.a(G1222), .O(gate480inter8));
  nand2 gate1970(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate1971(.a(s_203), .b(gate480inter3), .O(gate480inter10));
  nor2  gate1972(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate1973(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate1974(.a(gate480inter12), .b(gate480inter1), .O(G1289));

  xor2  gate1625(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate1626(.a(gate481inter0), .b(s_154), .O(gate481inter1));
  and2  gate1627(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate1628(.a(s_154), .O(gate481inter3));
  inv1  gate1629(.a(s_155), .O(gate481inter4));
  nand2 gate1630(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate1631(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate1632(.a(G32), .O(gate481inter7));
  inv1  gate1633(.a(G1225), .O(gate481inter8));
  nand2 gate1634(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate1635(.a(s_155), .b(gate481inter3), .O(gate481inter10));
  nor2  gate1636(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate1637(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate1638(.a(gate481inter12), .b(gate481inter1), .O(G1290));
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );

  xor2  gate1891(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate1892(.a(gate483inter0), .b(s_192), .O(gate483inter1));
  and2  gate1893(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate1894(.a(s_192), .O(gate483inter3));
  inv1  gate1895(.a(s_193), .O(gate483inter4));
  nand2 gate1896(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate1897(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate1898(.a(G1228), .O(gate483inter7));
  inv1  gate1899(.a(G1229), .O(gate483inter8));
  nand2 gate1900(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate1901(.a(s_193), .b(gate483inter3), .O(gate483inter10));
  nor2  gate1902(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate1903(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate1904(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate2591(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate2592(.a(gate490inter0), .b(s_292), .O(gate490inter1));
  and2  gate2593(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate2594(.a(s_292), .O(gate490inter3));
  inv1  gate2595(.a(s_293), .O(gate490inter4));
  nand2 gate2596(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate2597(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate2598(.a(G1242), .O(gate490inter7));
  inv1  gate2599(.a(G1243), .O(gate490inter8));
  nand2 gate2600(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate2601(.a(s_293), .b(gate490inter3), .O(gate490inter10));
  nor2  gate2602(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate2603(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate2604(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate1415(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1416(.a(gate494inter0), .b(s_124), .O(gate494inter1));
  and2  gate1417(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1418(.a(s_124), .O(gate494inter3));
  inv1  gate1419(.a(s_125), .O(gate494inter4));
  nand2 gate1420(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1421(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1422(.a(G1250), .O(gate494inter7));
  inv1  gate1423(.a(G1251), .O(gate494inter8));
  nand2 gate1424(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1425(.a(s_125), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1426(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1427(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1428(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate701(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate702(.a(gate496inter0), .b(s_22), .O(gate496inter1));
  and2  gate703(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate704(.a(s_22), .O(gate496inter3));
  inv1  gate705(.a(s_23), .O(gate496inter4));
  nand2 gate706(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate707(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate708(.a(G1254), .O(gate496inter7));
  inv1  gate709(.a(G1255), .O(gate496inter8));
  nand2 gate710(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate711(.a(s_23), .b(gate496inter3), .O(gate496inter10));
  nor2  gate712(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate713(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate714(.a(gate496inter12), .b(gate496inter1), .O(G1305));
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );

  xor2  gate967(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate968(.a(gate498inter0), .b(s_60), .O(gate498inter1));
  and2  gate969(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate970(.a(s_60), .O(gate498inter3));
  inv1  gate971(.a(s_61), .O(gate498inter4));
  nand2 gate972(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate973(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate974(.a(G1258), .O(gate498inter7));
  inv1  gate975(.a(G1259), .O(gate498inter8));
  nand2 gate976(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate977(.a(s_61), .b(gate498inter3), .O(gate498inter10));
  nor2  gate978(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate979(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate980(.a(gate498inter12), .b(gate498inter1), .O(G1307));
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate2311(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate2312(.a(gate501inter0), .b(s_252), .O(gate501inter1));
  and2  gate2313(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate2314(.a(s_252), .O(gate501inter3));
  inv1  gate2315(.a(s_253), .O(gate501inter4));
  nand2 gate2316(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate2317(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate2318(.a(G1264), .O(gate501inter7));
  inv1  gate2319(.a(G1265), .O(gate501inter8));
  nand2 gate2320(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate2321(.a(s_253), .b(gate501inter3), .O(gate501inter10));
  nor2  gate2322(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate2323(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate2324(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate589(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate590(.a(gate504inter0), .b(s_6), .O(gate504inter1));
  and2  gate591(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate592(.a(s_6), .O(gate504inter3));
  inv1  gate593(.a(s_7), .O(gate504inter4));
  nand2 gate594(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate595(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate596(.a(G1270), .O(gate504inter7));
  inv1  gate597(.a(G1271), .O(gate504inter8));
  nand2 gate598(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate599(.a(s_7), .b(gate504inter3), .O(gate504inter10));
  nor2  gate600(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate601(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate602(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate575(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate576(.a(gate506inter0), .b(s_4), .O(gate506inter1));
  and2  gate577(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate578(.a(s_4), .O(gate506inter3));
  inv1  gate579(.a(s_5), .O(gate506inter4));
  nand2 gate580(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate581(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate582(.a(G1274), .O(gate506inter7));
  inv1  gate583(.a(G1275), .O(gate506inter8));
  nand2 gate584(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate585(.a(s_5), .b(gate506inter3), .O(gate506inter10));
  nor2  gate586(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate587(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate588(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate547(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate548(.a(gate511inter0), .b(s_0), .O(gate511inter1));
  and2  gate549(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate550(.a(s_0), .O(gate511inter3));
  inv1  gate551(.a(s_1), .O(gate511inter4));
  nand2 gate552(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate553(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate554(.a(G1284), .O(gate511inter7));
  inv1  gate555(.a(G1285), .O(gate511inter8));
  nand2 gate556(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate557(.a(s_1), .b(gate511inter3), .O(gate511inter10));
  nor2  gate558(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate559(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate560(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate1373(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate1374(.a(gate514inter0), .b(s_118), .O(gate514inter1));
  and2  gate1375(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate1376(.a(s_118), .O(gate514inter3));
  inv1  gate1377(.a(s_119), .O(gate514inter4));
  nand2 gate1378(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate1379(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate1380(.a(G1290), .O(gate514inter7));
  inv1  gate1381(.a(G1291), .O(gate514inter8));
  nand2 gate1382(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate1383(.a(s_119), .b(gate514inter3), .O(gate514inter10));
  nor2  gate1384(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate1385(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate1386(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule