module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );

  xor2  gate645(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate646(.a(gate10inter0), .b(s_14), .O(gate10inter1));
  and2  gate647(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate648(.a(s_14), .O(gate10inter3));
  inv1  gate649(.a(s_15), .O(gate10inter4));
  nand2 gate650(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate651(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate652(.a(G3), .O(gate10inter7));
  inv1  gate653(.a(G4), .O(gate10inter8));
  nand2 gate654(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate655(.a(s_15), .b(gate10inter3), .O(gate10inter10));
  nor2  gate656(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate657(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate658(.a(gate10inter12), .b(gate10inter1), .O(G269));
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate1765(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate1766(.a(gate12inter0), .b(s_174), .O(gate12inter1));
  and2  gate1767(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate1768(.a(s_174), .O(gate12inter3));
  inv1  gate1769(.a(s_175), .O(gate12inter4));
  nand2 gate1770(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate1771(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate1772(.a(G7), .O(gate12inter7));
  inv1  gate1773(.a(G8), .O(gate12inter8));
  nand2 gate1774(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate1775(.a(s_175), .b(gate12inter3), .O(gate12inter10));
  nor2  gate1776(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate1777(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate1778(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );

  xor2  gate1149(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate1150(.a(gate14inter0), .b(s_86), .O(gate14inter1));
  and2  gate1151(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate1152(.a(s_86), .O(gate14inter3));
  inv1  gate1153(.a(s_87), .O(gate14inter4));
  nand2 gate1154(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate1155(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate1156(.a(G11), .O(gate14inter7));
  inv1  gate1157(.a(G12), .O(gate14inter8));
  nand2 gate1158(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate1159(.a(s_87), .b(gate14inter3), .O(gate14inter10));
  nor2  gate1160(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate1161(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate1162(.a(gate14inter12), .b(gate14inter1), .O(G281));

  xor2  gate1051(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate1052(.a(gate15inter0), .b(s_72), .O(gate15inter1));
  and2  gate1053(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate1054(.a(s_72), .O(gate15inter3));
  inv1  gate1055(.a(s_73), .O(gate15inter4));
  nand2 gate1056(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate1057(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate1058(.a(G13), .O(gate15inter7));
  inv1  gate1059(.a(G14), .O(gate15inter8));
  nand2 gate1060(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate1061(.a(s_73), .b(gate15inter3), .O(gate15inter10));
  nor2  gate1062(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate1063(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate1064(.a(gate15inter12), .b(gate15inter1), .O(G284));

  xor2  gate1233(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate1234(.a(gate16inter0), .b(s_98), .O(gate16inter1));
  and2  gate1235(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate1236(.a(s_98), .O(gate16inter3));
  inv1  gate1237(.a(s_99), .O(gate16inter4));
  nand2 gate1238(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate1239(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate1240(.a(G15), .O(gate16inter7));
  inv1  gate1241(.a(G16), .O(gate16inter8));
  nand2 gate1242(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate1243(.a(s_99), .b(gate16inter3), .O(gate16inter10));
  nor2  gate1244(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate1245(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate1246(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate1415(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate1416(.a(gate19inter0), .b(s_124), .O(gate19inter1));
  and2  gate1417(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate1418(.a(s_124), .O(gate19inter3));
  inv1  gate1419(.a(s_125), .O(gate19inter4));
  nand2 gate1420(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate1421(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate1422(.a(G21), .O(gate19inter7));
  inv1  gate1423(.a(G22), .O(gate19inter8));
  nand2 gate1424(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate1425(.a(s_125), .b(gate19inter3), .O(gate19inter10));
  nor2  gate1426(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate1427(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate1428(.a(gate19inter12), .b(gate19inter1), .O(G296));

  xor2  gate2045(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate2046(.a(gate20inter0), .b(s_214), .O(gate20inter1));
  and2  gate2047(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate2048(.a(s_214), .O(gate20inter3));
  inv1  gate2049(.a(s_215), .O(gate20inter4));
  nand2 gate2050(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate2051(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate2052(.a(G23), .O(gate20inter7));
  inv1  gate2053(.a(G24), .O(gate20inter8));
  nand2 gate2054(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate2055(.a(s_215), .b(gate20inter3), .O(gate20inter10));
  nor2  gate2056(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate2057(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate2058(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate1723(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate1724(.a(gate29inter0), .b(s_168), .O(gate29inter1));
  and2  gate1725(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate1726(.a(s_168), .O(gate29inter3));
  inv1  gate1727(.a(s_169), .O(gate29inter4));
  nand2 gate1728(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate1729(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate1730(.a(G3), .O(gate29inter7));
  inv1  gate1731(.a(G7), .O(gate29inter8));
  nand2 gate1732(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate1733(.a(s_169), .b(gate29inter3), .O(gate29inter10));
  nor2  gate1734(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate1735(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate1736(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate1639(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate1640(.a(gate31inter0), .b(s_156), .O(gate31inter1));
  and2  gate1641(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate1642(.a(s_156), .O(gate31inter3));
  inv1  gate1643(.a(s_157), .O(gate31inter4));
  nand2 gate1644(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate1645(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate1646(.a(G4), .O(gate31inter7));
  inv1  gate1647(.a(G8), .O(gate31inter8));
  nand2 gate1648(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate1649(.a(s_157), .b(gate31inter3), .O(gate31inter10));
  nor2  gate1650(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate1651(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate1652(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate1107(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate1108(.a(gate33inter0), .b(s_80), .O(gate33inter1));
  and2  gate1109(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate1110(.a(s_80), .O(gate33inter3));
  inv1  gate1111(.a(s_81), .O(gate33inter4));
  nand2 gate1112(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate1113(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate1114(.a(G17), .O(gate33inter7));
  inv1  gate1115(.a(G21), .O(gate33inter8));
  nand2 gate1116(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate1117(.a(s_81), .b(gate33inter3), .O(gate33inter10));
  nor2  gate1118(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate1119(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate1120(.a(gate33inter12), .b(gate33inter1), .O(G338));
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate1569(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate1570(.a(gate39inter0), .b(s_146), .O(gate39inter1));
  and2  gate1571(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate1572(.a(s_146), .O(gate39inter3));
  inv1  gate1573(.a(s_147), .O(gate39inter4));
  nand2 gate1574(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate1575(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate1576(.a(G20), .O(gate39inter7));
  inv1  gate1577(.a(G24), .O(gate39inter8));
  nand2 gate1578(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate1579(.a(s_147), .b(gate39inter3), .O(gate39inter10));
  nor2  gate1580(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate1581(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate1582(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate995(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate996(.a(gate44inter0), .b(s_64), .O(gate44inter1));
  and2  gate997(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate998(.a(s_64), .O(gate44inter3));
  inv1  gate999(.a(s_65), .O(gate44inter4));
  nand2 gate1000(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate1001(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate1002(.a(G4), .O(gate44inter7));
  inv1  gate1003(.a(G269), .O(gate44inter8));
  nand2 gate1004(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate1005(.a(s_65), .b(gate44inter3), .O(gate44inter10));
  nor2  gate1006(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate1007(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate1008(.a(gate44inter12), .b(gate44inter1), .O(G365));

  xor2  gate1471(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate1472(.a(gate45inter0), .b(s_132), .O(gate45inter1));
  and2  gate1473(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate1474(.a(s_132), .O(gate45inter3));
  inv1  gate1475(.a(s_133), .O(gate45inter4));
  nand2 gate1476(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate1477(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate1478(.a(G5), .O(gate45inter7));
  inv1  gate1479(.a(G272), .O(gate45inter8));
  nand2 gate1480(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate1481(.a(s_133), .b(gate45inter3), .O(gate45inter10));
  nor2  gate1482(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate1483(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate1484(.a(gate45inter12), .b(gate45inter1), .O(G366));
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );

  xor2  gate1709(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate1710(.a(gate48inter0), .b(s_166), .O(gate48inter1));
  and2  gate1711(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate1712(.a(s_166), .O(gate48inter3));
  inv1  gate1713(.a(s_167), .O(gate48inter4));
  nand2 gate1714(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate1715(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate1716(.a(G8), .O(gate48inter7));
  inv1  gate1717(.a(G275), .O(gate48inter8));
  nand2 gate1718(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate1719(.a(s_167), .b(gate48inter3), .O(gate48inter10));
  nor2  gate1720(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate1721(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate1722(.a(gate48inter12), .b(gate48inter1), .O(G369));
nand2 gate49( .a(G9), .b(G278), .O(G370) );

  xor2  gate1555(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate1556(.a(gate50inter0), .b(s_144), .O(gate50inter1));
  and2  gate1557(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate1558(.a(s_144), .O(gate50inter3));
  inv1  gate1559(.a(s_145), .O(gate50inter4));
  nand2 gate1560(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate1561(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate1562(.a(G10), .O(gate50inter7));
  inv1  gate1563(.a(G278), .O(gate50inter8));
  nand2 gate1564(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate1565(.a(s_145), .b(gate50inter3), .O(gate50inter10));
  nor2  gate1566(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate1567(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate1568(.a(gate50inter12), .b(gate50inter1), .O(G371));
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate603(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate604(.a(gate52inter0), .b(s_8), .O(gate52inter1));
  and2  gate605(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate606(.a(s_8), .O(gate52inter3));
  inv1  gate607(.a(s_9), .O(gate52inter4));
  nand2 gate608(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate609(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate610(.a(G12), .O(gate52inter7));
  inv1  gate611(.a(G281), .O(gate52inter8));
  nand2 gate612(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate613(.a(s_9), .b(gate52inter3), .O(gate52inter10));
  nor2  gate614(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate615(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate616(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate1079(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate1080(.a(gate55inter0), .b(s_76), .O(gate55inter1));
  and2  gate1081(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate1082(.a(s_76), .O(gate55inter3));
  inv1  gate1083(.a(s_77), .O(gate55inter4));
  nand2 gate1084(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate1085(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate1086(.a(G15), .O(gate55inter7));
  inv1  gate1087(.a(G287), .O(gate55inter8));
  nand2 gate1088(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate1089(.a(s_77), .b(gate55inter3), .O(gate55inter10));
  nor2  gate1090(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate1091(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate1092(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate561(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate562(.a(gate57inter0), .b(s_2), .O(gate57inter1));
  and2  gate563(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate564(.a(s_2), .O(gate57inter3));
  inv1  gate565(.a(s_3), .O(gate57inter4));
  nand2 gate566(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate567(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate568(.a(G17), .O(gate57inter7));
  inv1  gate569(.a(G290), .O(gate57inter8));
  nand2 gate570(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate571(.a(s_3), .b(gate57inter3), .O(gate57inter10));
  nor2  gate572(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate573(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate574(.a(gate57inter12), .b(gate57inter1), .O(G378));
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate1163(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate1164(.a(gate62inter0), .b(s_88), .O(gate62inter1));
  and2  gate1165(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate1166(.a(s_88), .O(gate62inter3));
  inv1  gate1167(.a(s_89), .O(gate62inter4));
  nand2 gate1168(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate1169(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate1170(.a(G22), .O(gate62inter7));
  inv1  gate1171(.a(G296), .O(gate62inter8));
  nand2 gate1172(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate1173(.a(s_89), .b(gate62inter3), .O(gate62inter10));
  nor2  gate1174(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate1175(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate1176(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );

  xor2  gate575(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate576(.a(gate64inter0), .b(s_4), .O(gate64inter1));
  and2  gate577(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate578(.a(s_4), .O(gate64inter3));
  inv1  gate579(.a(s_5), .O(gate64inter4));
  nand2 gate580(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate581(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate582(.a(G24), .O(gate64inter7));
  inv1  gate583(.a(G299), .O(gate64inter8));
  nand2 gate584(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate585(.a(s_5), .b(gate64inter3), .O(gate64inter10));
  nor2  gate586(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate587(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate588(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate1191(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate1192(.a(gate71inter0), .b(s_92), .O(gate71inter1));
  and2  gate1193(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate1194(.a(s_92), .O(gate71inter3));
  inv1  gate1195(.a(s_93), .O(gate71inter4));
  nand2 gate1196(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate1197(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate1198(.a(G31), .O(gate71inter7));
  inv1  gate1199(.a(G311), .O(gate71inter8));
  nand2 gate1200(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate1201(.a(s_93), .b(gate71inter3), .O(gate71inter10));
  nor2  gate1202(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate1203(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate1204(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );

  xor2  gate1821(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate1822(.a(gate79inter0), .b(s_182), .O(gate79inter1));
  and2  gate1823(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate1824(.a(s_182), .O(gate79inter3));
  inv1  gate1825(.a(s_183), .O(gate79inter4));
  nand2 gate1826(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate1827(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate1828(.a(G10), .O(gate79inter7));
  inv1  gate1829(.a(G323), .O(gate79inter8));
  nand2 gate1830(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate1831(.a(s_183), .b(gate79inter3), .O(gate79inter10));
  nor2  gate1832(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate1833(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate1834(.a(gate79inter12), .b(gate79inter1), .O(G400));
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate687(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate688(.a(gate82inter0), .b(s_20), .O(gate82inter1));
  and2  gate689(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate690(.a(s_20), .O(gate82inter3));
  inv1  gate691(.a(s_21), .O(gate82inter4));
  nand2 gate692(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate693(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate694(.a(G7), .O(gate82inter7));
  inv1  gate695(.a(G326), .O(gate82inter8));
  nand2 gate696(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate697(.a(s_21), .b(gate82inter3), .O(gate82inter10));
  nor2  gate698(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate699(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate700(.a(gate82inter12), .b(gate82inter1), .O(G403));

  xor2  gate631(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate632(.a(gate83inter0), .b(s_12), .O(gate83inter1));
  and2  gate633(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate634(.a(s_12), .O(gate83inter3));
  inv1  gate635(.a(s_13), .O(gate83inter4));
  nand2 gate636(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate637(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate638(.a(G11), .O(gate83inter7));
  inv1  gate639(.a(G329), .O(gate83inter8));
  nand2 gate640(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate641(.a(s_13), .b(gate83inter3), .O(gate83inter10));
  nor2  gate642(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate643(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate644(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate771(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate772(.a(gate94inter0), .b(s_32), .O(gate94inter1));
  and2  gate773(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate774(.a(s_32), .O(gate94inter3));
  inv1  gate775(.a(s_33), .O(gate94inter4));
  nand2 gate776(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate777(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate778(.a(G22), .O(gate94inter7));
  inv1  gate779(.a(G344), .O(gate94inter8));
  nand2 gate780(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate781(.a(s_33), .b(gate94inter3), .O(gate94inter10));
  nor2  gate782(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate783(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate784(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate953(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate954(.a(gate99inter0), .b(s_58), .O(gate99inter1));
  and2  gate955(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate956(.a(s_58), .O(gate99inter3));
  inv1  gate957(.a(s_59), .O(gate99inter4));
  nand2 gate958(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate959(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate960(.a(G27), .O(gate99inter7));
  inv1  gate961(.a(G353), .O(gate99inter8));
  nand2 gate962(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate963(.a(s_59), .b(gate99inter3), .O(gate99inter10));
  nor2  gate964(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate965(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate966(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );

  xor2  gate1863(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate1864(.a(gate101inter0), .b(s_188), .O(gate101inter1));
  and2  gate1865(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate1866(.a(s_188), .O(gate101inter3));
  inv1  gate1867(.a(s_189), .O(gate101inter4));
  nand2 gate1868(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate1869(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate1870(.a(G20), .O(gate101inter7));
  inv1  gate1871(.a(G356), .O(gate101inter8));
  nand2 gate1872(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate1873(.a(s_189), .b(gate101inter3), .O(gate101inter10));
  nor2  gate1874(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate1875(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate1876(.a(gate101inter12), .b(gate101inter1), .O(G422));

  xor2  gate799(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate800(.a(gate102inter0), .b(s_36), .O(gate102inter1));
  and2  gate801(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate802(.a(s_36), .O(gate102inter3));
  inv1  gate803(.a(s_37), .O(gate102inter4));
  nand2 gate804(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate805(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate806(.a(G24), .O(gate102inter7));
  inv1  gate807(.a(G356), .O(gate102inter8));
  nand2 gate808(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate809(.a(s_37), .b(gate102inter3), .O(gate102inter10));
  nor2  gate810(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate811(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate812(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate1807(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate1808(.a(gate107inter0), .b(s_180), .O(gate107inter1));
  and2  gate1809(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate1810(.a(s_180), .O(gate107inter3));
  inv1  gate1811(.a(s_181), .O(gate107inter4));
  nand2 gate1812(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate1813(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate1814(.a(G366), .O(gate107inter7));
  inv1  gate1815(.a(G367), .O(gate107inter8));
  nand2 gate1816(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate1817(.a(s_181), .b(gate107inter3), .O(gate107inter10));
  nor2  gate1818(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate1819(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate1820(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate1317(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate1318(.a(gate112inter0), .b(s_110), .O(gate112inter1));
  and2  gate1319(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate1320(.a(s_110), .O(gate112inter3));
  inv1  gate1321(.a(s_111), .O(gate112inter4));
  nand2 gate1322(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate1323(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate1324(.a(G376), .O(gate112inter7));
  inv1  gate1325(.a(G377), .O(gate112inter8));
  nand2 gate1326(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate1327(.a(s_111), .b(gate112inter3), .O(gate112inter10));
  nor2  gate1328(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate1329(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate1330(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate785(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate786(.a(gate116inter0), .b(s_34), .O(gate116inter1));
  and2  gate787(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate788(.a(s_34), .O(gate116inter3));
  inv1  gate789(.a(s_35), .O(gate116inter4));
  nand2 gate790(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate791(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate792(.a(G384), .O(gate116inter7));
  inv1  gate793(.a(G385), .O(gate116inter8));
  nand2 gate794(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate795(.a(s_35), .b(gate116inter3), .O(gate116inter10));
  nor2  gate796(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate797(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate798(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate869(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate870(.a(gate119inter0), .b(s_46), .O(gate119inter1));
  and2  gate871(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate872(.a(s_46), .O(gate119inter3));
  inv1  gate873(.a(s_47), .O(gate119inter4));
  nand2 gate874(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate875(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate876(.a(G390), .O(gate119inter7));
  inv1  gate877(.a(G391), .O(gate119inter8));
  nand2 gate878(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate879(.a(s_47), .b(gate119inter3), .O(gate119inter10));
  nor2  gate880(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate881(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate882(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate1443(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate1444(.a(gate121inter0), .b(s_128), .O(gate121inter1));
  and2  gate1445(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate1446(.a(s_128), .O(gate121inter3));
  inv1  gate1447(.a(s_129), .O(gate121inter4));
  nand2 gate1448(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate1449(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate1450(.a(G394), .O(gate121inter7));
  inv1  gate1451(.a(G395), .O(gate121inter8));
  nand2 gate1452(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate1453(.a(s_129), .b(gate121inter3), .O(gate121inter10));
  nor2  gate1454(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate1455(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate1456(.a(gate121inter12), .b(gate121inter1), .O(G474));

  xor2  gate1373(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate1374(.a(gate122inter0), .b(s_118), .O(gate122inter1));
  and2  gate1375(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate1376(.a(s_118), .O(gate122inter3));
  inv1  gate1377(.a(s_119), .O(gate122inter4));
  nand2 gate1378(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate1379(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate1380(.a(G396), .O(gate122inter7));
  inv1  gate1381(.a(G397), .O(gate122inter8));
  nand2 gate1382(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate1383(.a(s_119), .b(gate122inter3), .O(gate122inter10));
  nor2  gate1384(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate1385(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate1386(.a(gate122inter12), .b(gate122inter1), .O(G477));
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );

  xor2  gate1275(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate1276(.a(gate129inter0), .b(s_104), .O(gate129inter1));
  and2  gate1277(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate1278(.a(s_104), .O(gate129inter3));
  inv1  gate1279(.a(s_105), .O(gate129inter4));
  nand2 gate1280(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate1281(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate1282(.a(G410), .O(gate129inter7));
  inv1  gate1283(.a(G411), .O(gate129inter8));
  nand2 gate1284(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate1285(.a(s_105), .b(gate129inter3), .O(gate129inter10));
  nor2  gate1286(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate1287(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate1288(.a(gate129inter12), .b(gate129inter1), .O(G498));
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate1681(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate1682(.a(gate132inter0), .b(s_162), .O(gate132inter1));
  and2  gate1683(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate1684(.a(s_162), .O(gate132inter3));
  inv1  gate1685(.a(s_163), .O(gate132inter4));
  nand2 gate1686(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate1687(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate1688(.a(G416), .O(gate132inter7));
  inv1  gate1689(.a(G417), .O(gate132inter8));
  nand2 gate1690(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate1691(.a(s_163), .b(gate132inter3), .O(gate132inter10));
  nor2  gate1692(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate1693(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate1694(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate1751(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate1752(.a(gate138inter0), .b(s_172), .O(gate138inter1));
  and2  gate1753(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate1754(.a(s_172), .O(gate138inter3));
  inv1  gate1755(.a(s_173), .O(gate138inter4));
  nand2 gate1756(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate1757(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate1758(.a(G432), .O(gate138inter7));
  inv1  gate1759(.a(G435), .O(gate138inter8));
  nand2 gate1760(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate1761(.a(s_173), .b(gate138inter3), .O(gate138inter10));
  nor2  gate1762(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate1763(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate1764(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );

  xor2  gate2073(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate2074(.a(gate145inter0), .b(s_218), .O(gate145inter1));
  and2  gate2075(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate2076(.a(s_218), .O(gate145inter3));
  inv1  gate2077(.a(s_219), .O(gate145inter4));
  nand2 gate2078(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate2079(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate2080(.a(G474), .O(gate145inter7));
  inv1  gate2081(.a(G477), .O(gate145inter8));
  nand2 gate2082(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate2083(.a(s_219), .b(gate145inter3), .O(gate145inter10));
  nor2  gate2084(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate2085(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate2086(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate1583(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate1584(.a(gate151inter0), .b(s_148), .O(gate151inter1));
  and2  gate1585(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate1586(.a(s_148), .O(gate151inter3));
  inv1  gate1587(.a(s_149), .O(gate151inter4));
  nand2 gate1588(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate1589(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate1590(.a(G510), .O(gate151inter7));
  inv1  gate1591(.a(G513), .O(gate151inter8));
  nand2 gate1592(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate1593(.a(s_149), .b(gate151inter3), .O(gate151inter10));
  nor2  gate1594(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate1595(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate1596(.a(gate151inter12), .b(gate151inter1), .O(G564));

  xor2  gate547(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate548(.a(gate152inter0), .b(s_0), .O(gate152inter1));
  and2  gate549(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate550(.a(s_0), .O(gate152inter3));
  inv1  gate551(.a(s_1), .O(gate152inter4));
  nand2 gate552(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate553(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate554(.a(G516), .O(gate152inter7));
  inv1  gate555(.a(G519), .O(gate152inter8));
  nand2 gate556(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate557(.a(s_1), .b(gate152inter3), .O(gate152inter10));
  nor2  gate558(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate559(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate560(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate2031(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate2032(.a(gate155inter0), .b(s_212), .O(gate155inter1));
  and2  gate2033(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate2034(.a(s_212), .O(gate155inter3));
  inv1  gate2035(.a(s_213), .O(gate155inter4));
  nand2 gate2036(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate2037(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate2038(.a(G432), .O(gate155inter7));
  inv1  gate2039(.a(G525), .O(gate155inter8));
  nand2 gate2040(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate2041(.a(s_213), .b(gate155inter3), .O(gate155inter10));
  nor2  gate2042(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate2043(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate2044(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate1919(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate1920(.a(gate157inter0), .b(s_196), .O(gate157inter1));
  and2  gate1921(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate1922(.a(s_196), .O(gate157inter3));
  inv1  gate1923(.a(s_197), .O(gate157inter4));
  nand2 gate1924(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate1925(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate1926(.a(G438), .O(gate157inter7));
  inv1  gate1927(.a(G528), .O(gate157inter8));
  nand2 gate1928(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate1929(.a(s_197), .b(gate157inter3), .O(gate157inter10));
  nor2  gate1930(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate1931(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate1932(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate1037(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate1038(.a(gate164inter0), .b(s_70), .O(gate164inter1));
  and2  gate1039(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate1040(.a(s_70), .O(gate164inter3));
  inv1  gate1041(.a(s_71), .O(gate164inter4));
  nand2 gate1042(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate1043(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate1044(.a(G459), .O(gate164inter7));
  inv1  gate1045(.a(G537), .O(gate164inter8));
  nand2 gate1046(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate1047(.a(s_71), .b(gate164inter3), .O(gate164inter10));
  nor2  gate1048(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate1049(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate1050(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );

  xor2  gate701(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate702(.a(gate168inter0), .b(s_22), .O(gate168inter1));
  and2  gate703(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate704(.a(s_22), .O(gate168inter3));
  inv1  gate705(.a(s_23), .O(gate168inter4));
  nand2 gate706(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate707(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate708(.a(G471), .O(gate168inter7));
  inv1  gate709(.a(G543), .O(gate168inter8));
  nand2 gate710(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate711(.a(s_23), .b(gate168inter3), .O(gate168inter10));
  nor2  gate712(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate713(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate714(.a(gate168inter12), .b(gate168inter1), .O(G585));
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate1485(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate1486(.a(gate170inter0), .b(s_134), .O(gate170inter1));
  and2  gate1487(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate1488(.a(s_134), .O(gate170inter3));
  inv1  gate1489(.a(s_135), .O(gate170inter4));
  nand2 gate1490(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate1491(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate1492(.a(G477), .O(gate170inter7));
  inv1  gate1493(.a(G546), .O(gate170inter8));
  nand2 gate1494(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate1495(.a(s_135), .b(gate170inter3), .O(gate170inter10));
  nor2  gate1496(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate1497(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate1498(.a(gate170inter12), .b(gate170inter1), .O(G587));

  xor2  gate1933(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate1934(.a(gate171inter0), .b(s_198), .O(gate171inter1));
  and2  gate1935(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate1936(.a(s_198), .O(gate171inter3));
  inv1  gate1937(.a(s_199), .O(gate171inter4));
  nand2 gate1938(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate1939(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate1940(.a(G480), .O(gate171inter7));
  inv1  gate1941(.a(G549), .O(gate171inter8));
  nand2 gate1942(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate1943(.a(s_199), .b(gate171inter3), .O(gate171inter10));
  nor2  gate1944(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate1945(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate1946(.a(gate171inter12), .b(gate171inter1), .O(G588));
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate911(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate912(.a(gate174inter0), .b(s_52), .O(gate174inter1));
  and2  gate913(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate914(.a(s_52), .O(gate174inter3));
  inv1  gate915(.a(s_53), .O(gate174inter4));
  nand2 gate916(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate917(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate918(.a(G489), .O(gate174inter7));
  inv1  gate919(.a(G552), .O(gate174inter8));
  nand2 gate920(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate921(.a(s_53), .b(gate174inter3), .O(gate174inter10));
  nor2  gate922(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate923(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate924(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate1429(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate1430(.a(gate178inter0), .b(s_126), .O(gate178inter1));
  and2  gate1431(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate1432(.a(s_126), .O(gate178inter3));
  inv1  gate1433(.a(s_127), .O(gate178inter4));
  nand2 gate1434(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate1435(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate1436(.a(G501), .O(gate178inter7));
  inv1  gate1437(.a(G558), .O(gate178inter8));
  nand2 gate1438(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate1439(.a(s_127), .b(gate178inter3), .O(gate178inter10));
  nor2  gate1440(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate1441(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate1442(.a(gate178inter12), .b(gate178inter1), .O(G595));
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );

  xor2  gate1065(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate1066(.a(gate182inter0), .b(s_74), .O(gate182inter1));
  and2  gate1067(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate1068(.a(s_74), .O(gate182inter3));
  inv1  gate1069(.a(s_75), .O(gate182inter4));
  nand2 gate1070(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate1071(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate1072(.a(G513), .O(gate182inter7));
  inv1  gate1073(.a(G564), .O(gate182inter8));
  nand2 gate1074(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate1075(.a(s_75), .b(gate182inter3), .O(gate182inter10));
  nor2  gate1076(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate1077(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate1078(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate1359(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate1360(.a(gate187inter0), .b(s_116), .O(gate187inter1));
  and2  gate1361(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate1362(.a(s_116), .O(gate187inter3));
  inv1  gate1363(.a(s_117), .O(gate187inter4));
  nand2 gate1364(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate1365(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate1366(.a(G574), .O(gate187inter7));
  inv1  gate1367(.a(G575), .O(gate187inter8));
  nand2 gate1368(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate1369(.a(s_117), .b(gate187inter3), .O(gate187inter10));
  nor2  gate1370(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate1371(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate1372(.a(gate187inter12), .b(gate187inter1), .O(G612));
nand2 gate188( .a(G576), .b(G577), .O(G617) );

  xor2  gate1093(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate1094(.a(gate189inter0), .b(s_78), .O(gate189inter1));
  and2  gate1095(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate1096(.a(s_78), .O(gate189inter3));
  inv1  gate1097(.a(s_79), .O(gate189inter4));
  nand2 gate1098(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate1099(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate1100(.a(G578), .O(gate189inter7));
  inv1  gate1101(.a(G579), .O(gate189inter8));
  nand2 gate1102(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate1103(.a(s_79), .b(gate189inter3), .O(gate189inter10));
  nor2  gate1104(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate1105(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate1106(.a(gate189inter12), .b(gate189inter1), .O(G622));

  xor2  gate715(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate716(.a(gate190inter0), .b(s_24), .O(gate190inter1));
  and2  gate717(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate718(.a(s_24), .O(gate190inter3));
  inv1  gate719(.a(s_25), .O(gate190inter4));
  nand2 gate720(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate721(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate722(.a(G580), .O(gate190inter7));
  inv1  gate723(.a(G581), .O(gate190inter8));
  nand2 gate724(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate725(.a(s_25), .b(gate190inter3), .O(gate190inter10));
  nor2  gate726(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate727(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate728(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );

  xor2  gate1401(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate1402(.a(gate192inter0), .b(s_122), .O(gate192inter1));
  and2  gate1403(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate1404(.a(s_122), .O(gate192inter3));
  inv1  gate1405(.a(s_123), .O(gate192inter4));
  nand2 gate1406(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate1407(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate1408(.a(G584), .O(gate192inter7));
  inv1  gate1409(.a(G585), .O(gate192inter8));
  nand2 gate1410(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate1411(.a(s_123), .b(gate192inter3), .O(gate192inter10));
  nor2  gate1412(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate1413(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate1414(.a(gate192inter12), .b(gate192inter1), .O(G637));

  xor2  gate1877(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate1878(.a(gate193inter0), .b(s_190), .O(gate193inter1));
  and2  gate1879(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate1880(.a(s_190), .O(gate193inter3));
  inv1  gate1881(.a(s_191), .O(gate193inter4));
  nand2 gate1882(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate1883(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate1884(.a(G586), .O(gate193inter7));
  inv1  gate1885(.a(G587), .O(gate193inter8));
  nand2 gate1886(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate1887(.a(s_191), .b(gate193inter3), .O(gate193inter10));
  nor2  gate1888(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate1889(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate1890(.a(gate193inter12), .b(gate193inter1), .O(G642));

  xor2  gate659(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate660(.a(gate194inter0), .b(s_16), .O(gate194inter1));
  and2  gate661(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate662(.a(s_16), .O(gate194inter3));
  inv1  gate663(.a(s_17), .O(gate194inter4));
  nand2 gate664(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate665(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate666(.a(G588), .O(gate194inter7));
  inv1  gate667(.a(G589), .O(gate194inter8));
  nand2 gate668(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate669(.a(s_17), .b(gate194inter3), .O(gate194inter10));
  nor2  gate670(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate671(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate672(.a(gate194inter12), .b(gate194inter1), .O(G645));
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate1793(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate1794(.a(gate196inter0), .b(s_178), .O(gate196inter1));
  and2  gate1795(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate1796(.a(s_178), .O(gate196inter3));
  inv1  gate1797(.a(s_179), .O(gate196inter4));
  nand2 gate1798(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate1799(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate1800(.a(G592), .O(gate196inter7));
  inv1  gate1801(.a(G593), .O(gate196inter8));
  nand2 gate1802(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate1803(.a(s_179), .b(gate196inter3), .O(gate196inter10));
  nor2  gate1804(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate1805(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate1806(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );

  xor2  gate1331(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate1332(.a(gate199inter0), .b(s_112), .O(gate199inter1));
  and2  gate1333(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate1334(.a(s_112), .O(gate199inter3));
  inv1  gate1335(.a(s_113), .O(gate199inter4));
  nand2 gate1336(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate1337(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate1338(.a(G598), .O(gate199inter7));
  inv1  gate1339(.a(G599), .O(gate199inter8));
  nand2 gate1340(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate1341(.a(s_113), .b(gate199inter3), .O(gate199inter10));
  nor2  gate1342(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate1343(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate1344(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );

  xor2  gate729(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate730(.a(gate202inter0), .b(s_26), .O(gate202inter1));
  and2  gate731(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate732(.a(s_26), .O(gate202inter3));
  inv1  gate733(.a(s_27), .O(gate202inter4));
  nand2 gate734(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate735(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate736(.a(G612), .O(gate202inter7));
  inv1  gate737(.a(G617), .O(gate202inter8));
  nand2 gate738(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate739(.a(s_27), .b(gate202inter3), .O(gate202inter10));
  nor2  gate740(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate741(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate742(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );

  xor2  gate673(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate674(.a(gate207inter0), .b(s_18), .O(gate207inter1));
  and2  gate675(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate676(.a(s_18), .O(gate207inter3));
  inv1  gate677(.a(s_19), .O(gate207inter4));
  nand2 gate678(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate679(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate680(.a(G622), .O(gate207inter7));
  inv1  gate681(.a(G632), .O(gate207inter8));
  nand2 gate682(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate683(.a(s_19), .b(gate207inter3), .O(gate207inter10));
  nor2  gate684(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate685(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate686(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );

  xor2  gate2003(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate2004(.a(gate217inter0), .b(s_208), .O(gate217inter1));
  and2  gate2005(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate2006(.a(s_208), .O(gate217inter3));
  inv1  gate2007(.a(s_209), .O(gate217inter4));
  nand2 gate2008(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate2009(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate2010(.a(G622), .O(gate217inter7));
  inv1  gate2011(.a(G678), .O(gate217inter8));
  nand2 gate2012(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate2013(.a(s_209), .b(gate217inter3), .O(gate217inter10));
  nor2  gate2014(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate2015(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate2016(.a(gate217inter12), .b(gate217inter1), .O(G698));

  xor2  gate617(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate618(.a(gate218inter0), .b(s_10), .O(gate218inter1));
  and2  gate619(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate620(.a(s_10), .O(gate218inter3));
  inv1  gate621(.a(s_11), .O(gate218inter4));
  nand2 gate622(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate623(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate624(.a(G627), .O(gate218inter7));
  inv1  gate625(.a(G678), .O(gate218inter8));
  nand2 gate626(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate627(.a(s_11), .b(gate218inter3), .O(gate218inter10));
  nor2  gate628(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate629(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate630(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate1023(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate1024(.a(gate220inter0), .b(s_68), .O(gate220inter1));
  and2  gate1025(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate1026(.a(s_68), .O(gate220inter3));
  inv1  gate1027(.a(s_69), .O(gate220inter4));
  nand2 gate1028(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate1029(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate1030(.a(G637), .O(gate220inter7));
  inv1  gate1031(.a(G681), .O(gate220inter8));
  nand2 gate1032(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate1033(.a(s_69), .b(gate220inter3), .O(gate220inter10));
  nor2  gate1034(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate1035(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate1036(.a(gate220inter12), .b(gate220inter1), .O(G701));
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate1891(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate1892(.a(gate224inter0), .b(s_192), .O(gate224inter1));
  and2  gate1893(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate1894(.a(s_192), .O(gate224inter3));
  inv1  gate1895(.a(s_193), .O(gate224inter4));
  nand2 gate1896(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate1897(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate1898(.a(G637), .O(gate224inter7));
  inv1  gate1899(.a(G687), .O(gate224inter8));
  nand2 gate1900(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate1901(.a(s_193), .b(gate224inter3), .O(gate224inter10));
  nor2  gate1902(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate1903(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate1904(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );

  xor2  gate1457(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate1458(.a(gate232inter0), .b(s_130), .O(gate232inter1));
  and2  gate1459(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate1460(.a(s_130), .O(gate232inter3));
  inv1  gate1461(.a(s_131), .O(gate232inter4));
  nand2 gate1462(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate1463(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate1464(.a(G704), .O(gate232inter7));
  inv1  gate1465(.a(G705), .O(gate232inter8));
  nand2 gate1466(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate1467(.a(s_131), .b(gate232inter3), .O(gate232inter10));
  nor2  gate1468(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate1469(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate1470(.a(gate232inter12), .b(gate232inter1), .O(G727));
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate1289(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate1290(.a(gate237inter0), .b(s_106), .O(gate237inter1));
  and2  gate1291(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate1292(.a(s_106), .O(gate237inter3));
  inv1  gate1293(.a(s_107), .O(gate237inter4));
  nand2 gate1294(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1295(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1296(.a(G254), .O(gate237inter7));
  inv1  gate1297(.a(G706), .O(gate237inter8));
  nand2 gate1298(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1299(.a(s_107), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1300(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1301(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1302(.a(gate237inter12), .b(gate237inter1), .O(G742));

  xor2  gate743(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate744(.a(gate238inter0), .b(s_28), .O(gate238inter1));
  and2  gate745(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate746(.a(s_28), .O(gate238inter3));
  inv1  gate747(.a(s_29), .O(gate238inter4));
  nand2 gate748(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate749(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate750(.a(G257), .O(gate238inter7));
  inv1  gate751(.a(G709), .O(gate238inter8));
  nand2 gate752(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate753(.a(s_29), .b(gate238inter3), .O(gate238inter10));
  nor2  gate754(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate755(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate756(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate925(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate926(.a(gate243inter0), .b(s_54), .O(gate243inter1));
  and2  gate927(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate928(.a(s_54), .O(gate243inter3));
  inv1  gate929(.a(s_55), .O(gate243inter4));
  nand2 gate930(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate931(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate932(.a(G245), .O(gate243inter7));
  inv1  gate933(.a(G733), .O(gate243inter8));
  nand2 gate934(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate935(.a(s_55), .b(gate243inter3), .O(gate243inter10));
  nor2  gate936(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate937(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate938(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate1625(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate1626(.a(gate248inter0), .b(s_154), .O(gate248inter1));
  and2  gate1627(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate1628(.a(s_154), .O(gate248inter3));
  inv1  gate1629(.a(s_155), .O(gate248inter4));
  nand2 gate1630(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate1631(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate1632(.a(G727), .O(gate248inter7));
  inv1  gate1633(.a(G739), .O(gate248inter8));
  nand2 gate1634(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate1635(.a(s_155), .b(gate248inter3), .O(gate248inter10));
  nor2  gate1636(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate1637(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate1638(.a(gate248inter12), .b(gate248inter1), .O(G761));

  xor2  gate1219(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate1220(.a(gate249inter0), .b(s_96), .O(gate249inter1));
  and2  gate1221(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate1222(.a(s_96), .O(gate249inter3));
  inv1  gate1223(.a(s_97), .O(gate249inter4));
  nand2 gate1224(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate1225(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate1226(.a(G254), .O(gate249inter7));
  inv1  gate1227(.a(G742), .O(gate249inter8));
  nand2 gate1228(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate1229(.a(s_97), .b(gate249inter3), .O(gate249inter10));
  nor2  gate1230(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate1231(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate1232(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate1905(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate1906(.a(gate258inter0), .b(s_194), .O(gate258inter1));
  and2  gate1907(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate1908(.a(s_194), .O(gate258inter3));
  inv1  gate1909(.a(s_195), .O(gate258inter4));
  nand2 gate1910(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate1911(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate1912(.a(G756), .O(gate258inter7));
  inv1  gate1913(.a(G757), .O(gate258inter8));
  nand2 gate1914(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate1915(.a(s_195), .b(gate258inter3), .O(gate258inter10));
  nor2  gate1916(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate1917(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate1918(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate1975(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate1976(.a(gate262inter0), .b(s_204), .O(gate262inter1));
  and2  gate1977(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate1978(.a(s_204), .O(gate262inter3));
  inv1  gate1979(.a(s_205), .O(gate262inter4));
  nand2 gate1980(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate1981(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate1982(.a(G764), .O(gate262inter7));
  inv1  gate1983(.a(G765), .O(gate262inter8));
  nand2 gate1984(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate1985(.a(s_205), .b(gate262inter3), .O(gate262inter10));
  nor2  gate1986(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate1987(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate1988(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );

  xor2  gate1541(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate1542(.a(gate264inter0), .b(s_142), .O(gate264inter1));
  and2  gate1543(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate1544(.a(s_142), .O(gate264inter3));
  inv1  gate1545(.a(s_143), .O(gate264inter4));
  nand2 gate1546(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate1547(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate1548(.a(G768), .O(gate264inter7));
  inv1  gate1549(.a(G769), .O(gate264inter8));
  nand2 gate1550(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate1551(.a(s_143), .b(gate264inter3), .O(gate264inter10));
  nor2  gate1552(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate1553(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate1554(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate1205(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate1206(.a(gate266inter0), .b(s_94), .O(gate266inter1));
  and2  gate1207(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate1208(.a(s_94), .O(gate266inter3));
  inv1  gate1209(.a(s_95), .O(gate266inter4));
  nand2 gate1210(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate1211(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate1212(.a(G645), .O(gate266inter7));
  inv1  gate1213(.a(G773), .O(gate266inter8));
  nand2 gate1214(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate1215(.a(s_95), .b(gate266inter3), .O(gate266inter10));
  nor2  gate1216(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate1217(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate1218(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate1387(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate1388(.a(gate268inter0), .b(s_120), .O(gate268inter1));
  and2  gate1389(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate1390(.a(s_120), .O(gate268inter3));
  inv1  gate1391(.a(s_121), .O(gate268inter4));
  nand2 gate1392(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1393(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1394(.a(G651), .O(gate268inter7));
  inv1  gate1395(.a(G779), .O(gate268inter8));
  nand2 gate1396(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1397(.a(s_121), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1398(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1399(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1400(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate1247(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate1248(.a(gate279inter0), .b(s_100), .O(gate279inter1));
  and2  gate1249(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate1250(.a(s_100), .O(gate279inter3));
  inv1  gate1251(.a(s_101), .O(gate279inter4));
  nand2 gate1252(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate1253(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate1254(.a(G651), .O(gate279inter7));
  inv1  gate1255(.a(G803), .O(gate279inter8));
  nand2 gate1256(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate1257(.a(s_101), .b(gate279inter3), .O(gate279inter10));
  nor2  gate1258(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate1259(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate1260(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate813(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate814(.a(gate283inter0), .b(s_38), .O(gate283inter1));
  and2  gate815(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate816(.a(s_38), .O(gate283inter3));
  inv1  gate817(.a(s_39), .O(gate283inter4));
  nand2 gate818(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate819(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate820(.a(G657), .O(gate283inter7));
  inv1  gate821(.a(G809), .O(gate283inter8));
  nand2 gate822(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate823(.a(s_39), .b(gate283inter3), .O(gate283inter10));
  nor2  gate824(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate825(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate826(.a(gate283inter12), .b(gate283inter1), .O(G828));

  xor2  gate841(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate842(.a(gate284inter0), .b(s_42), .O(gate284inter1));
  and2  gate843(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate844(.a(s_42), .O(gate284inter3));
  inv1  gate845(.a(s_43), .O(gate284inter4));
  nand2 gate846(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate847(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate848(.a(G785), .O(gate284inter7));
  inv1  gate849(.a(G809), .O(gate284inter8));
  nand2 gate850(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate851(.a(s_43), .b(gate284inter3), .O(gate284inter10));
  nor2  gate852(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate853(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate854(.a(gate284inter12), .b(gate284inter1), .O(G829));
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate1121(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate1122(.a(gate286inter0), .b(s_82), .O(gate286inter1));
  and2  gate1123(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate1124(.a(s_82), .O(gate286inter3));
  inv1  gate1125(.a(s_83), .O(gate286inter4));
  nand2 gate1126(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate1127(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate1128(.a(G788), .O(gate286inter7));
  inv1  gate1129(.a(G812), .O(gate286inter8));
  nand2 gate1130(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate1131(.a(s_83), .b(gate286inter3), .O(gate286inter10));
  nor2  gate1132(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate1133(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate1134(.a(gate286inter12), .b(gate286inter1), .O(G831));
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate2017(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate2018(.a(gate295inter0), .b(s_210), .O(gate295inter1));
  and2  gate2019(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate2020(.a(s_210), .O(gate295inter3));
  inv1  gate2021(.a(s_211), .O(gate295inter4));
  nand2 gate2022(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate2023(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate2024(.a(G830), .O(gate295inter7));
  inv1  gate2025(.a(G831), .O(gate295inter8));
  nand2 gate2026(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate2027(.a(s_211), .b(gate295inter3), .O(gate295inter10));
  nor2  gate2028(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate2029(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate2030(.a(gate295inter12), .b(gate295inter1), .O(G912));
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate1135(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate1136(.a(gate388inter0), .b(s_84), .O(gate388inter1));
  and2  gate1137(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate1138(.a(s_84), .O(gate388inter3));
  inv1  gate1139(.a(s_85), .O(gate388inter4));
  nand2 gate1140(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate1141(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate1142(.a(G2), .O(gate388inter7));
  inv1  gate1143(.a(G1039), .O(gate388inter8));
  nand2 gate1144(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate1145(.a(s_85), .b(gate388inter3), .O(gate388inter10));
  nor2  gate1146(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate1147(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate1148(.a(gate388inter12), .b(gate388inter1), .O(G1135));

  xor2  gate1303(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate1304(.a(gate389inter0), .b(s_108), .O(gate389inter1));
  and2  gate1305(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate1306(.a(s_108), .O(gate389inter3));
  inv1  gate1307(.a(s_109), .O(gate389inter4));
  nand2 gate1308(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate1309(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate1310(.a(G3), .O(gate389inter7));
  inv1  gate1311(.a(G1042), .O(gate389inter8));
  nand2 gate1312(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate1313(.a(s_109), .b(gate389inter3), .O(gate389inter10));
  nor2  gate1314(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate1315(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate1316(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate1989(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate1990(.a(gate400inter0), .b(s_206), .O(gate400inter1));
  and2  gate1991(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate1992(.a(s_206), .O(gate400inter3));
  inv1  gate1993(.a(s_207), .O(gate400inter4));
  nand2 gate1994(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate1995(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate1996(.a(G14), .O(gate400inter7));
  inv1  gate1997(.a(G1075), .O(gate400inter8));
  nand2 gate1998(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate1999(.a(s_207), .b(gate400inter3), .O(gate400inter10));
  nor2  gate2000(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate2001(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate2002(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate1513(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate1514(.a(gate402inter0), .b(s_138), .O(gate402inter1));
  and2  gate1515(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate1516(.a(s_138), .O(gate402inter3));
  inv1  gate1517(.a(s_139), .O(gate402inter4));
  nand2 gate1518(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate1519(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate1520(.a(G16), .O(gate402inter7));
  inv1  gate1521(.a(G1081), .O(gate402inter8));
  nand2 gate1522(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate1523(.a(s_139), .b(gate402inter3), .O(gate402inter10));
  nor2  gate1524(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate1525(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate1526(.a(gate402inter12), .b(gate402inter1), .O(G1177));
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );

  xor2  gate855(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate856(.a(gate405inter0), .b(s_44), .O(gate405inter1));
  and2  gate857(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate858(.a(s_44), .O(gate405inter3));
  inv1  gate859(.a(s_45), .O(gate405inter4));
  nand2 gate860(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate861(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate862(.a(G19), .O(gate405inter7));
  inv1  gate863(.a(G1090), .O(gate405inter8));
  nand2 gate864(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate865(.a(s_45), .b(gate405inter3), .O(gate405inter10));
  nor2  gate866(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate867(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate868(.a(gate405inter12), .b(gate405inter1), .O(G1186));
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate1961(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate1962(.a(gate407inter0), .b(s_202), .O(gate407inter1));
  and2  gate1963(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate1964(.a(s_202), .O(gate407inter3));
  inv1  gate1965(.a(s_203), .O(gate407inter4));
  nand2 gate1966(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate1967(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate1968(.a(G21), .O(gate407inter7));
  inv1  gate1969(.a(G1096), .O(gate407inter8));
  nand2 gate1970(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate1971(.a(s_203), .b(gate407inter3), .O(gate407inter10));
  nor2  gate1972(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate1973(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate1974(.a(gate407inter12), .b(gate407inter1), .O(G1192));

  xor2  gate589(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate590(.a(gate408inter0), .b(s_6), .O(gate408inter1));
  and2  gate591(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate592(.a(s_6), .O(gate408inter3));
  inv1  gate593(.a(s_7), .O(gate408inter4));
  nand2 gate594(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate595(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate596(.a(G22), .O(gate408inter7));
  inv1  gate597(.a(G1099), .O(gate408inter8));
  nand2 gate598(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate599(.a(s_7), .b(gate408inter3), .O(gate408inter10));
  nor2  gate600(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate601(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate602(.a(gate408inter12), .b(gate408inter1), .O(G1195));
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate1737(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate1738(.a(gate413inter0), .b(s_170), .O(gate413inter1));
  and2  gate1739(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate1740(.a(s_170), .O(gate413inter3));
  inv1  gate1741(.a(s_171), .O(gate413inter4));
  nand2 gate1742(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1743(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1744(.a(G27), .O(gate413inter7));
  inv1  gate1745(.a(G1114), .O(gate413inter8));
  nand2 gate1746(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1747(.a(s_171), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1748(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1749(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1750(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate939(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate940(.a(gate421inter0), .b(s_56), .O(gate421inter1));
  and2  gate941(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate942(.a(s_56), .O(gate421inter3));
  inv1  gate943(.a(s_57), .O(gate421inter4));
  nand2 gate944(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate945(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate946(.a(G2), .O(gate421inter7));
  inv1  gate947(.a(G1135), .O(gate421inter8));
  nand2 gate948(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate949(.a(s_57), .b(gate421inter3), .O(gate421inter10));
  nor2  gate950(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate951(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate952(.a(gate421inter12), .b(gate421inter1), .O(G1230));
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate1597(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate1598(.a(gate425inter0), .b(s_150), .O(gate425inter1));
  and2  gate1599(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate1600(.a(s_150), .O(gate425inter3));
  inv1  gate1601(.a(s_151), .O(gate425inter4));
  nand2 gate1602(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1603(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1604(.a(G4), .O(gate425inter7));
  inv1  gate1605(.a(G1141), .O(gate425inter8));
  nand2 gate1606(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1607(.a(s_151), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1608(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1609(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1610(.a(gate425inter12), .b(gate425inter1), .O(G1234));

  xor2  gate1009(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate1010(.a(gate426inter0), .b(s_66), .O(gate426inter1));
  and2  gate1011(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate1012(.a(s_66), .O(gate426inter3));
  inv1  gate1013(.a(s_67), .O(gate426inter4));
  nand2 gate1014(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate1015(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate1016(.a(G1045), .O(gate426inter7));
  inv1  gate1017(.a(G1141), .O(gate426inter8));
  nand2 gate1018(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate1019(.a(s_67), .b(gate426inter3), .O(gate426inter10));
  nor2  gate1020(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate1021(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate1022(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate1261(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate1262(.a(gate431inter0), .b(s_102), .O(gate431inter1));
  and2  gate1263(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate1264(.a(s_102), .O(gate431inter3));
  inv1  gate1265(.a(s_103), .O(gate431inter4));
  nand2 gate1266(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate1267(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate1268(.a(G7), .O(gate431inter7));
  inv1  gate1269(.a(G1150), .O(gate431inter8));
  nand2 gate1270(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate1271(.a(s_103), .b(gate431inter3), .O(gate431inter10));
  nor2  gate1272(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate1273(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate1274(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate1499(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate1500(.a(gate441inter0), .b(s_136), .O(gate441inter1));
  and2  gate1501(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate1502(.a(s_136), .O(gate441inter3));
  inv1  gate1503(.a(s_137), .O(gate441inter4));
  nand2 gate1504(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate1505(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate1506(.a(G12), .O(gate441inter7));
  inv1  gate1507(.a(G1165), .O(gate441inter8));
  nand2 gate1508(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate1509(.a(s_137), .b(gate441inter3), .O(gate441inter10));
  nor2  gate1510(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate1511(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate1512(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate967(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate968(.a(gate443inter0), .b(s_60), .O(gate443inter1));
  and2  gate969(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate970(.a(s_60), .O(gate443inter3));
  inv1  gate971(.a(s_61), .O(gate443inter4));
  nand2 gate972(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate973(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate974(.a(G13), .O(gate443inter7));
  inv1  gate975(.a(G1168), .O(gate443inter8));
  nand2 gate976(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate977(.a(s_61), .b(gate443inter3), .O(gate443inter10));
  nor2  gate978(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate979(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate980(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );

  xor2  gate1345(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate1346(.a(gate446inter0), .b(s_114), .O(gate446inter1));
  and2  gate1347(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate1348(.a(s_114), .O(gate446inter3));
  inv1  gate1349(.a(s_115), .O(gate446inter4));
  nand2 gate1350(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate1351(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate1352(.a(G1075), .O(gate446inter7));
  inv1  gate1353(.a(G1171), .O(gate446inter8));
  nand2 gate1354(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate1355(.a(s_115), .b(gate446inter3), .O(gate446inter10));
  nor2  gate1356(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate1357(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate1358(.a(gate446inter12), .b(gate446inter1), .O(G1255));
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );

  xor2  gate1653(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate1654(.a(gate451inter0), .b(s_158), .O(gate451inter1));
  and2  gate1655(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate1656(.a(s_158), .O(gate451inter3));
  inv1  gate1657(.a(s_159), .O(gate451inter4));
  nand2 gate1658(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate1659(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate1660(.a(G17), .O(gate451inter7));
  inv1  gate1661(.a(G1180), .O(gate451inter8));
  nand2 gate1662(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate1663(.a(s_159), .b(gate451inter3), .O(gate451inter10));
  nor2  gate1664(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate1665(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate1666(.a(gate451inter12), .b(gate451inter1), .O(G1260));

  xor2  gate897(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate898(.a(gate452inter0), .b(s_50), .O(gate452inter1));
  and2  gate899(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate900(.a(s_50), .O(gate452inter3));
  inv1  gate901(.a(s_51), .O(gate452inter4));
  nand2 gate902(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate903(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate904(.a(G1084), .O(gate452inter7));
  inv1  gate905(.a(G1180), .O(gate452inter8));
  nand2 gate906(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate907(.a(s_51), .b(gate452inter3), .O(gate452inter10));
  nor2  gate908(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate909(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate910(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate1779(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate1780(.a(gate463inter0), .b(s_176), .O(gate463inter1));
  and2  gate1781(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate1782(.a(s_176), .O(gate463inter3));
  inv1  gate1783(.a(s_177), .O(gate463inter4));
  nand2 gate1784(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate1785(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate1786(.a(G23), .O(gate463inter7));
  inv1  gate1787(.a(G1198), .O(gate463inter8));
  nand2 gate1788(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate1789(.a(s_177), .b(gate463inter3), .O(gate463inter10));
  nor2  gate1790(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate1791(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate1792(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate1527(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate1528(.a(gate466inter0), .b(s_140), .O(gate466inter1));
  and2  gate1529(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate1530(.a(s_140), .O(gate466inter3));
  inv1  gate1531(.a(s_141), .O(gate466inter4));
  nand2 gate1532(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate1533(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate1534(.a(G1105), .O(gate466inter7));
  inv1  gate1535(.a(G1201), .O(gate466inter8));
  nand2 gate1536(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate1537(.a(s_141), .b(gate466inter3), .O(gate466inter10));
  nor2  gate1538(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate1539(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate1540(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );

  xor2  gate827(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate828(.a(gate468inter0), .b(s_40), .O(gate468inter1));
  and2  gate829(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate830(.a(s_40), .O(gate468inter3));
  inv1  gate831(.a(s_41), .O(gate468inter4));
  nand2 gate832(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate833(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate834(.a(G1108), .O(gate468inter7));
  inv1  gate835(.a(G1204), .O(gate468inter8));
  nand2 gate836(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate837(.a(s_41), .b(gate468inter3), .O(gate468inter10));
  nor2  gate838(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate839(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate840(.a(gate468inter12), .b(gate468inter1), .O(G1277));

  xor2  gate883(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate884(.a(gate469inter0), .b(s_48), .O(gate469inter1));
  and2  gate885(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate886(.a(s_48), .O(gate469inter3));
  inv1  gate887(.a(s_49), .O(gate469inter4));
  nand2 gate888(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate889(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate890(.a(G26), .O(gate469inter7));
  inv1  gate891(.a(G1207), .O(gate469inter8));
  nand2 gate892(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate893(.a(s_49), .b(gate469inter3), .O(gate469inter10));
  nor2  gate894(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate895(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate896(.a(gate469inter12), .b(gate469inter1), .O(G1278));
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate1667(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate1668(.a(gate475inter0), .b(s_160), .O(gate475inter1));
  and2  gate1669(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate1670(.a(s_160), .O(gate475inter3));
  inv1  gate1671(.a(s_161), .O(gate475inter4));
  nand2 gate1672(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate1673(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate1674(.a(G29), .O(gate475inter7));
  inv1  gate1675(.a(G1216), .O(gate475inter8));
  nand2 gate1676(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate1677(.a(s_161), .b(gate475inter3), .O(gate475inter10));
  nor2  gate1678(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate1679(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate1680(.a(gate475inter12), .b(gate475inter1), .O(G1284));

  xor2  gate1611(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate1612(.a(gate476inter0), .b(s_152), .O(gate476inter1));
  and2  gate1613(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate1614(.a(s_152), .O(gate476inter3));
  inv1  gate1615(.a(s_153), .O(gate476inter4));
  nand2 gate1616(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate1617(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate1618(.a(G1120), .O(gate476inter7));
  inv1  gate1619(.a(G1216), .O(gate476inter8));
  nand2 gate1620(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate1621(.a(s_153), .b(gate476inter3), .O(gate476inter10));
  nor2  gate1622(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate1623(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate1624(.a(gate476inter12), .b(gate476inter1), .O(G1285));

  xor2  gate981(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate982(.a(gate477inter0), .b(s_62), .O(gate477inter1));
  and2  gate983(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate984(.a(s_62), .O(gate477inter3));
  inv1  gate985(.a(s_63), .O(gate477inter4));
  nand2 gate986(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate987(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate988(.a(G30), .O(gate477inter7));
  inv1  gate989(.a(G1219), .O(gate477inter8));
  nand2 gate990(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate991(.a(s_63), .b(gate477inter3), .O(gate477inter10));
  nor2  gate992(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate993(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate994(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );

  xor2  gate1835(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate1836(.a(gate479inter0), .b(s_184), .O(gate479inter1));
  and2  gate1837(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate1838(.a(s_184), .O(gate479inter3));
  inv1  gate1839(.a(s_185), .O(gate479inter4));
  nand2 gate1840(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate1841(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate1842(.a(G31), .O(gate479inter7));
  inv1  gate1843(.a(G1222), .O(gate479inter8));
  nand2 gate1844(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate1845(.a(s_185), .b(gate479inter3), .O(gate479inter10));
  nor2  gate1846(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate1847(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate1848(.a(gate479inter12), .b(gate479inter1), .O(G1288));

  xor2  gate2087(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate2088(.a(gate480inter0), .b(s_220), .O(gate480inter1));
  and2  gate2089(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate2090(.a(s_220), .O(gate480inter3));
  inv1  gate2091(.a(s_221), .O(gate480inter4));
  nand2 gate2092(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate2093(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate2094(.a(G1126), .O(gate480inter7));
  inv1  gate2095(.a(G1222), .O(gate480inter8));
  nand2 gate2096(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate2097(.a(s_221), .b(gate480inter3), .O(gate480inter10));
  nor2  gate2098(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate2099(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate2100(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );

  xor2  gate1695(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate1696(.a(gate483inter0), .b(s_164), .O(gate483inter1));
  and2  gate1697(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate1698(.a(s_164), .O(gate483inter3));
  inv1  gate1699(.a(s_165), .O(gate483inter4));
  nand2 gate1700(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate1701(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate1702(.a(G1228), .O(gate483inter7));
  inv1  gate1703(.a(G1229), .O(gate483inter8));
  nand2 gate1704(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate1705(.a(s_165), .b(gate483inter3), .O(gate483inter10));
  nor2  gate1706(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate1707(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate1708(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate1849(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate1850(.a(gate489inter0), .b(s_186), .O(gate489inter1));
  and2  gate1851(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate1852(.a(s_186), .O(gate489inter3));
  inv1  gate1853(.a(s_187), .O(gate489inter4));
  nand2 gate1854(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate1855(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate1856(.a(G1240), .O(gate489inter7));
  inv1  gate1857(.a(G1241), .O(gate489inter8));
  nand2 gate1858(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate1859(.a(s_187), .b(gate489inter3), .O(gate489inter10));
  nor2  gate1860(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate1861(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate1862(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate757(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate758(.a(gate494inter0), .b(s_30), .O(gate494inter1));
  and2  gate759(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate760(.a(s_30), .O(gate494inter3));
  inv1  gate761(.a(s_31), .O(gate494inter4));
  nand2 gate762(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate763(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate764(.a(G1250), .O(gate494inter7));
  inv1  gate765(.a(G1251), .O(gate494inter8));
  nand2 gate766(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate767(.a(s_31), .b(gate494inter3), .O(gate494inter10));
  nor2  gate768(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate769(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate770(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate1177(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate1178(.a(gate504inter0), .b(s_90), .O(gate504inter1));
  and2  gate1179(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate1180(.a(s_90), .O(gate504inter3));
  inv1  gate1181(.a(s_91), .O(gate504inter4));
  nand2 gate1182(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate1183(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate1184(.a(G1270), .O(gate504inter7));
  inv1  gate1185(.a(G1271), .O(gate504inter8));
  nand2 gate1186(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate1187(.a(s_91), .b(gate504inter3), .O(gate504inter10));
  nor2  gate1188(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate1189(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate1190(.a(gate504inter12), .b(gate504inter1), .O(G1313));

  xor2  gate2059(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate2060(.a(gate505inter0), .b(s_216), .O(gate505inter1));
  and2  gate2061(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate2062(.a(s_216), .O(gate505inter3));
  inv1  gate2063(.a(s_217), .O(gate505inter4));
  nand2 gate2064(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate2065(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate2066(.a(G1272), .O(gate505inter7));
  inv1  gate2067(.a(G1273), .O(gate505inter8));
  nand2 gate2068(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate2069(.a(s_217), .b(gate505inter3), .O(gate505inter10));
  nor2  gate2070(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate2071(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate2072(.a(gate505inter12), .b(gate505inter1), .O(G1314));
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate1947(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate1948(.a(gate511inter0), .b(s_200), .O(gate511inter1));
  and2  gate1949(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate1950(.a(s_200), .O(gate511inter3));
  inv1  gate1951(.a(s_201), .O(gate511inter4));
  nand2 gate1952(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate1953(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate1954(.a(G1284), .O(gate511inter7));
  inv1  gate1955(.a(G1285), .O(gate511inter8));
  nand2 gate1956(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate1957(.a(s_201), .b(gate511inter3), .O(gate511inter10));
  nor2  gate1958(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate1959(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate1960(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule