module c432 (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
             N430,N431,N432);
input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
      N99,N102,N105,N108,N112,N115;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91;
output N223,N329,N370,N421,N430,N431,N432;
wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12;


inv1 gate1( .a(N1), .O(N118) );
inv1 gate2( .a(N4), .O(N119) );
inv1 gate3( .a(N11), .O(N122) );
inv1 gate4( .a(N17), .O(N123) );
inv1 gate5( .a(N24), .O(N126) );
inv1 gate6( .a(N30), .O(N127) );
inv1 gate7( .a(N37), .O(N130) );
inv1 gate8( .a(N43), .O(N131) );
inv1 gate9( .a(N50), .O(N134) );
inv1 gate10( .a(N56), .O(N135) );
inv1 gate11( .a(N63), .O(N138) );
inv1 gate12( .a(N69), .O(N139) );
inv1 gate13( .a(N76), .O(N142) );
inv1 gate14( .a(N82), .O(N143) );
inv1 gate15( .a(N89), .O(N146) );
inv1 gate16( .a(N95), .O(N147) );
inv1 gate17( .a(N102), .O(N150) );
inv1 gate18( .a(N108), .O(N151) );
nand2 gate19( .a(N118), .b(N4), .O(N154) );
nor2 gate20( .a(N8), .b(N119), .O(N157) );

  xor2  gate385(.a(N119), .b(N14), .O(gate21inter0));
  nand2 gate386(.a(gate21inter0), .b(s_32), .O(gate21inter1));
  and2  gate387(.a(N119), .b(N14), .O(gate21inter2));
  inv1  gate388(.a(s_32), .O(gate21inter3));
  inv1  gate389(.a(s_33), .O(gate21inter4));
  nand2 gate390(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate391(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate392(.a(N14), .O(gate21inter7));
  inv1  gate393(.a(N119), .O(gate21inter8));
  nand2 gate394(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate395(.a(s_33), .b(gate21inter3), .O(gate21inter10));
  nor2  gate396(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate397(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate398(.a(gate21inter12), .b(gate21inter1), .O(N158));

  xor2  gate301(.a(N17), .b(N122), .O(gate22inter0));
  nand2 gate302(.a(gate22inter0), .b(s_20), .O(gate22inter1));
  and2  gate303(.a(N17), .b(N122), .O(gate22inter2));
  inv1  gate304(.a(s_20), .O(gate22inter3));
  inv1  gate305(.a(s_21), .O(gate22inter4));
  nand2 gate306(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate307(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate308(.a(N122), .O(gate22inter7));
  inv1  gate309(.a(N17), .O(gate22inter8));
  nand2 gate310(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate311(.a(s_21), .b(gate22inter3), .O(gate22inter10));
  nor2  gate312(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate313(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate314(.a(gate22inter12), .b(gate22inter1), .O(N159));
nand2 gate23( .a(N126), .b(N30), .O(N162) );
nand2 gate24( .a(N130), .b(N43), .O(N165) );
nand2 gate25( .a(N134), .b(N56), .O(N168) );

  xor2  gate259(.a(N69), .b(N138), .O(gate26inter0));
  nand2 gate260(.a(gate26inter0), .b(s_14), .O(gate26inter1));
  and2  gate261(.a(N69), .b(N138), .O(gate26inter2));
  inv1  gate262(.a(s_14), .O(gate26inter3));
  inv1  gate263(.a(s_15), .O(gate26inter4));
  nand2 gate264(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate265(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate266(.a(N138), .O(gate26inter7));
  inv1  gate267(.a(N69), .O(gate26inter8));
  nand2 gate268(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate269(.a(s_15), .b(gate26inter3), .O(gate26inter10));
  nor2  gate270(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate271(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate272(.a(gate26inter12), .b(gate26inter1), .O(N171));
nand2 gate27( .a(N142), .b(N82), .O(N174) );

  xor2  gate413(.a(N95), .b(N146), .O(gate28inter0));
  nand2 gate414(.a(gate28inter0), .b(s_36), .O(gate28inter1));
  and2  gate415(.a(N95), .b(N146), .O(gate28inter2));
  inv1  gate416(.a(s_36), .O(gate28inter3));
  inv1  gate417(.a(s_37), .O(gate28inter4));
  nand2 gate418(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate419(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate420(.a(N146), .O(gate28inter7));
  inv1  gate421(.a(N95), .O(gate28inter8));
  nand2 gate422(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate423(.a(s_37), .b(gate28inter3), .O(gate28inter10));
  nor2  gate424(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate425(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate426(.a(gate28inter12), .b(gate28inter1), .O(N177));
nand2 gate29( .a(N150), .b(N108), .O(N180) );

  xor2  gate735(.a(N123), .b(N21), .O(gate30inter0));
  nand2 gate736(.a(gate30inter0), .b(s_82), .O(gate30inter1));
  and2  gate737(.a(N123), .b(N21), .O(gate30inter2));
  inv1  gate738(.a(s_82), .O(gate30inter3));
  inv1  gate739(.a(s_83), .O(gate30inter4));
  nand2 gate740(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate741(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate742(.a(N21), .O(gate30inter7));
  inv1  gate743(.a(N123), .O(gate30inter8));
  nand2 gate744(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate745(.a(s_83), .b(gate30inter3), .O(gate30inter10));
  nor2  gate746(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate747(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate748(.a(gate30inter12), .b(gate30inter1), .O(N183));

  xor2  gate273(.a(N123), .b(N27), .O(gate31inter0));
  nand2 gate274(.a(gate31inter0), .b(s_16), .O(gate31inter1));
  and2  gate275(.a(N123), .b(N27), .O(gate31inter2));
  inv1  gate276(.a(s_16), .O(gate31inter3));
  inv1  gate277(.a(s_17), .O(gate31inter4));
  nand2 gate278(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate279(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate280(.a(N27), .O(gate31inter7));
  inv1  gate281(.a(N123), .O(gate31inter8));
  nand2 gate282(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate283(.a(s_17), .b(gate31inter3), .O(gate31inter10));
  nor2  gate284(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate285(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate286(.a(gate31inter12), .b(gate31inter1), .O(N184));
nor2 gate32( .a(N34), .b(N127), .O(N185) );
nor2 gate33( .a(N40), .b(N127), .O(N186) );

  xor2  gate623(.a(N131), .b(N47), .O(gate34inter0));
  nand2 gate624(.a(gate34inter0), .b(s_66), .O(gate34inter1));
  and2  gate625(.a(N131), .b(N47), .O(gate34inter2));
  inv1  gate626(.a(s_66), .O(gate34inter3));
  inv1  gate627(.a(s_67), .O(gate34inter4));
  nand2 gate628(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate629(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate630(.a(N47), .O(gate34inter7));
  inv1  gate631(.a(N131), .O(gate34inter8));
  nand2 gate632(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate633(.a(s_67), .b(gate34inter3), .O(gate34inter10));
  nor2  gate634(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate635(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate636(.a(gate34inter12), .b(gate34inter1), .O(N187));

  xor2  gate791(.a(N131), .b(N53), .O(gate35inter0));
  nand2 gate792(.a(gate35inter0), .b(s_90), .O(gate35inter1));
  and2  gate793(.a(N131), .b(N53), .O(gate35inter2));
  inv1  gate794(.a(s_90), .O(gate35inter3));
  inv1  gate795(.a(s_91), .O(gate35inter4));
  nand2 gate796(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate797(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate798(.a(N53), .O(gate35inter7));
  inv1  gate799(.a(N131), .O(gate35inter8));
  nand2 gate800(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate801(.a(s_91), .b(gate35inter3), .O(gate35inter10));
  nor2  gate802(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate803(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate804(.a(gate35inter12), .b(gate35inter1), .O(N188));
nor2 gate36( .a(N60), .b(N135), .O(N189) );

  xor2  gate357(.a(N135), .b(N66), .O(gate37inter0));
  nand2 gate358(.a(gate37inter0), .b(s_28), .O(gate37inter1));
  and2  gate359(.a(N135), .b(N66), .O(gate37inter2));
  inv1  gate360(.a(s_28), .O(gate37inter3));
  inv1  gate361(.a(s_29), .O(gate37inter4));
  nand2 gate362(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate363(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate364(.a(N66), .O(gate37inter7));
  inv1  gate365(.a(N135), .O(gate37inter8));
  nand2 gate366(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate367(.a(s_29), .b(gate37inter3), .O(gate37inter10));
  nor2  gate368(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate369(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate370(.a(gate37inter12), .b(gate37inter1), .O(N190));

  xor2  gate329(.a(N139), .b(N73), .O(gate38inter0));
  nand2 gate330(.a(gate38inter0), .b(s_24), .O(gate38inter1));
  and2  gate331(.a(N139), .b(N73), .O(gate38inter2));
  inv1  gate332(.a(s_24), .O(gate38inter3));
  inv1  gate333(.a(s_25), .O(gate38inter4));
  nand2 gate334(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate335(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate336(.a(N73), .O(gate38inter7));
  inv1  gate337(.a(N139), .O(gate38inter8));
  nand2 gate338(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate339(.a(s_25), .b(gate38inter3), .O(gate38inter10));
  nor2  gate340(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate341(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate342(.a(gate38inter12), .b(gate38inter1), .O(N191));

  xor2  gate595(.a(N139), .b(N79), .O(gate39inter0));
  nand2 gate596(.a(gate39inter0), .b(s_62), .O(gate39inter1));
  and2  gate597(.a(N139), .b(N79), .O(gate39inter2));
  inv1  gate598(.a(s_62), .O(gate39inter3));
  inv1  gate599(.a(s_63), .O(gate39inter4));
  nand2 gate600(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate601(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate602(.a(N79), .O(gate39inter7));
  inv1  gate603(.a(N139), .O(gate39inter8));
  nand2 gate604(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate605(.a(s_63), .b(gate39inter3), .O(gate39inter10));
  nor2  gate606(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate607(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate608(.a(gate39inter12), .b(gate39inter1), .O(N192));

  xor2  gate693(.a(N143), .b(N86), .O(gate40inter0));
  nand2 gate694(.a(gate40inter0), .b(s_76), .O(gate40inter1));
  and2  gate695(.a(N143), .b(N86), .O(gate40inter2));
  inv1  gate696(.a(s_76), .O(gate40inter3));
  inv1  gate697(.a(s_77), .O(gate40inter4));
  nand2 gate698(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate699(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate700(.a(N86), .O(gate40inter7));
  inv1  gate701(.a(N143), .O(gate40inter8));
  nand2 gate702(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate703(.a(s_77), .b(gate40inter3), .O(gate40inter10));
  nor2  gate704(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate705(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate706(.a(gate40inter12), .b(gate40inter1), .O(N193));

  xor2  gate371(.a(N143), .b(N92), .O(gate41inter0));
  nand2 gate372(.a(gate41inter0), .b(s_30), .O(gate41inter1));
  and2  gate373(.a(N143), .b(N92), .O(gate41inter2));
  inv1  gate374(.a(s_30), .O(gate41inter3));
  inv1  gate375(.a(s_31), .O(gate41inter4));
  nand2 gate376(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate377(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate378(.a(N92), .O(gate41inter7));
  inv1  gate379(.a(N143), .O(gate41inter8));
  nand2 gate380(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate381(.a(s_31), .b(gate41inter3), .O(gate41inter10));
  nor2  gate382(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate383(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate384(.a(gate41inter12), .b(gate41inter1), .O(N194));
nor2 gate42( .a(N99), .b(N147), .O(N195) );
nor2 gate43( .a(N105), .b(N147), .O(N196) );
nor2 gate44( .a(N112), .b(N151), .O(N197) );
nor2 gate45( .a(N115), .b(N151), .O(N198) );
and9 gate46( .a(N154), .b(N159), .c(N162), .d(N165), .e(N168), .f(N171), .g(N174), .h(N177), .i(N180), .O(N199) );
inv1 gate47( .a(N199), .O(N203) );
inv1 gate48( .a(N199), .O(N213) );
inv1 gate49( .a(N199), .O(N223) );
xor2 gate50( .a(N203), .b(N154), .O(N224) );
xor2 gate51( .a(N203), .b(N159), .O(N227) );

  xor2  gate763(.a(N162), .b(N203), .O(gate52inter0));
  nand2 gate764(.a(gate52inter0), .b(s_86), .O(gate52inter1));
  and2  gate765(.a(N162), .b(N203), .O(gate52inter2));
  inv1  gate766(.a(s_86), .O(gate52inter3));
  inv1  gate767(.a(s_87), .O(gate52inter4));
  nand2 gate768(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate769(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate770(.a(N203), .O(gate52inter7));
  inv1  gate771(.a(N162), .O(gate52inter8));
  nand2 gate772(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate773(.a(s_87), .b(gate52inter3), .O(gate52inter10));
  nor2  gate774(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate775(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate776(.a(gate52inter12), .b(gate52inter1), .O(N230));

  xor2  gate637(.a(N165), .b(N203), .O(gate53inter0));
  nand2 gate638(.a(gate53inter0), .b(s_68), .O(gate53inter1));
  and2  gate639(.a(N165), .b(N203), .O(gate53inter2));
  inv1  gate640(.a(s_68), .O(gate53inter3));
  inv1  gate641(.a(s_69), .O(gate53inter4));
  nand2 gate642(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate643(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate644(.a(N203), .O(gate53inter7));
  inv1  gate645(.a(N165), .O(gate53inter8));
  nand2 gate646(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate647(.a(s_69), .b(gate53inter3), .O(gate53inter10));
  nor2  gate648(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate649(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate650(.a(gate53inter12), .b(gate53inter1), .O(N233));
xor2 gate54( .a(N203), .b(N168), .O(N236) );
xor2 gate55( .a(N203), .b(N171), .O(N239) );
nand2 gate56( .a(N1), .b(N213), .O(N242) );
xor2 gate57( .a(N203), .b(N174), .O(N243) );
nand2 gate58( .a(N213), .b(N11), .O(N246) );
xor2 gate59( .a(N203), .b(N177), .O(N247) );

  xor2  gate231(.a(N24), .b(N213), .O(gate60inter0));
  nand2 gate232(.a(gate60inter0), .b(s_10), .O(gate60inter1));
  and2  gate233(.a(N24), .b(N213), .O(gate60inter2));
  inv1  gate234(.a(s_10), .O(gate60inter3));
  inv1  gate235(.a(s_11), .O(gate60inter4));
  nand2 gate236(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate237(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate238(.a(N213), .O(gate60inter7));
  inv1  gate239(.a(N24), .O(gate60inter8));
  nand2 gate240(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate241(.a(s_11), .b(gate60inter3), .O(gate60inter10));
  nor2  gate242(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate243(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate244(.a(gate60inter12), .b(gate60inter1), .O(N250));

  xor2  gate427(.a(N180), .b(N203), .O(gate61inter0));
  nand2 gate428(.a(gate61inter0), .b(s_38), .O(gate61inter1));
  and2  gate429(.a(N180), .b(N203), .O(gate61inter2));
  inv1  gate430(.a(s_38), .O(gate61inter3));
  inv1  gate431(.a(s_39), .O(gate61inter4));
  nand2 gate432(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate433(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate434(.a(N203), .O(gate61inter7));
  inv1  gate435(.a(N180), .O(gate61inter8));
  nand2 gate436(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate437(.a(s_39), .b(gate61inter3), .O(gate61inter10));
  nor2  gate438(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate439(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate440(.a(gate61inter12), .b(gate61inter1), .O(N251));
nand2 gate62( .a(N213), .b(N37), .O(N254) );
nand2 gate63( .a(N213), .b(N50), .O(N255) );

  xor2  gate525(.a(N63), .b(N213), .O(gate64inter0));
  nand2 gate526(.a(gate64inter0), .b(s_52), .O(gate64inter1));
  and2  gate527(.a(N63), .b(N213), .O(gate64inter2));
  inv1  gate528(.a(s_52), .O(gate64inter3));
  inv1  gate529(.a(s_53), .O(gate64inter4));
  nand2 gate530(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate531(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate532(.a(N213), .O(gate64inter7));
  inv1  gate533(.a(N63), .O(gate64inter8));
  nand2 gate534(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate535(.a(s_53), .b(gate64inter3), .O(gate64inter10));
  nor2  gate536(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate537(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate538(.a(gate64inter12), .b(gate64inter1), .O(N256));
nand2 gate65( .a(N213), .b(N76), .O(N257) );

  xor2  gate189(.a(N89), .b(N213), .O(gate66inter0));
  nand2 gate190(.a(gate66inter0), .b(s_4), .O(gate66inter1));
  and2  gate191(.a(N89), .b(N213), .O(gate66inter2));
  inv1  gate192(.a(s_4), .O(gate66inter3));
  inv1  gate193(.a(s_5), .O(gate66inter4));
  nand2 gate194(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate195(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate196(.a(N213), .O(gate66inter7));
  inv1  gate197(.a(N89), .O(gate66inter8));
  nand2 gate198(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate199(.a(s_5), .b(gate66inter3), .O(gate66inter10));
  nor2  gate200(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate201(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate202(.a(gate66inter12), .b(gate66inter1), .O(N258));
nand2 gate67( .a(N213), .b(N102), .O(N259) );

  xor2  gate217(.a(N157), .b(N224), .O(gate68inter0));
  nand2 gate218(.a(gate68inter0), .b(s_8), .O(gate68inter1));
  and2  gate219(.a(N157), .b(N224), .O(gate68inter2));
  inv1  gate220(.a(s_8), .O(gate68inter3));
  inv1  gate221(.a(s_9), .O(gate68inter4));
  nand2 gate222(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate223(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate224(.a(N224), .O(gate68inter7));
  inv1  gate225(.a(N157), .O(gate68inter8));
  nand2 gate226(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate227(.a(s_9), .b(gate68inter3), .O(gate68inter10));
  nor2  gate228(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate229(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate230(.a(gate68inter12), .b(gate68inter1), .O(N260));
nand2 gate69( .a(N224), .b(N158), .O(N263) );

  xor2  gate651(.a(N183), .b(N227), .O(gate70inter0));
  nand2 gate652(.a(gate70inter0), .b(s_70), .O(gate70inter1));
  and2  gate653(.a(N183), .b(N227), .O(gate70inter2));
  inv1  gate654(.a(s_70), .O(gate70inter3));
  inv1  gate655(.a(s_71), .O(gate70inter4));
  nand2 gate656(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate657(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate658(.a(N227), .O(gate70inter7));
  inv1  gate659(.a(N183), .O(gate70inter8));
  nand2 gate660(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate661(.a(s_71), .b(gate70inter3), .O(gate70inter10));
  nor2  gate662(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate663(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate664(.a(gate70inter12), .b(gate70inter1), .O(N264));

  xor2  gate707(.a(N185), .b(N230), .O(gate71inter0));
  nand2 gate708(.a(gate71inter0), .b(s_78), .O(gate71inter1));
  and2  gate709(.a(N185), .b(N230), .O(gate71inter2));
  inv1  gate710(.a(s_78), .O(gate71inter3));
  inv1  gate711(.a(s_79), .O(gate71inter4));
  nand2 gate712(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate713(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate714(.a(N230), .O(gate71inter7));
  inv1  gate715(.a(N185), .O(gate71inter8));
  nand2 gate716(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate717(.a(s_79), .b(gate71inter3), .O(gate71inter10));
  nor2  gate718(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate719(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate720(.a(gate71inter12), .b(gate71inter1), .O(N267));
nand2 gate72( .a(N233), .b(N187), .O(N270) );

  xor2  gate553(.a(N189), .b(N236), .O(gate73inter0));
  nand2 gate554(.a(gate73inter0), .b(s_56), .O(gate73inter1));
  and2  gate555(.a(N189), .b(N236), .O(gate73inter2));
  inv1  gate556(.a(s_56), .O(gate73inter3));
  inv1  gate557(.a(s_57), .O(gate73inter4));
  nand2 gate558(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate559(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate560(.a(N236), .O(gate73inter7));
  inv1  gate561(.a(N189), .O(gate73inter8));
  nand2 gate562(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate563(.a(s_57), .b(gate73inter3), .O(gate73inter10));
  nor2  gate564(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate565(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate566(.a(gate73inter12), .b(gate73inter1), .O(N273));
nand2 gate74( .a(N239), .b(N191), .O(N276) );

  xor2  gate567(.a(N193), .b(N243), .O(gate75inter0));
  nand2 gate568(.a(gate75inter0), .b(s_58), .O(gate75inter1));
  and2  gate569(.a(N193), .b(N243), .O(gate75inter2));
  inv1  gate570(.a(s_58), .O(gate75inter3));
  inv1  gate571(.a(s_59), .O(gate75inter4));
  nand2 gate572(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate573(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate574(.a(N243), .O(gate75inter7));
  inv1  gate575(.a(N193), .O(gate75inter8));
  nand2 gate576(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate577(.a(s_59), .b(gate75inter3), .O(gate75inter10));
  nor2  gate578(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate579(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate580(.a(gate75inter12), .b(gate75inter1), .O(N279));
nand2 gate76( .a(N247), .b(N195), .O(N282) );

  xor2  gate511(.a(N197), .b(N251), .O(gate77inter0));
  nand2 gate512(.a(gate77inter0), .b(s_50), .O(gate77inter1));
  and2  gate513(.a(N197), .b(N251), .O(gate77inter2));
  inv1  gate514(.a(s_50), .O(gate77inter3));
  inv1  gate515(.a(s_51), .O(gate77inter4));
  nand2 gate516(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate517(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate518(.a(N251), .O(gate77inter7));
  inv1  gate519(.a(N197), .O(gate77inter8));
  nand2 gate520(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate521(.a(s_51), .b(gate77inter3), .O(gate77inter10));
  nor2  gate522(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate523(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate524(.a(gate77inter12), .b(gate77inter1), .O(N285));
nand2 gate78( .a(N227), .b(N184), .O(N288) );

  xor2  gate679(.a(N186), .b(N230), .O(gate79inter0));
  nand2 gate680(.a(gate79inter0), .b(s_74), .O(gate79inter1));
  and2  gate681(.a(N186), .b(N230), .O(gate79inter2));
  inv1  gate682(.a(s_74), .O(gate79inter3));
  inv1  gate683(.a(s_75), .O(gate79inter4));
  nand2 gate684(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate685(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate686(.a(N230), .O(gate79inter7));
  inv1  gate687(.a(N186), .O(gate79inter8));
  nand2 gate688(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate689(.a(s_75), .b(gate79inter3), .O(gate79inter10));
  nor2  gate690(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate691(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate692(.a(gate79inter12), .b(gate79inter1), .O(N289));

  xor2  gate175(.a(N188), .b(N233), .O(gate80inter0));
  nand2 gate176(.a(gate80inter0), .b(s_2), .O(gate80inter1));
  and2  gate177(.a(N188), .b(N233), .O(gate80inter2));
  inv1  gate178(.a(s_2), .O(gate80inter3));
  inv1  gate179(.a(s_3), .O(gate80inter4));
  nand2 gate180(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate181(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate182(.a(N233), .O(gate80inter7));
  inv1  gate183(.a(N188), .O(gate80inter8));
  nand2 gate184(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate185(.a(s_3), .b(gate80inter3), .O(gate80inter10));
  nor2  gate186(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate187(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate188(.a(gate80inter12), .b(gate80inter1), .O(N290));
nand2 gate81( .a(N236), .b(N190), .O(N291) );
nand2 gate82( .a(N239), .b(N192), .O(N292) );
nand2 gate83( .a(N243), .b(N194), .O(N293) );

  xor2  gate245(.a(N196), .b(N247), .O(gate84inter0));
  nand2 gate246(.a(gate84inter0), .b(s_12), .O(gate84inter1));
  and2  gate247(.a(N196), .b(N247), .O(gate84inter2));
  inv1  gate248(.a(s_12), .O(gate84inter3));
  inv1  gate249(.a(s_13), .O(gate84inter4));
  nand2 gate250(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate251(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate252(.a(N247), .O(gate84inter7));
  inv1  gate253(.a(N196), .O(gate84inter8));
  nand2 gate254(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate255(.a(s_13), .b(gate84inter3), .O(gate84inter10));
  nor2  gate256(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate257(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate258(.a(gate84inter12), .b(gate84inter1), .O(N294));

  xor2  gate287(.a(N198), .b(N251), .O(gate85inter0));
  nand2 gate288(.a(gate85inter0), .b(s_18), .O(gate85inter1));
  and2  gate289(.a(N198), .b(N251), .O(gate85inter2));
  inv1  gate290(.a(s_18), .O(gate85inter3));
  inv1  gate291(.a(s_19), .O(gate85inter4));
  nand2 gate292(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate293(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate294(.a(N251), .O(gate85inter7));
  inv1  gate295(.a(N198), .O(gate85inter8));
  nand2 gate296(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate297(.a(s_19), .b(gate85inter3), .O(gate85inter10));
  nor2  gate298(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate299(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate300(.a(gate85inter12), .b(gate85inter1), .O(N295));
and9 gate86( .a(N260), .b(N264), .c(N267), .d(N270), .e(N273), .f(N276), .g(N279), .h(N282), .i(N285), .O(N296) );
inv1 gate87( .a(N263), .O(N300) );
inv1 gate88( .a(N288), .O(N301) );
inv1 gate89( .a(N289), .O(N302) );
inv1 gate90( .a(N290), .O(N303) );
inv1 gate91( .a(N291), .O(N304) );
inv1 gate92( .a(N292), .O(N305) );
inv1 gate93( .a(N293), .O(N306) );
inv1 gate94( .a(N294), .O(N307) );
inv1 gate95( .a(N295), .O(N308) );
inv1 gate96( .a(N296), .O(N309) );
inv1 gate97( .a(N296), .O(N319) );
inv1 gate98( .a(N296), .O(N329) );

  xor2  gate721(.a(N260), .b(N309), .O(gate99inter0));
  nand2 gate722(.a(gate99inter0), .b(s_80), .O(gate99inter1));
  and2  gate723(.a(N260), .b(N309), .O(gate99inter2));
  inv1  gate724(.a(s_80), .O(gate99inter3));
  inv1  gate725(.a(s_81), .O(gate99inter4));
  nand2 gate726(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate727(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate728(.a(N309), .O(gate99inter7));
  inv1  gate729(.a(N260), .O(gate99inter8));
  nand2 gate730(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate731(.a(s_81), .b(gate99inter3), .O(gate99inter10));
  nor2  gate732(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate733(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate734(.a(gate99inter12), .b(gate99inter1), .O(N330));
xor2 gate100( .a(N309), .b(N264), .O(N331) );

  xor2  gate777(.a(N267), .b(N309), .O(gate101inter0));
  nand2 gate778(.a(gate101inter0), .b(s_88), .O(gate101inter1));
  and2  gate779(.a(N267), .b(N309), .O(gate101inter2));
  inv1  gate780(.a(s_88), .O(gate101inter3));
  inv1  gate781(.a(s_89), .O(gate101inter4));
  nand2 gate782(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate783(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate784(.a(N309), .O(gate101inter7));
  inv1  gate785(.a(N267), .O(gate101inter8));
  nand2 gate786(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate787(.a(s_89), .b(gate101inter3), .O(gate101inter10));
  nor2  gate788(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate789(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate790(.a(gate101inter12), .b(gate101inter1), .O(N332));

  xor2  gate665(.a(N270), .b(N309), .O(gate102inter0));
  nand2 gate666(.a(gate102inter0), .b(s_72), .O(gate102inter1));
  and2  gate667(.a(N270), .b(N309), .O(gate102inter2));
  inv1  gate668(.a(s_72), .O(gate102inter3));
  inv1  gate669(.a(s_73), .O(gate102inter4));
  nand2 gate670(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate671(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate672(.a(N309), .O(gate102inter7));
  inv1  gate673(.a(N270), .O(gate102inter8));
  nand2 gate674(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate675(.a(s_73), .b(gate102inter3), .O(gate102inter10));
  nor2  gate676(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate677(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate678(.a(gate102inter12), .b(gate102inter1), .O(N333));

  xor2  gate203(.a(N319), .b(N8), .O(gate103inter0));
  nand2 gate204(.a(gate103inter0), .b(s_6), .O(gate103inter1));
  and2  gate205(.a(N319), .b(N8), .O(gate103inter2));
  inv1  gate206(.a(s_6), .O(gate103inter3));
  inv1  gate207(.a(s_7), .O(gate103inter4));
  nand2 gate208(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate209(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate210(.a(N8), .O(gate103inter7));
  inv1  gate211(.a(N319), .O(gate103inter8));
  nand2 gate212(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate213(.a(s_7), .b(gate103inter3), .O(gate103inter10));
  nor2  gate214(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate215(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate216(.a(gate103inter12), .b(gate103inter1), .O(N334));
xor2 gate104( .a(N309), .b(N273), .O(N335) );
nand2 gate105( .a(N319), .b(N21), .O(N336) );
xor2 gate106( .a(N309), .b(N276), .O(N337) );
nand2 gate107( .a(N319), .b(N34), .O(N338) );

  xor2  gate161(.a(N279), .b(N309), .O(gate108inter0));
  nand2 gate162(.a(gate108inter0), .b(s_0), .O(gate108inter1));
  and2  gate163(.a(N279), .b(N309), .O(gate108inter2));
  inv1  gate164(.a(s_0), .O(gate108inter3));
  inv1  gate165(.a(s_1), .O(gate108inter4));
  nand2 gate166(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate167(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate168(.a(N309), .O(gate108inter7));
  inv1  gate169(.a(N279), .O(gate108inter8));
  nand2 gate170(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate171(.a(s_1), .b(gate108inter3), .O(gate108inter10));
  nor2  gate172(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate173(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate174(.a(gate108inter12), .b(gate108inter1), .O(N339));

  xor2  gate749(.a(N47), .b(N319), .O(gate109inter0));
  nand2 gate750(.a(gate109inter0), .b(s_84), .O(gate109inter1));
  and2  gate751(.a(N47), .b(N319), .O(gate109inter2));
  inv1  gate752(.a(s_84), .O(gate109inter3));
  inv1  gate753(.a(s_85), .O(gate109inter4));
  nand2 gate754(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate755(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate756(.a(N319), .O(gate109inter7));
  inv1  gate757(.a(N47), .O(gate109inter8));
  nand2 gate758(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate759(.a(s_85), .b(gate109inter3), .O(gate109inter10));
  nor2  gate760(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate761(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate762(.a(gate109inter12), .b(gate109inter1), .O(N340));
xor2 gate110( .a(N309), .b(N282), .O(N341) );
nand2 gate111( .a(N319), .b(N60), .O(N342) );
xor2 gate112( .a(N309), .b(N285), .O(N343) );
nand2 gate113( .a(N319), .b(N73), .O(N344) );
nand2 gate114( .a(N319), .b(N86), .O(N345) );

  xor2  gate609(.a(N99), .b(N319), .O(gate115inter0));
  nand2 gate610(.a(gate115inter0), .b(s_64), .O(gate115inter1));
  and2  gate611(.a(N99), .b(N319), .O(gate115inter2));
  inv1  gate612(.a(s_64), .O(gate115inter3));
  inv1  gate613(.a(s_65), .O(gate115inter4));
  nand2 gate614(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate615(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate616(.a(N319), .O(gate115inter7));
  inv1  gate617(.a(N99), .O(gate115inter8));
  nand2 gate618(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate619(.a(s_65), .b(gate115inter3), .O(gate115inter10));
  nor2  gate620(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate621(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate622(.a(gate115inter12), .b(gate115inter1), .O(N346));

  xor2  gate581(.a(N112), .b(N319), .O(gate116inter0));
  nand2 gate582(.a(gate116inter0), .b(s_60), .O(gate116inter1));
  and2  gate583(.a(N112), .b(N319), .O(gate116inter2));
  inv1  gate584(.a(s_60), .O(gate116inter3));
  inv1  gate585(.a(s_61), .O(gate116inter4));
  nand2 gate586(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate587(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate588(.a(N319), .O(gate116inter7));
  inv1  gate589(.a(N112), .O(gate116inter8));
  nand2 gate590(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate591(.a(s_61), .b(gate116inter3), .O(gate116inter10));
  nor2  gate592(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate593(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate594(.a(gate116inter12), .b(gate116inter1), .O(N347));
nand2 gate117( .a(N330), .b(N300), .O(N348) );

  xor2  gate399(.a(N301), .b(N331), .O(gate118inter0));
  nand2 gate400(.a(gate118inter0), .b(s_34), .O(gate118inter1));
  and2  gate401(.a(N301), .b(N331), .O(gate118inter2));
  inv1  gate402(.a(s_34), .O(gate118inter3));
  inv1  gate403(.a(s_35), .O(gate118inter4));
  nand2 gate404(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate405(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate406(.a(N331), .O(gate118inter7));
  inv1  gate407(.a(N301), .O(gate118inter8));
  nand2 gate408(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate409(.a(s_35), .b(gate118inter3), .O(gate118inter10));
  nor2  gate410(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate411(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate412(.a(gate118inter12), .b(gate118inter1), .O(N349));
nand2 gate119( .a(N332), .b(N302), .O(N350) );
nand2 gate120( .a(N333), .b(N303), .O(N351) );

  xor2  gate315(.a(N304), .b(N335), .O(gate121inter0));
  nand2 gate316(.a(gate121inter0), .b(s_22), .O(gate121inter1));
  and2  gate317(.a(N304), .b(N335), .O(gate121inter2));
  inv1  gate318(.a(s_22), .O(gate121inter3));
  inv1  gate319(.a(s_23), .O(gate121inter4));
  nand2 gate320(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate321(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate322(.a(N335), .O(gate121inter7));
  inv1  gate323(.a(N304), .O(gate121inter8));
  nand2 gate324(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate325(.a(s_23), .b(gate121inter3), .O(gate121inter10));
  nor2  gate326(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate327(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate328(.a(gate121inter12), .b(gate121inter1), .O(N352));
nand2 gate122( .a(N337), .b(N305), .O(N353) );
nand2 gate123( .a(N339), .b(N306), .O(N354) );

  xor2  gate343(.a(N307), .b(N341), .O(gate124inter0));
  nand2 gate344(.a(gate124inter0), .b(s_26), .O(gate124inter1));
  and2  gate345(.a(N307), .b(N341), .O(gate124inter2));
  inv1  gate346(.a(s_26), .O(gate124inter3));
  inv1  gate347(.a(s_27), .O(gate124inter4));
  nand2 gate348(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate349(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate350(.a(N341), .O(gate124inter7));
  inv1  gate351(.a(N307), .O(gate124inter8));
  nand2 gate352(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate353(.a(s_27), .b(gate124inter3), .O(gate124inter10));
  nor2  gate354(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate355(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate356(.a(gate124inter12), .b(gate124inter1), .O(N355));

  xor2  gate539(.a(N308), .b(N343), .O(gate125inter0));
  nand2 gate540(.a(gate125inter0), .b(s_54), .O(gate125inter1));
  and2  gate541(.a(N308), .b(N343), .O(gate125inter2));
  inv1  gate542(.a(s_54), .O(gate125inter3));
  inv1  gate543(.a(s_55), .O(gate125inter4));
  nand2 gate544(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate545(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate546(.a(N343), .O(gate125inter7));
  inv1  gate547(.a(N308), .O(gate125inter8));
  nand2 gate548(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate549(.a(s_55), .b(gate125inter3), .O(gate125inter10));
  nor2  gate550(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate551(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate552(.a(gate125inter12), .b(gate125inter1), .O(N356));
and9 gate126( .a(N348), .b(N349), .c(N350), .d(N351), .e(N352), .f(N353), .g(N354), .h(N355), .i(N356), .O(N357) );
inv1 gate127( .a(N357), .O(N360) );
inv1 gate128( .a(N357), .O(N370) );
nand2 gate129( .a(N14), .b(N360), .O(N371) );
nand2 gate130( .a(N360), .b(N27), .O(N372) );
nand2 gate131( .a(N360), .b(N40), .O(N373) );

  xor2  gate469(.a(N53), .b(N360), .O(gate132inter0));
  nand2 gate470(.a(gate132inter0), .b(s_44), .O(gate132inter1));
  and2  gate471(.a(N53), .b(N360), .O(gate132inter2));
  inv1  gate472(.a(s_44), .O(gate132inter3));
  inv1  gate473(.a(s_45), .O(gate132inter4));
  nand2 gate474(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate475(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate476(.a(N360), .O(gate132inter7));
  inv1  gate477(.a(N53), .O(gate132inter8));
  nand2 gate478(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate479(.a(s_45), .b(gate132inter3), .O(gate132inter10));
  nor2  gate480(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate481(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate482(.a(gate132inter12), .b(gate132inter1), .O(N374));
nand2 gate133( .a(N360), .b(N66), .O(N375) );
nand2 gate134( .a(N360), .b(N79), .O(N376) );

  xor2  gate483(.a(N92), .b(N360), .O(gate135inter0));
  nand2 gate484(.a(gate135inter0), .b(s_46), .O(gate135inter1));
  and2  gate485(.a(N92), .b(N360), .O(gate135inter2));
  inv1  gate486(.a(s_46), .O(gate135inter3));
  inv1  gate487(.a(s_47), .O(gate135inter4));
  nand2 gate488(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate489(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate490(.a(N360), .O(gate135inter7));
  inv1  gate491(.a(N92), .O(gate135inter8));
  nand2 gate492(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate493(.a(s_47), .b(gate135inter3), .O(gate135inter10));
  nor2  gate494(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate495(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate496(.a(gate135inter12), .b(gate135inter1), .O(N377));
nand2 gate136( .a(N360), .b(N105), .O(N378) );

  xor2  gate441(.a(N115), .b(N360), .O(gate137inter0));
  nand2 gate442(.a(gate137inter0), .b(s_40), .O(gate137inter1));
  and2  gate443(.a(N115), .b(N360), .O(gate137inter2));
  inv1  gate444(.a(s_40), .O(gate137inter3));
  inv1  gate445(.a(s_41), .O(gate137inter4));
  nand2 gate446(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate447(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate448(.a(N360), .O(gate137inter7));
  inv1  gate449(.a(N115), .O(gate137inter8));
  nand2 gate450(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate451(.a(s_41), .b(gate137inter3), .O(gate137inter10));
  nor2  gate452(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate453(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate454(.a(gate137inter12), .b(gate137inter1), .O(N379));
nand4 gate138( .a(N4), .b(N242), .c(N334), .d(N371), .O(N380) );
nand4 gate139( .a(N246), .b(N336), .c(N372), .d(N17), .O(N381) );
nand4 gate140( .a(N250), .b(N338), .c(N373), .d(N30), .O(N386) );
nand4 gate141( .a(N254), .b(N340), .c(N374), .d(N43), .O(N393) );
nand4 gate142( .a(N255), .b(N342), .c(N375), .d(N56), .O(N399) );
nand4 gate143( .a(N256), .b(N344), .c(N376), .d(N69), .O(N404) );
nand4 gate144( .a(N257), .b(N345), .c(N377), .d(N82), .O(N407) );
nand4 gate145( .a(N258), .b(N346), .c(N378), .d(N95), .O(N411) );
nand4 gate146( .a(N259), .b(N347), .c(N379), .d(N108), .O(N414) );
inv1 gate147( .a(N380), .O(N415) );
and8 gate148( .a(N381), .b(N386), .c(N393), .d(N399), .e(N404), .f(N407), .g(N411), .h(N414), .O(N416) );
inv1 gate149( .a(N393), .O(N417) );
inv1 gate150( .a(N404), .O(N418) );
inv1 gate151( .a(N407), .O(N419) );
inv1 gate152( .a(N411), .O(N420) );

  xor2  gate497(.a(N416), .b(N415), .O(gate153inter0));
  nand2 gate498(.a(gate153inter0), .b(s_48), .O(gate153inter1));
  and2  gate499(.a(N416), .b(N415), .O(gate153inter2));
  inv1  gate500(.a(s_48), .O(gate153inter3));
  inv1  gate501(.a(s_49), .O(gate153inter4));
  nand2 gate502(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate503(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate504(.a(N415), .O(gate153inter7));
  inv1  gate505(.a(N416), .O(gate153inter8));
  nand2 gate506(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate507(.a(s_49), .b(gate153inter3), .O(gate153inter10));
  nor2  gate508(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate509(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate510(.a(gate153inter12), .b(gate153inter1), .O(N421));

  xor2  gate455(.a(N417), .b(N386), .O(gate154inter0));
  nand2 gate456(.a(gate154inter0), .b(s_42), .O(gate154inter1));
  and2  gate457(.a(N417), .b(N386), .O(gate154inter2));
  inv1  gate458(.a(s_42), .O(gate154inter3));
  inv1  gate459(.a(s_43), .O(gate154inter4));
  nand2 gate460(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate461(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate462(.a(N386), .O(gate154inter7));
  inv1  gate463(.a(N417), .O(gate154inter8));
  nand2 gate464(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate465(.a(s_43), .b(gate154inter3), .O(gate154inter10));
  nor2  gate466(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate467(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate468(.a(gate154inter12), .b(gate154inter1), .O(N422));
nand4 gate155( .a(N386), .b(N393), .c(N418), .d(N399), .O(N425) );
nand3 gate156( .a(N399), .b(N393), .c(N419), .O(N428) );
nand4 gate157( .a(N386), .b(N393), .c(N407), .d(N420), .O(N429) );
nand4 gate158( .a(N381), .b(N386), .c(N422), .d(N399), .O(N430) );
nand4 gate159( .a(N381), .b(N386), .c(N425), .d(N428), .O(N431) );
nand4 gate160( .a(N381), .b(N422), .c(N425), .d(N429), .O(N432) );

endmodule