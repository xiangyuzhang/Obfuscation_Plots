module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate813(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate814(.a(gate9inter0), .b(s_38), .O(gate9inter1));
  and2  gate815(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate816(.a(s_38), .O(gate9inter3));
  inv1  gate817(.a(s_39), .O(gate9inter4));
  nand2 gate818(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate819(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate820(.a(G1), .O(gate9inter7));
  inv1  gate821(.a(G2), .O(gate9inter8));
  nand2 gate822(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate823(.a(s_39), .b(gate9inter3), .O(gate9inter10));
  nor2  gate824(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate825(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate826(.a(gate9inter12), .b(gate9inter1), .O(G266));

  xor2  gate1471(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate1472(.a(gate10inter0), .b(s_132), .O(gate10inter1));
  and2  gate1473(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate1474(.a(s_132), .O(gate10inter3));
  inv1  gate1475(.a(s_133), .O(gate10inter4));
  nand2 gate1476(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate1477(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate1478(.a(G3), .O(gate10inter7));
  inv1  gate1479(.a(G4), .O(gate10inter8));
  nand2 gate1480(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate1481(.a(s_133), .b(gate10inter3), .O(gate10inter10));
  nor2  gate1482(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate1483(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate1484(.a(gate10inter12), .b(gate10inter1), .O(G269));
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );

  xor2  gate1415(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate1416(.a(gate14inter0), .b(s_124), .O(gate14inter1));
  and2  gate1417(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate1418(.a(s_124), .O(gate14inter3));
  inv1  gate1419(.a(s_125), .O(gate14inter4));
  nand2 gate1420(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate1421(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate1422(.a(G11), .O(gate14inter7));
  inv1  gate1423(.a(G12), .O(gate14inter8));
  nand2 gate1424(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate1425(.a(s_125), .b(gate14inter3), .O(gate14inter10));
  nor2  gate1426(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate1427(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate1428(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate743(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate744(.a(gate16inter0), .b(s_28), .O(gate16inter1));
  and2  gate745(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate746(.a(s_28), .O(gate16inter3));
  inv1  gate747(.a(s_29), .O(gate16inter4));
  nand2 gate748(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate749(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate750(.a(G15), .O(gate16inter7));
  inv1  gate751(.a(G16), .O(gate16inter8));
  nand2 gate752(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate753(.a(s_29), .b(gate16inter3), .O(gate16inter10));
  nor2  gate754(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate755(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate756(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate547(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate548(.a(gate27inter0), .b(s_0), .O(gate27inter1));
  and2  gate549(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate550(.a(s_0), .O(gate27inter3));
  inv1  gate551(.a(s_1), .O(gate27inter4));
  nand2 gate552(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate553(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate554(.a(G2), .O(gate27inter7));
  inv1  gate555(.a(G6), .O(gate27inter8));
  nand2 gate556(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate557(.a(s_1), .b(gate27inter3), .O(gate27inter10));
  nor2  gate558(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate559(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate560(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );

  xor2  gate841(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate842(.a(gate30inter0), .b(s_42), .O(gate30inter1));
  and2  gate843(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate844(.a(s_42), .O(gate30inter3));
  inv1  gate845(.a(s_43), .O(gate30inter4));
  nand2 gate846(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate847(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate848(.a(G11), .O(gate30inter7));
  inv1  gate849(.a(G15), .O(gate30inter8));
  nand2 gate850(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate851(.a(s_43), .b(gate30inter3), .O(gate30inter10));
  nor2  gate852(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate853(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate854(.a(gate30inter12), .b(gate30inter1), .O(G329));
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate771(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate772(.a(gate34inter0), .b(s_32), .O(gate34inter1));
  and2  gate773(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate774(.a(s_32), .O(gate34inter3));
  inv1  gate775(.a(s_33), .O(gate34inter4));
  nand2 gate776(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate777(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate778(.a(G25), .O(gate34inter7));
  inv1  gate779(.a(G29), .O(gate34inter8));
  nand2 gate780(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate781(.a(s_33), .b(gate34inter3), .O(gate34inter10));
  nor2  gate782(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate783(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate784(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate1485(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1486(.a(gate36inter0), .b(s_134), .O(gate36inter1));
  and2  gate1487(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1488(.a(s_134), .O(gate36inter3));
  inv1  gate1489(.a(s_135), .O(gate36inter4));
  nand2 gate1490(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1491(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1492(.a(G26), .O(gate36inter7));
  inv1  gate1493(.a(G30), .O(gate36inter8));
  nand2 gate1494(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1495(.a(s_135), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1496(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1497(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1498(.a(gate36inter12), .b(gate36inter1), .O(G347));

  xor2  gate575(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate576(.a(gate37inter0), .b(s_4), .O(gate37inter1));
  and2  gate577(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate578(.a(s_4), .O(gate37inter3));
  inv1  gate579(.a(s_5), .O(gate37inter4));
  nand2 gate580(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate581(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate582(.a(G19), .O(gate37inter7));
  inv1  gate583(.a(G23), .O(gate37inter8));
  nand2 gate584(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate585(.a(s_5), .b(gate37inter3), .O(gate37inter10));
  nor2  gate586(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate587(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate588(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate1023(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate1024(.a(gate51inter0), .b(s_68), .O(gate51inter1));
  and2  gate1025(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate1026(.a(s_68), .O(gate51inter3));
  inv1  gate1027(.a(s_69), .O(gate51inter4));
  nand2 gate1028(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate1029(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate1030(.a(G11), .O(gate51inter7));
  inv1  gate1031(.a(G281), .O(gate51inter8));
  nand2 gate1032(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate1033(.a(s_69), .b(gate51inter3), .O(gate51inter10));
  nor2  gate1034(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate1035(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate1036(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );

  xor2  gate1457(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate1458(.a(gate61inter0), .b(s_130), .O(gate61inter1));
  and2  gate1459(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate1460(.a(s_130), .O(gate61inter3));
  inv1  gate1461(.a(s_131), .O(gate61inter4));
  nand2 gate1462(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate1463(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate1464(.a(G21), .O(gate61inter7));
  inv1  gate1465(.a(G296), .O(gate61inter8));
  nand2 gate1466(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate1467(.a(s_131), .b(gate61inter3), .O(gate61inter10));
  nor2  gate1468(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate1469(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate1470(.a(gate61inter12), .b(gate61inter1), .O(G382));
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate925(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate926(.a(gate63inter0), .b(s_54), .O(gate63inter1));
  and2  gate927(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate928(.a(s_54), .O(gate63inter3));
  inv1  gate929(.a(s_55), .O(gate63inter4));
  nand2 gate930(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate931(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate932(.a(G23), .O(gate63inter7));
  inv1  gate933(.a(G299), .O(gate63inter8));
  nand2 gate934(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate935(.a(s_55), .b(gate63inter3), .O(gate63inter10));
  nor2  gate936(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate937(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate938(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate1345(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate1346(.a(gate69inter0), .b(s_114), .O(gate69inter1));
  and2  gate1347(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate1348(.a(s_114), .O(gate69inter3));
  inv1  gate1349(.a(s_115), .O(gate69inter4));
  nand2 gate1350(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate1351(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate1352(.a(G29), .O(gate69inter7));
  inv1  gate1353(.a(G308), .O(gate69inter8));
  nand2 gate1354(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate1355(.a(s_115), .b(gate69inter3), .O(gate69inter10));
  nor2  gate1356(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate1357(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate1358(.a(gate69inter12), .b(gate69inter1), .O(G390));
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );

  xor2  gate883(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate884(.a(gate84inter0), .b(s_48), .O(gate84inter1));
  and2  gate885(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate886(.a(s_48), .O(gate84inter3));
  inv1  gate887(.a(s_49), .O(gate84inter4));
  nand2 gate888(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate889(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate890(.a(G15), .O(gate84inter7));
  inv1  gate891(.a(G329), .O(gate84inter8));
  nand2 gate892(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate893(.a(s_49), .b(gate84inter3), .O(gate84inter10));
  nor2  gate894(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate895(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate896(.a(gate84inter12), .b(gate84inter1), .O(G405));
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate687(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate688(.a(gate91inter0), .b(s_20), .O(gate91inter1));
  and2  gate689(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate690(.a(s_20), .O(gate91inter3));
  inv1  gate691(.a(s_21), .O(gate91inter4));
  nand2 gate692(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate693(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate694(.a(G25), .O(gate91inter7));
  inv1  gate695(.a(G341), .O(gate91inter8));
  nand2 gate696(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate697(.a(s_21), .b(gate91inter3), .O(gate91inter10));
  nor2  gate698(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate699(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate700(.a(gate91inter12), .b(gate91inter1), .O(G412));

  xor2  gate1233(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate1234(.a(gate92inter0), .b(s_98), .O(gate92inter1));
  and2  gate1235(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate1236(.a(s_98), .O(gate92inter3));
  inv1  gate1237(.a(s_99), .O(gate92inter4));
  nand2 gate1238(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate1239(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate1240(.a(G29), .O(gate92inter7));
  inv1  gate1241(.a(G341), .O(gate92inter8));
  nand2 gate1242(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate1243(.a(s_99), .b(gate92inter3), .O(gate92inter10));
  nor2  gate1244(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate1245(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate1246(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate1065(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate1066(.a(gate95inter0), .b(s_74), .O(gate95inter1));
  and2  gate1067(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate1068(.a(s_74), .O(gate95inter3));
  inv1  gate1069(.a(s_75), .O(gate95inter4));
  nand2 gate1070(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate1071(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate1072(.a(G26), .O(gate95inter7));
  inv1  gate1073(.a(G347), .O(gate95inter8));
  nand2 gate1074(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate1075(.a(s_75), .b(gate95inter3), .O(gate95inter10));
  nor2  gate1076(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate1077(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate1078(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate1149(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate1150(.a(gate99inter0), .b(s_86), .O(gate99inter1));
  and2  gate1151(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate1152(.a(s_86), .O(gate99inter3));
  inv1  gate1153(.a(s_87), .O(gate99inter4));
  nand2 gate1154(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate1155(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate1156(.a(G27), .O(gate99inter7));
  inv1  gate1157(.a(G353), .O(gate99inter8));
  nand2 gate1158(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate1159(.a(s_87), .b(gate99inter3), .O(gate99inter10));
  nor2  gate1160(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate1161(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate1162(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );

  xor2  gate631(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate632(.a(gate101inter0), .b(s_12), .O(gate101inter1));
  and2  gate633(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate634(.a(s_12), .O(gate101inter3));
  inv1  gate635(.a(s_13), .O(gate101inter4));
  nand2 gate636(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate637(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate638(.a(G20), .O(gate101inter7));
  inv1  gate639(.a(G356), .O(gate101inter8));
  nand2 gate640(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate641(.a(s_13), .b(gate101inter3), .O(gate101inter10));
  nor2  gate642(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate643(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate644(.a(gate101inter12), .b(gate101inter1), .O(G422));
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate897(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate898(.a(gate106inter0), .b(s_50), .O(gate106inter1));
  and2  gate899(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate900(.a(s_50), .O(gate106inter3));
  inv1  gate901(.a(s_51), .O(gate106inter4));
  nand2 gate902(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate903(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate904(.a(G364), .O(gate106inter7));
  inv1  gate905(.a(G365), .O(gate106inter8));
  nand2 gate906(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate907(.a(s_51), .b(gate106inter3), .O(gate106inter10));
  nor2  gate908(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate909(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate910(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );

  xor2  gate1275(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate1276(.a(gate114inter0), .b(s_104), .O(gate114inter1));
  and2  gate1277(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate1278(.a(s_104), .O(gate114inter3));
  inv1  gate1279(.a(s_105), .O(gate114inter4));
  nand2 gate1280(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate1281(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate1282(.a(G380), .O(gate114inter7));
  inv1  gate1283(.a(G381), .O(gate114inter8));
  nand2 gate1284(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate1285(.a(s_105), .b(gate114inter3), .O(gate114inter10));
  nor2  gate1286(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate1287(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate1288(.a(gate114inter12), .b(gate114inter1), .O(G453));
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate953(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate954(.a(gate131inter0), .b(s_58), .O(gate131inter1));
  and2  gate955(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate956(.a(s_58), .O(gate131inter3));
  inv1  gate957(.a(s_59), .O(gate131inter4));
  nand2 gate958(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate959(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate960(.a(G414), .O(gate131inter7));
  inv1  gate961(.a(G415), .O(gate131inter8));
  nand2 gate962(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate963(.a(s_59), .b(gate131inter3), .O(gate131inter10));
  nor2  gate964(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate965(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate966(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate1289(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate1290(.a(gate137inter0), .b(s_106), .O(gate137inter1));
  and2  gate1291(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate1292(.a(s_106), .O(gate137inter3));
  inv1  gate1293(.a(s_107), .O(gate137inter4));
  nand2 gate1294(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate1295(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate1296(.a(G426), .O(gate137inter7));
  inv1  gate1297(.a(G429), .O(gate137inter8));
  nand2 gate1298(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate1299(.a(s_107), .b(gate137inter3), .O(gate137inter10));
  nor2  gate1300(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate1301(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate1302(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );

  xor2  gate995(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate996(.a(gate140inter0), .b(s_64), .O(gate140inter1));
  and2  gate997(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate998(.a(s_64), .O(gate140inter3));
  inv1  gate999(.a(s_65), .O(gate140inter4));
  nand2 gate1000(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate1001(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate1002(.a(G444), .O(gate140inter7));
  inv1  gate1003(.a(G447), .O(gate140inter8));
  nand2 gate1004(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate1005(.a(s_65), .b(gate140inter3), .O(gate140inter10));
  nor2  gate1006(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate1007(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate1008(.a(gate140inter12), .b(gate140inter1), .O(G531));
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate1009(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate1010(.a(gate153inter0), .b(s_66), .O(gate153inter1));
  and2  gate1011(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate1012(.a(s_66), .O(gate153inter3));
  inv1  gate1013(.a(s_67), .O(gate153inter4));
  nand2 gate1014(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate1015(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate1016(.a(G426), .O(gate153inter7));
  inv1  gate1017(.a(G522), .O(gate153inter8));
  nand2 gate1018(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate1019(.a(s_67), .b(gate153inter3), .O(gate153inter10));
  nor2  gate1020(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate1021(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate1022(.a(gate153inter12), .b(gate153inter1), .O(G570));
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate855(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate856(.a(gate156inter0), .b(s_44), .O(gate156inter1));
  and2  gate857(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate858(.a(s_44), .O(gate156inter3));
  inv1  gate859(.a(s_45), .O(gate156inter4));
  nand2 gate860(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate861(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate862(.a(G435), .O(gate156inter7));
  inv1  gate863(.a(G525), .O(gate156inter8));
  nand2 gate864(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate865(.a(s_45), .b(gate156inter3), .O(gate156inter10));
  nor2  gate866(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate867(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate868(.a(gate156inter12), .b(gate156inter1), .O(G573));

  xor2  gate1219(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate1220(.a(gate157inter0), .b(s_96), .O(gate157inter1));
  and2  gate1221(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate1222(.a(s_96), .O(gate157inter3));
  inv1  gate1223(.a(s_97), .O(gate157inter4));
  nand2 gate1224(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate1225(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate1226(.a(G438), .O(gate157inter7));
  inv1  gate1227(.a(G528), .O(gate157inter8));
  nand2 gate1228(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate1229(.a(s_97), .b(gate157inter3), .O(gate157inter10));
  nor2  gate1230(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate1231(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate1232(.a(gate157inter12), .b(gate157inter1), .O(G574));

  xor2  gate715(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate716(.a(gate158inter0), .b(s_24), .O(gate158inter1));
  and2  gate717(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate718(.a(s_24), .O(gate158inter3));
  inv1  gate719(.a(s_25), .O(gate158inter4));
  nand2 gate720(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate721(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate722(.a(G441), .O(gate158inter7));
  inv1  gate723(.a(G528), .O(gate158inter8));
  nand2 gate724(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate725(.a(s_25), .b(gate158inter3), .O(gate158inter10));
  nor2  gate726(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate727(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate728(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate1373(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate1374(.a(gate160inter0), .b(s_118), .O(gate160inter1));
  and2  gate1375(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate1376(.a(s_118), .O(gate160inter3));
  inv1  gate1377(.a(s_119), .O(gate160inter4));
  nand2 gate1378(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate1379(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate1380(.a(G447), .O(gate160inter7));
  inv1  gate1381(.a(G531), .O(gate160inter8));
  nand2 gate1382(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate1383(.a(s_119), .b(gate160inter3), .O(gate160inter10));
  nor2  gate1384(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate1385(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate1386(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );

  xor2  gate603(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate604(.a(gate166inter0), .b(s_8), .O(gate166inter1));
  and2  gate605(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate606(.a(s_8), .O(gate166inter3));
  inv1  gate607(.a(s_9), .O(gate166inter4));
  nand2 gate608(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate609(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate610(.a(G465), .O(gate166inter7));
  inv1  gate611(.a(G540), .O(gate166inter8));
  nand2 gate612(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate613(.a(s_9), .b(gate166inter3), .O(gate166inter10));
  nor2  gate614(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate615(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate616(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );

  xor2  gate939(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate940(.a(gate168inter0), .b(s_56), .O(gate168inter1));
  and2  gate941(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate942(.a(s_56), .O(gate168inter3));
  inv1  gate943(.a(s_57), .O(gate168inter4));
  nand2 gate944(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate945(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate946(.a(G471), .O(gate168inter7));
  inv1  gate947(.a(G543), .O(gate168inter8));
  nand2 gate948(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate949(.a(s_57), .b(gate168inter3), .O(gate168inter10));
  nor2  gate950(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate951(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate952(.a(gate168inter12), .b(gate168inter1), .O(G585));
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate1191(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate1192(.a(gate178inter0), .b(s_92), .O(gate178inter1));
  and2  gate1193(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate1194(.a(s_92), .O(gate178inter3));
  inv1  gate1195(.a(s_93), .O(gate178inter4));
  nand2 gate1196(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate1197(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate1198(.a(G501), .O(gate178inter7));
  inv1  gate1199(.a(G558), .O(gate178inter8));
  nand2 gate1200(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate1201(.a(s_93), .b(gate178inter3), .O(gate178inter10));
  nor2  gate1202(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate1203(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate1204(.a(gate178inter12), .b(gate178inter1), .O(G595));
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate701(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate702(.a(gate181inter0), .b(s_22), .O(gate181inter1));
  and2  gate703(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate704(.a(s_22), .O(gate181inter3));
  inv1  gate705(.a(s_23), .O(gate181inter4));
  nand2 gate706(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate707(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate708(.a(G510), .O(gate181inter7));
  inv1  gate709(.a(G564), .O(gate181inter8));
  nand2 gate710(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate711(.a(s_23), .b(gate181inter3), .O(gate181inter10));
  nor2  gate712(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate713(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate714(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate1513(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate1514(.a(gate185inter0), .b(s_138), .O(gate185inter1));
  and2  gate1515(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate1516(.a(s_138), .O(gate185inter3));
  inv1  gate1517(.a(s_139), .O(gate185inter4));
  nand2 gate1518(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate1519(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate1520(.a(G570), .O(gate185inter7));
  inv1  gate1521(.a(G571), .O(gate185inter8));
  nand2 gate1522(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate1523(.a(s_139), .b(gate185inter3), .O(gate185inter10));
  nor2  gate1524(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate1525(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate1526(.a(gate185inter12), .b(gate185inter1), .O(G602));
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );

  xor2  gate1569(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate1570(.a(gate189inter0), .b(s_146), .O(gate189inter1));
  and2  gate1571(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate1572(.a(s_146), .O(gate189inter3));
  inv1  gate1573(.a(s_147), .O(gate189inter4));
  nand2 gate1574(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate1575(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate1576(.a(G578), .O(gate189inter7));
  inv1  gate1577(.a(G579), .O(gate189inter8));
  nand2 gate1578(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate1579(.a(s_147), .b(gate189inter3), .O(gate189inter10));
  nor2  gate1580(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate1581(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate1582(.a(gate189inter12), .b(gate189inter1), .O(G622));
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate1317(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate1318(.a(gate195inter0), .b(s_110), .O(gate195inter1));
  and2  gate1319(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate1320(.a(s_110), .O(gate195inter3));
  inv1  gate1321(.a(s_111), .O(gate195inter4));
  nand2 gate1322(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate1323(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate1324(.a(G590), .O(gate195inter7));
  inv1  gate1325(.a(G591), .O(gate195inter8));
  nand2 gate1326(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate1327(.a(s_111), .b(gate195inter3), .O(gate195inter10));
  nor2  gate1328(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate1329(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate1330(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate1331(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate1332(.a(gate197inter0), .b(s_112), .O(gate197inter1));
  and2  gate1333(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate1334(.a(s_112), .O(gate197inter3));
  inv1  gate1335(.a(s_113), .O(gate197inter4));
  nand2 gate1336(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate1337(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate1338(.a(G594), .O(gate197inter7));
  inv1  gate1339(.a(G595), .O(gate197inter8));
  nand2 gate1340(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate1341(.a(s_113), .b(gate197inter3), .O(gate197inter10));
  nor2  gate1342(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate1343(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate1344(.a(gate197inter12), .b(gate197inter1), .O(G654));

  xor2  gate1443(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate1444(.a(gate198inter0), .b(s_128), .O(gate198inter1));
  and2  gate1445(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate1446(.a(s_128), .O(gate198inter3));
  inv1  gate1447(.a(s_129), .O(gate198inter4));
  nand2 gate1448(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate1449(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate1450(.a(G596), .O(gate198inter7));
  inv1  gate1451(.a(G597), .O(gate198inter8));
  nand2 gate1452(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate1453(.a(s_129), .b(gate198inter3), .O(gate198inter10));
  nor2  gate1454(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate1455(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate1456(.a(gate198inter12), .b(gate198inter1), .O(G657));
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate561(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate562(.a(gate218inter0), .b(s_2), .O(gate218inter1));
  and2  gate563(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate564(.a(s_2), .O(gate218inter3));
  inv1  gate565(.a(s_3), .O(gate218inter4));
  nand2 gate566(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate567(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate568(.a(G627), .O(gate218inter7));
  inv1  gate569(.a(G678), .O(gate218inter8));
  nand2 gate570(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate571(.a(s_3), .b(gate218inter3), .O(gate218inter10));
  nor2  gate572(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate573(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate574(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );

  xor2  gate729(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate730(.a(gate221inter0), .b(s_26), .O(gate221inter1));
  and2  gate731(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate732(.a(s_26), .O(gate221inter3));
  inv1  gate733(.a(s_27), .O(gate221inter4));
  nand2 gate734(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate735(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate736(.a(G622), .O(gate221inter7));
  inv1  gate737(.a(G684), .O(gate221inter8));
  nand2 gate738(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate739(.a(s_27), .b(gate221inter3), .O(gate221inter10));
  nor2  gate740(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate741(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate742(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate589(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate590(.a(gate224inter0), .b(s_6), .O(gate224inter1));
  and2  gate591(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate592(.a(s_6), .O(gate224inter3));
  inv1  gate593(.a(s_7), .O(gate224inter4));
  nand2 gate594(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate595(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate596(.a(G637), .O(gate224inter7));
  inv1  gate597(.a(G687), .O(gate224inter8));
  nand2 gate598(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate599(.a(s_7), .b(gate224inter3), .O(gate224inter10));
  nor2  gate600(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate601(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate602(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );

  xor2  gate1359(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate1360(.a(gate235inter0), .b(s_116), .O(gate235inter1));
  and2  gate1361(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate1362(.a(s_116), .O(gate235inter3));
  inv1  gate1363(.a(s_117), .O(gate235inter4));
  nand2 gate1364(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate1365(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate1366(.a(G248), .O(gate235inter7));
  inv1  gate1367(.a(G724), .O(gate235inter8));
  nand2 gate1368(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate1369(.a(s_117), .b(gate235inter3), .O(gate235inter10));
  nor2  gate1370(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate1371(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate1372(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );

  xor2  gate967(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate968(.a(gate238inter0), .b(s_60), .O(gate238inter1));
  and2  gate969(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate970(.a(s_60), .O(gate238inter3));
  inv1  gate971(.a(s_61), .O(gate238inter4));
  nand2 gate972(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate973(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate974(.a(G257), .O(gate238inter7));
  inv1  gate975(.a(G709), .O(gate238inter8));
  nand2 gate976(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate977(.a(s_61), .b(gate238inter3), .O(gate238inter10));
  nor2  gate978(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate979(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate980(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate869(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate870(.a(gate240inter0), .b(s_46), .O(gate240inter1));
  and2  gate871(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate872(.a(s_46), .O(gate240inter3));
  inv1  gate873(.a(s_47), .O(gate240inter4));
  nand2 gate874(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate875(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate876(.a(G263), .O(gate240inter7));
  inv1  gate877(.a(G715), .O(gate240inter8));
  nand2 gate878(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate879(.a(s_47), .b(gate240inter3), .O(gate240inter10));
  nor2  gate880(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate881(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate882(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );

  xor2  gate1555(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate1556(.a(gate247inter0), .b(s_144), .O(gate247inter1));
  and2  gate1557(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate1558(.a(s_144), .O(gate247inter3));
  inv1  gate1559(.a(s_145), .O(gate247inter4));
  nand2 gate1560(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate1561(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate1562(.a(G251), .O(gate247inter7));
  inv1  gate1563(.a(G739), .O(gate247inter8));
  nand2 gate1564(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate1565(.a(s_145), .b(gate247inter3), .O(gate247inter10));
  nor2  gate1566(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate1567(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate1568(.a(gate247inter12), .b(gate247inter1), .O(G760));
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate1401(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate1402(.a(gate249inter0), .b(s_122), .O(gate249inter1));
  and2  gate1403(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate1404(.a(s_122), .O(gate249inter3));
  inv1  gate1405(.a(s_123), .O(gate249inter4));
  nand2 gate1406(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate1407(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate1408(.a(G254), .O(gate249inter7));
  inv1  gate1409(.a(G742), .O(gate249inter8));
  nand2 gate1410(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate1411(.a(s_123), .b(gate249inter3), .O(gate249inter10));
  nor2  gate1412(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate1413(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate1414(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate799(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate800(.a(gate253inter0), .b(s_36), .O(gate253inter1));
  and2  gate801(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate802(.a(s_36), .O(gate253inter3));
  inv1  gate803(.a(s_37), .O(gate253inter4));
  nand2 gate804(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate805(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate806(.a(G260), .O(gate253inter7));
  inv1  gate807(.a(G748), .O(gate253inter8));
  nand2 gate808(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate809(.a(s_37), .b(gate253inter3), .O(gate253inter10));
  nor2  gate810(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate811(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate812(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate757(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate758(.a(gate257inter0), .b(s_30), .O(gate257inter1));
  and2  gate759(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate760(.a(s_30), .O(gate257inter3));
  inv1  gate761(.a(s_31), .O(gate257inter4));
  nand2 gate762(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate763(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate764(.a(G754), .O(gate257inter7));
  inv1  gate765(.a(G755), .O(gate257inter8));
  nand2 gate766(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate767(.a(s_31), .b(gate257inter3), .O(gate257inter10));
  nor2  gate768(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate769(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate770(.a(gate257inter12), .b(gate257inter1), .O(G770));

  xor2  gate981(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate982(.a(gate258inter0), .b(s_62), .O(gate258inter1));
  and2  gate983(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate984(.a(s_62), .O(gate258inter3));
  inv1  gate985(.a(s_63), .O(gate258inter4));
  nand2 gate986(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate987(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate988(.a(G756), .O(gate258inter7));
  inv1  gate989(.a(G757), .O(gate258inter8));
  nand2 gate990(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate991(.a(s_63), .b(gate258inter3), .O(gate258inter10));
  nor2  gate992(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate993(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate994(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate1597(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate1598(.a(gate261inter0), .b(s_150), .O(gate261inter1));
  and2  gate1599(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate1600(.a(s_150), .O(gate261inter3));
  inv1  gate1601(.a(s_151), .O(gate261inter4));
  nand2 gate1602(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate1603(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate1604(.a(G762), .O(gate261inter7));
  inv1  gate1605(.a(G763), .O(gate261inter8));
  nand2 gate1606(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate1607(.a(s_151), .b(gate261inter3), .O(gate261inter10));
  nor2  gate1608(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate1609(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate1610(.a(gate261inter12), .b(gate261inter1), .O(G782));
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate1499(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate1500(.a(gate268inter0), .b(s_136), .O(gate268inter1));
  and2  gate1501(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate1502(.a(s_136), .O(gate268inter3));
  inv1  gate1503(.a(s_137), .O(gate268inter4));
  nand2 gate1504(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1505(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1506(.a(G651), .O(gate268inter7));
  inv1  gate1507(.a(G779), .O(gate268inter8));
  nand2 gate1508(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1509(.a(s_137), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1510(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1511(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1512(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );

  xor2  gate1429(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate1430(.a(gate273inter0), .b(s_126), .O(gate273inter1));
  and2  gate1431(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate1432(.a(s_126), .O(gate273inter3));
  inv1  gate1433(.a(s_127), .O(gate273inter4));
  nand2 gate1434(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate1435(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate1436(.a(G642), .O(gate273inter7));
  inv1  gate1437(.a(G794), .O(gate273inter8));
  nand2 gate1438(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate1439(.a(s_127), .b(gate273inter3), .O(gate273inter10));
  nor2  gate1440(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate1441(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate1442(.a(gate273inter12), .b(gate273inter1), .O(G818));
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate1205(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate1206(.a(gate278inter0), .b(s_94), .O(gate278inter1));
  and2  gate1207(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate1208(.a(s_94), .O(gate278inter3));
  inv1  gate1209(.a(s_95), .O(gate278inter4));
  nand2 gate1210(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate1211(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate1212(.a(G776), .O(gate278inter7));
  inv1  gate1213(.a(G800), .O(gate278inter8));
  nand2 gate1214(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate1215(.a(s_95), .b(gate278inter3), .O(gate278inter10));
  nor2  gate1216(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate1217(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate1218(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate1037(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate1038(.a(gate285inter0), .b(s_70), .O(gate285inter1));
  and2  gate1039(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate1040(.a(s_70), .O(gate285inter3));
  inv1  gate1041(.a(s_71), .O(gate285inter4));
  nand2 gate1042(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate1043(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate1044(.a(G660), .O(gate285inter7));
  inv1  gate1045(.a(G812), .O(gate285inter8));
  nand2 gate1046(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate1047(.a(s_71), .b(gate285inter3), .O(gate285inter10));
  nor2  gate1048(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate1049(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate1050(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate645(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate646(.a(gate390inter0), .b(s_14), .O(gate390inter1));
  and2  gate647(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate648(.a(s_14), .O(gate390inter3));
  inv1  gate649(.a(s_15), .O(gate390inter4));
  nand2 gate650(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate651(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate652(.a(G4), .O(gate390inter7));
  inv1  gate653(.a(G1045), .O(gate390inter8));
  nand2 gate654(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate655(.a(s_15), .b(gate390inter3), .O(gate390inter10));
  nor2  gate656(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate657(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate658(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate1051(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate1052(.a(gate406inter0), .b(s_72), .O(gate406inter1));
  and2  gate1053(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate1054(.a(s_72), .O(gate406inter3));
  inv1  gate1055(.a(s_73), .O(gate406inter4));
  nand2 gate1056(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate1057(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate1058(.a(G20), .O(gate406inter7));
  inv1  gate1059(.a(G1093), .O(gate406inter8));
  nand2 gate1060(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate1061(.a(s_73), .b(gate406inter3), .O(gate406inter10));
  nor2  gate1062(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate1063(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate1064(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate785(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate786(.a(gate409inter0), .b(s_34), .O(gate409inter1));
  and2  gate787(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate788(.a(s_34), .O(gate409inter3));
  inv1  gate789(.a(s_35), .O(gate409inter4));
  nand2 gate790(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate791(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate792(.a(G23), .O(gate409inter7));
  inv1  gate793(.a(G1102), .O(gate409inter8));
  nand2 gate794(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate795(.a(s_35), .b(gate409inter3), .O(gate409inter10));
  nor2  gate796(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate797(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate798(.a(gate409inter12), .b(gate409inter1), .O(G1198));
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );

  xor2  gate1107(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate1108(.a(gate412inter0), .b(s_80), .O(gate412inter1));
  and2  gate1109(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate1110(.a(s_80), .O(gate412inter3));
  inv1  gate1111(.a(s_81), .O(gate412inter4));
  nand2 gate1112(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate1113(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate1114(.a(G26), .O(gate412inter7));
  inv1  gate1115(.a(G1111), .O(gate412inter8));
  nand2 gate1116(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate1117(.a(s_81), .b(gate412inter3), .O(gate412inter10));
  nor2  gate1118(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate1119(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate1120(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );

  xor2  gate617(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate618(.a(gate414inter0), .b(s_10), .O(gate414inter1));
  and2  gate619(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate620(.a(s_10), .O(gate414inter3));
  inv1  gate621(.a(s_11), .O(gate414inter4));
  nand2 gate622(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate623(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate624(.a(G28), .O(gate414inter7));
  inv1  gate625(.a(G1117), .O(gate414inter8));
  nand2 gate626(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate627(.a(s_11), .b(gate414inter3), .O(gate414inter10));
  nor2  gate628(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate629(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate630(.a(gate414inter12), .b(gate414inter1), .O(G1213));
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );

  xor2  gate827(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate828(.a(gate416inter0), .b(s_40), .O(gate416inter1));
  and2  gate829(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate830(.a(s_40), .O(gate416inter3));
  inv1  gate831(.a(s_41), .O(gate416inter4));
  nand2 gate832(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate833(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate834(.a(G30), .O(gate416inter7));
  inv1  gate835(.a(G1123), .O(gate416inter8));
  nand2 gate836(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate837(.a(s_41), .b(gate416inter3), .O(gate416inter10));
  nor2  gate838(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate839(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate840(.a(gate416inter12), .b(gate416inter1), .O(G1219));

  xor2  gate1261(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate1262(.a(gate417inter0), .b(s_102), .O(gate417inter1));
  and2  gate1263(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate1264(.a(s_102), .O(gate417inter3));
  inv1  gate1265(.a(s_103), .O(gate417inter4));
  nand2 gate1266(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate1267(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate1268(.a(G31), .O(gate417inter7));
  inv1  gate1269(.a(G1126), .O(gate417inter8));
  nand2 gate1270(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate1271(.a(s_103), .b(gate417inter3), .O(gate417inter10));
  nor2  gate1272(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate1273(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate1274(.a(gate417inter12), .b(gate417inter1), .O(G1222));

  xor2  gate1163(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate1164(.a(gate418inter0), .b(s_88), .O(gate418inter1));
  and2  gate1165(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate1166(.a(s_88), .O(gate418inter3));
  inv1  gate1167(.a(s_89), .O(gate418inter4));
  nand2 gate1168(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate1169(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate1170(.a(G32), .O(gate418inter7));
  inv1  gate1171(.a(G1129), .O(gate418inter8));
  nand2 gate1172(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate1173(.a(s_89), .b(gate418inter3), .O(gate418inter10));
  nor2  gate1174(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate1175(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate1176(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );

  xor2  gate1303(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate1304(.a(gate423inter0), .b(s_108), .O(gate423inter1));
  and2  gate1305(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate1306(.a(s_108), .O(gate423inter3));
  inv1  gate1307(.a(s_109), .O(gate423inter4));
  nand2 gate1308(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate1309(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate1310(.a(G3), .O(gate423inter7));
  inv1  gate1311(.a(G1138), .O(gate423inter8));
  nand2 gate1312(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate1313(.a(s_109), .b(gate423inter3), .O(gate423inter10));
  nor2  gate1314(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate1315(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate1316(.a(gate423inter12), .b(gate423inter1), .O(G1232));
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate1583(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate1584(.a(gate425inter0), .b(s_148), .O(gate425inter1));
  and2  gate1585(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate1586(.a(s_148), .O(gate425inter3));
  inv1  gate1587(.a(s_149), .O(gate425inter4));
  nand2 gate1588(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1589(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1590(.a(G4), .O(gate425inter7));
  inv1  gate1591(.a(G1141), .O(gate425inter8));
  nand2 gate1592(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1593(.a(s_149), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1594(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1595(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1596(.a(gate425inter12), .b(gate425inter1), .O(G1234));
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate1177(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate1178(.a(gate442inter0), .b(s_90), .O(gate442inter1));
  and2  gate1179(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate1180(.a(s_90), .O(gate442inter3));
  inv1  gate1181(.a(s_91), .O(gate442inter4));
  nand2 gate1182(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate1183(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate1184(.a(G1069), .O(gate442inter7));
  inv1  gate1185(.a(G1165), .O(gate442inter8));
  nand2 gate1186(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate1187(.a(s_91), .b(gate442inter3), .O(gate442inter10));
  nor2  gate1188(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate1189(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate1190(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );

  xor2  gate1527(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate1528(.a(gate449inter0), .b(s_140), .O(gate449inter1));
  and2  gate1529(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate1530(.a(s_140), .O(gate449inter3));
  inv1  gate1531(.a(s_141), .O(gate449inter4));
  nand2 gate1532(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate1533(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate1534(.a(G16), .O(gate449inter7));
  inv1  gate1535(.a(G1177), .O(gate449inter8));
  nand2 gate1536(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate1537(.a(s_141), .b(gate449inter3), .O(gate449inter10));
  nor2  gate1538(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate1539(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate1540(.a(gate449inter12), .b(gate449inter1), .O(G1258));

  xor2  gate911(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate912(.a(gate450inter0), .b(s_52), .O(gate450inter1));
  and2  gate913(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate914(.a(s_52), .O(gate450inter3));
  inv1  gate915(.a(s_53), .O(gate450inter4));
  nand2 gate916(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate917(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate918(.a(G1081), .O(gate450inter7));
  inv1  gate919(.a(G1177), .O(gate450inter8));
  nand2 gate920(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate921(.a(s_53), .b(gate450inter3), .O(gate450inter10));
  nor2  gate922(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate923(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate924(.a(gate450inter12), .b(gate450inter1), .O(G1259));
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate1121(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate1122(.a(gate453inter0), .b(s_82), .O(gate453inter1));
  and2  gate1123(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate1124(.a(s_82), .O(gate453inter3));
  inv1  gate1125(.a(s_83), .O(gate453inter4));
  nand2 gate1126(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate1127(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate1128(.a(G18), .O(gate453inter7));
  inv1  gate1129(.a(G1183), .O(gate453inter8));
  nand2 gate1130(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate1131(.a(s_83), .b(gate453inter3), .O(gate453inter10));
  nor2  gate1132(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate1133(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate1134(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate1387(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate1388(.a(gate463inter0), .b(s_120), .O(gate463inter1));
  and2  gate1389(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate1390(.a(s_120), .O(gate463inter3));
  inv1  gate1391(.a(s_121), .O(gate463inter4));
  nand2 gate1392(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate1393(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate1394(.a(G23), .O(gate463inter7));
  inv1  gate1395(.a(G1198), .O(gate463inter8));
  nand2 gate1396(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate1397(.a(s_121), .b(gate463inter3), .O(gate463inter10));
  nor2  gate1398(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate1399(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate1400(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate659(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate660(.a(gate477inter0), .b(s_16), .O(gate477inter1));
  and2  gate661(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate662(.a(s_16), .O(gate477inter3));
  inv1  gate663(.a(s_17), .O(gate477inter4));
  nand2 gate664(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate665(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate666(.a(G30), .O(gate477inter7));
  inv1  gate667(.a(G1219), .O(gate477inter8));
  nand2 gate668(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate669(.a(s_17), .b(gate477inter3), .O(gate477inter10));
  nor2  gate670(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate671(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate672(.a(gate477inter12), .b(gate477inter1), .O(G1286));

  xor2  gate1247(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate1248(.a(gate478inter0), .b(s_100), .O(gate478inter1));
  and2  gate1249(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate1250(.a(s_100), .O(gate478inter3));
  inv1  gate1251(.a(s_101), .O(gate478inter4));
  nand2 gate1252(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate1253(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate1254(.a(G1123), .O(gate478inter7));
  inv1  gate1255(.a(G1219), .O(gate478inter8));
  nand2 gate1256(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate1257(.a(s_101), .b(gate478inter3), .O(gate478inter10));
  nor2  gate1258(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate1259(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate1260(.a(gate478inter12), .b(gate478inter1), .O(G1287));
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate1093(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate1094(.a(gate492inter0), .b(s_78), .O(gate492inter1));
  and2  gate1095(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate1096(.a(s_78), .O(gate492inter3));
  inv1  gate1097(.a(s_79), .O(gate492inter4));
  nand2 gate1098(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate1099(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate1100(.a(G1246), .O(gate492inter7));
  inv1  gate1101(.a(G1247), .O(gate492inter8));
  nand2 gate1102(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate1103(.a(s_79), .b(gate492inter3), .O(gate492inter10));
  nor2  gate1104(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate1105(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate1106(.a(gate492inter12), .b(gate492inter1), .O(G1301));
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate1079(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1080(.a(gate494inter0), .b(s_76), .O(gate494inter1));
  and2  gate1081(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1082(.a(s_76), .O(gate494inter3));
  inv1  gate1083(.a(s_77), .O(gate494inter4));
  nand2 gate1084(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1085(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1086(.a(G1250), .O(gate494inter7));
  inv1  gate1087(.a(G1251), .O(gate494inter8));
  nand2 gate1088(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1089(.a(s_77), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1090(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1091(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1092(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate1135(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate1136(.a(gate497inter0), .b(s_84), .O(gate497inter1));
  and2  gate1137(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate1138(.a(s_84), .O(gate497inter3));
  inv1  gate1139(.a(s_85), .O(gate497inter4));
  nand2 gate1140(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate1141(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate1142(.a(G1256), .O(gate497inter7));
  inv1  gate1143(.a(G1257), .O(gate497inter8));
  nand2 gate1144(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate1145(.a(s_85), .b(gate497inter3), .O(gate497inter10));
  nor2  gate1146(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate1147(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate1148(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate1541(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate1542(.a(gate502inter0), .b(s_142), .O(gate502inter1));
  and2  gate1543(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate1544(.a(s_142), .O(gate502inter3));
  inv1  gate1545(.a(s_143), .O(gate502inter4));
  nand2 gate1546(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate1547(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate1548(.a(G1266), .O(gate502inter7));
  inv1  gate1549(.a(G1267), .O(gate502inter8));
  nand2 gate1550(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate1551(.a(s_143), .b(gate502inter3), .O(gate502inter10));
  nor2  gate1552(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate1553(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate1554(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );

  xor2  gate673(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate674(.a(gate505inter0), .b(s_18), .O(gate505inter1));
  and2  gate675(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate676(.a(s_18), .O(gate505inter3));
  inv1  gate677(.a(s_19), .O(gate505inter4));
  nand2 gate678(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate679(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate680(.a(G1272), .O(gate505inter7));
  inv1  gate681(.a(G1273), .O(gate505inter8));
  nand2 gate682(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate683(.a(s_19), .b(gate505inter3), .O(gate505inter10));
  nor2  gate684(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate685(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate686(.a(gate505inter12), .b(gate505inter1), .O(G1314));
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule