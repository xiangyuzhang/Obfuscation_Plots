module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate1177(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate1178(.a(gate11inter0), .b(s_90), .O(gate11inter1));
  and2  gate1179(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate1180(.a(s_90), .O(gate11inter3));
  inv1  gate1181(.a(s_91), .O(gate11inter4));
  nand2 gate1182(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate1183(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate1184(.a(G5), .O(gate11inter7));
  inv1  gate1185(.a(G6), .O(gate11inter8));
  nand2 gate1186(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate1187(.a(s_91), .b(gate11inter3), .O(gate11inter10));
  nor2  gate1188(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate1189(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate1190(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate1499(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate1500(.a(gate13inter0), .b(s_136), .O(gate13inter1));
  and2  gate1501(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate1502(.a(s_136), .O(gate13inter3));
  inv1  gate1503(.a(s_137), .O(gate13inter4));
  nand2 gate1504(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate1505(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate1506(.a(G9), .O(gate13inter7));
  inv1  gate1507(.a(G10), .O(gate13inter8));
  nand2 gate1508(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate1509(.a(s_137), .b(gate13inter3), .O(gate13inter10));
  nor2  gate1510(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate1511(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate1512(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate1863(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate1864(.a(gate17inter0), .b(s_188), .O(gate17inter1));
  and2  gate1865(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate1866(.a(s_188), .O(gate17inter3));
  inv1  gate1867(.a(s_189), .O(gate17inter4));
  nand2 gate1868(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate1869(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate1870(.a(G17), .O(gate17inter7));
  inv1  gate1871(.a(G18), .O(gate17inter8));
  nand2 gate1872(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate1873(.a(s_189), .b(gate17inter3), .O(gate17inter10));
  nor2  gate1874(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate1875(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate1876(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate561(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate562(.a(gate23inter0), .b(s_2), .O(gate23inter1));
  and2  gate563(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate564(.a(s_2), .O(gate23inter3));
  inv1  gate565(.a(s_3), .O(gate23inter4));
  nand2 gate566(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate567(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate568(.a(G29), .O(gate23inter7));
  inv1  gate569(.a(G30), .O(gate23inter8));
  nand2 gate570(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate571(.a(s_3), .b(gate23inter3), .O(gate23inter10));
  nor2  gate572(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate573(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate574(.a(gate23inter12), .b(gate23inter1), .O(G308));

  xor2  gate1247(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate1248(.a(gate24inter0), .b(s_100), .O(gate24inter1));
  and2  gate1249(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate1250(.a(s_100), .O(gate24inter3));
  inv1  gate1251(.a(s_101), .O(gate24inter4));
  nand2 gate1252(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate1253(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate1254(.a(G31), .O(gate24inter7));
  inv1  gate1255(.a(G32), .O(gate24inter8));
  nand2 gate1256(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate1257(.a(s_101), .b(gate24inter3), .O(gate24inter10));
  nor2  gate1258(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate1259(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate1260(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate1121(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1122(.a(gate36inter0), .b(s_82), .O(gate36inter1));
  and2  gate1123(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1124(.a(s_82), .O(gate36inter3));
  inv1  gate1125(.a(s_83), .O(gate36inter4));
  nand2 gate1126(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1127(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1128(.a(G26), .O(gate36inter7));
  inv1  gate1129(.a(G30), .O(gate36inter8));
  nand2 gate1130(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1131(.a(s_83), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1132(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1133(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1134(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate687(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate688(.a(gate46inter0), .b(s_20), .O(gate46inter1));
  and2  gate689(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate690(.a(s_20), .O(gate46inter3));
  inv1  gate691(.a(s_21), .O(gate46inter4));
  nand2 gate692(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate693(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate694(.a(G6), .O(gate46inter7));
  inv1  gate695(.a(G272), .O(gate46inter8));
  nand2 gate696(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate697(.a(s_21), .b(gate46inter3), .O(gate46inter10));
  nor2  gate698(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate699(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate700(.a(gate46inter12), .b(gate46inter1), .O(G367));

  xor2  gate1779(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate1780(.a(gate47inter0), .b(s_176), .O(gate47inter1));
  and2  gate1781(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate1782(.a(s_176), .O(gate47inter3));
  inv1  gate1783(.a(s_177), .O(gate47inter4));
  nand2 gate1784(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate1785(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate1786(.a(G7), .O(gate47inter7));
  inv1  gate1787(.a(G275), .O(gate47inter8));
  nand2 gate1788(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate1789(.a(s_177), .b(gate47inter3), .O(gate47inter10));
  nor2  gate1790(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate1791(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate1792(.a(gate47inter12), .b(gate47inter1), .O(G368));
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate841(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate842(.a(gate57inter0), .b(s_42), .O(gate57inter1));
  and2  gate843(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate844(.a(s_42), .O(gate57inter3));
  inv1  gate845(.a(s_43), .O(gate57inter4));
  nand2 gate846(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate847(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate848(.a(G17), .O(gate57inter7));
  inv1  gate849(.a(G290), .O(gate57inter8));
  nand2 gate850(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate851(.a(s_43), .b(gate57inter3), .O(gate57inter10));
  nor2  gate852(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate853(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate854(.a(gate57inter12), .b(gate57inter1), .O(G378));
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate1513(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate1514(.a(gate60inter0), .b(s_138), .O(gate60inter1));
  and2  gate1515(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate1516(.a(s_138), .O(gate60inter3));
  inv1  gate1517(.a(s_139), .O(gate60inter4));
  nand2 gate1518(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate1519(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate1520(.a(G20), .O(gate60inter7));
  inv1  gate1521(.a(G293), .O(gate60inter8));
  nand2 gate1522(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate1523(.a(s_139), .b(gate60inter3), .O(gate60inter10));
  nor2  gate1524(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate1525(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate1526(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate1597(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate1598(.a(gate63inter0), .b(s_150), .O(gate63inter1));
  and2  gate1599(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate1600(.a(s_150), .O(gate63inter3));
  inv1  gate1601(.a(s_151), .O(gate63inter4));
  nand2 gate1602(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate1603(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate1604(.a(G23), .O(gate63inter7));
  inv1  gate1605(.a(G299), .O(gate63inter8));
  nand2 gate1606(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate1607(.a(s_151), .b(gate63inter3), .O(gate63inter10));
  nor2  gate1608(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate1609(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate1610(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate1751(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate1752(.a(gate66inter0), .b(s_172), .O(gate66inter1));
  and2  gate1753(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate1754(.a(s_172), .O(gate66inter3));
  inv1  gate1755(.a(s_173), .O(gate66inter4));
  nand2 gate1756(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate1757(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate1758(.a(G26), .O(gate66inter7));
  inv1  gate1759(.a(G302), .O(gate66inter8));
  nand2 gate1760(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate1761(.a(s_173), .b(gate66inter3), .O(gate66inter10));
  nor2  gate1762(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate1763(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate1764(.a(gate66inter12), .b(gate66inter1), .O(G387));

  xor2  gate939(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate940(.a(gate67inter0), .b(s_56), .O(gate67inter1));
  and2  gate941(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate942(.a(s_56), .O(gate67inter3));
  inv1  gate943(.a(s_57), .O(gate67inter4));
  nand2 gate944(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate945(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate946(.a(G27), .O(gate67inter7));
  inv1  gate947(.a(G305), .O(gate67inter8));
  nand2 gate948(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate949(.a(s_57), .b(gate67inter3), .O(gate67inter10));
  nor2  gate950(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate951(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate952(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );

  xor2  gate1303(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate1304(.a(gate72inter0), .b(s_108), .O(gate72inter1));
  and2  gate1305(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate1306(.a(s_108), .O(gate72inter3));
  inv1  gate1307(.a(s_109), .O(gate72inter4));
  nand2 gate1308(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate1309(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate1310(.a(G32), .O(gate72inter7));
  inv1  gate1311(.a(G311), .O(gate72inter8));
  nand2 gate1312(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate1313(.a(s_109), .b(gate72inter3), .O(gate72inter10));
  nor2  gate1314(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate1315(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate1316(.a(gate72inter12), .b(gate72inter1), .O(G393));

  xor2  gate1681(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate1682(.a(gate73inter0), .b(s_162), .O(gate73inter1));
  and2  gate1683(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate1684(.a(s_162), .O(gate73inter3));
  inv1  gate1685(.a(s_163), .O(gate73inter4));
  nand2 gate1686(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate1687(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate1688(.a(G1), .O(gate73inter7));
  inv1  gate1689(.a(G314), .O(gate73inter8));
  nand2 gate1690(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate1691(.a(s_163), .b(gate73inter3), .O(gate73inter10));
  nor2  gate1692(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate1693(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate1694(.a(gate73inter12), .b(gate73inter1), .O(G394));
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate1807(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate1808(.a(gate75inter0), .b(s_180), .O(gate75inter1));
  and2  gate1809(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate1810(.a(s_180), .O(gate75inter3));
  inv1  gate1811(.a(s_181), .O(gate75inter4));
  nand2 gate1812(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate1813(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate1814(.a(G9), .O(gate75inter7));
  inv1  gate1815(.a(G317), .O(gate75inter8));
  nand2 gate1816(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate1817(.a(s_181), .b(gate75inter3), .O(gate75inter10));
  nor2  gate1818(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate1819(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate1820(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate1765(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate1766(.a(gate96inter0), .b(s_174), .O(gate96inter1));
  and2  gate1767(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate1768(.a(s_174), .O(gate96inter3));
  inv1  gate1769(.a(s_175), .O(gate96inter4));
  nand2 gate1770(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate1771(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate1772(.a(G30), .O(gate96inter7));
  inv1  gate1773(.a(G347), .O(gate96inter8));
  nand2 gate1774(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate1775(.a(s_175), .b(gate96inter3), .O(gate96inter10));
  nor2  gate1776(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate1777(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate1778(.a(gate96inter12), .b(gate96inter1), .O(G417));
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate1387(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate1388(.a(gate100inter0), .b(s_120), .O(gate100inter1));
  and2  gate1389(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate1390(.a(s_120), .O(gate100inter3));
  inv1  gate1391(.a(s_121), .O(gate100inter4));
  nand2 gate1392(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate1393(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate1394(.a(G31), .O(gate100inter7));
  inv1  gate1395(.a(G353), .O(gate100inter8));
  nand2 gate1396(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate1397(.a(s_121), .b(gate100inter3), .O(gate100inter10));
  nor2  gate1398(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate1399(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate1400(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );

  xor2  gate659(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate660(.a(gate103inter0), .b(s_16), .O(gate103inter1));
  and2  gate661(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate662(.a(s_16), .O(gate103inter3));
  inv1  gate663(.a(s_17), .O(gate103inter4));
  nand2 gate664(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate665(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate666(.a(G28), .O(gate103inter7));
  inv1  gate667(.a(G359), .O(gate103inter8));
  nand2 gate668(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate669(.a(s_17), .b(gate103inter3), .O(gate103inter10));
  nor2  gate670(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate671(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate672(.a(gate103inter12), .b(gate103inter1), .O(G424));

  xor2  gate1149(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate1150(.a(gate104inter0), .b(s_86), .O(gate104inter1));
  and2  gate1151(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate1152(.a(s_86), .O(gate104inter3));
  inv1  gate1153(.a(s_87), .O(gate104inter4));
  nand2 gate1154(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate1155(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate1156(.a(G32), .O(gate104inter7));
  inv1  gate1157(.a(G359), .O(gate104inter8));
  nand2 gate1158(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate1159(.a(s_87), .b(gate104inter3), .O(gate104inter10));
  nor2  gate1160(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate1161(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate1162(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );

  xor2  gate953(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate954(.a(gate111inter0), .b(s_58), .O(gate111inter1));
  and2  gate955(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate956(.a(s_58), .O(gate111inter3));
  inv1  gate957(.a(s_59), .O(gate111inter4));
  nand2 gate958(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate959(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate960(.a(G374), .O(gate111inter7));
  inv1  gate961(.a(G375), .O(gate111inter8));
  nand2 gate962(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate963(.a(s_59), .b(gate111inter3), .O(gate111inter10));
  nor2  gate964(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate965(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate966(.a(gate111inter12), .b(gate111inter1), .O(G444));
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate855(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate856(.a(gate117inter0), .b(s_44), .O(gate117inter1));
  and2  gate857(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate858(.a(s_44), .O(gate117inter3));
  inv1  gate859(.a(s_45), .O(gate117inter4));
  nand2 gate860(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate861(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate862(.a(G386), .O(gate117inter7));
  inv1  gate863(.a(G387), .O(gate117inter8));
  nand2 gate864(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate865(.a(s_45), .b(gate117inter3), .O(gate117inter10));
  nor2  gate866(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate867(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate868(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate1037(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate1038(.a(gate119inter0), .b(s_70), .O(gate119inter1));
  and2  gate1039(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate1040(.a(s_70), .O(gate119inter3));
  inv1  gate1041(.a(s_71), .O(gate119inter4));
  nand2 gate1042(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate1043(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate1044(.a(G390), .O(gate119inter7));
  inv1  gate1045(.a(G391), .O(gate119inter8));
  nand2 gate1046(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate1047(.a(s_71), .b(gate119inter3), .O(gate119inter10));
  nor2  gate1048(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate1049(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate1050(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate1051(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate1052(.a(gate126inter0), .b(s_72), .O(gate126inter1));
  and2  gate1053(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate1054(.a(s_72), .O(gate126inter3));
  inv1  gate1055(.a(s_73), .O(gate126inter4));
  nand2 gate1056(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate1057(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate1058(.a(G404), .O(gate126inter7));
  inv1  gate1059(.a(G405), .O(gate126inter8));
  nand2 gate1060(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate1061(.a(s_73), .b(gate126inter3), .O(gate126inter10));
  nor2  gate1062(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate1063(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate1064(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate827(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate828(.a(gate130inter0), .b(s_40), .O(gate130inter1));
  and2  gate829(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate830(.a(s_40), .O(gate130inter3));
  inv1  gate831(.a(s_41), .O(gate130inter4));
  nand2 gate832(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate833(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate834(.a(G412), .O(gate130inter7));
  inv1  gate835(.a(G413), .O(gate130inter8));
  nand2 gate836(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate837(.a(s_41), .b(gate130inter3), .O(gate130inter10));
  nor2  gate838(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate839(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate840(.a(gate130inter12), .b(gate130inter1), .O(G501));
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate883(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate884(.a(gate132inter0), .b(s_48), .O(gate132inter1));
  and2  gate885(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate886(.a(s_48), .O(gate132inter3));
  inv1  gate887(.a(s_49), .O(gate132inter4));
  nand2 gate888(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate889(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate890(.a(G416), .O(gate132inter7));
  inv1  gate891(.a(G417), .O(gate132inter8));
  nand2 gate892(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate893(.a(s_49), .b(gate132inter3), .O(gate132inter10));
  nor2  gate894(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate895(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate896(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate1065(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate1066(.a(gate138inter0), .b(s_74), .O(gate138inter1));
  and2  gate1067(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate1068(.a(s_74), .O(gate138inter3));
  inv1  gate1069(.a(s_75), .O(gate138inter4));
  nand2 gate1070(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate1071(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate1072(.a(G432), .O(gate138inter7));
  inv1  gate1073(.a(G435), .O(gate138inter8));
  nand2 gate1074(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate1075(.a(s_75), .b(gate138inter3), .O(gate138inter10));
  nor2  gate1076(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate1077(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate1078(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate1667(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate1668(.a(gate150inter0), .b(s_160), .O(gate150inter1));
  and2  gate1669(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate1670(.a(s_160), .O(gate150inter3));
  inv1  gate1671(.a(s_161), .O(gate150inter4));
  nand2 gate1672(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate1673(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate1674(.a(G504), .O(gate150inter7));
  inv1  gate1675(.a(G507), .O(gate150inter8));
  nand2 gate1676(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate1677(.a(s_161), .b(gate150inter3), .O(gate150inter10));
  nor2  gate1678(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate1679(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate1680(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate1527(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate1528(.a(gate159inter0), .b(s_140), .O(gate159inter1));
  and2  gate1529(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate1530(.a(s_140), .O(gate159inter3));
  inv1  gate1531(.a(s_141), .O(gate159inter4));
  nand2 gate1532(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate1533(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate1534(.a(G444), .O(gate159inter7));
  inv1  gate1535(.a(G531), .O(gate159inter8));
  nand2 gate1536(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate1537(.a(s_141), .b(gate159inter3), .O(gate159inter10));
  nor2  gate1538(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate1539(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate1540(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate1695(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate1696(.a(gate165inter0), .b(s_164), .O(gate165inter1));
  and2  gate1697(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate1698(.a(s_164), .O(gate165inter3));
  inv1  gate1699(.a(s_165), .O(gate165inter4));
  nand2 gate1700(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate1701(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate1702(.a(G462), .O(gate165inter7));
  inv1  gate1703(.a(G540), .O(gate165inter8));
  nand2 gate1704(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate1705(.a(s_165), .b(gate165inter3), .O(gate165inter10));
  nor2  gate1706(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate1707(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate1708(.a(gate165inter12), .b(gate165inter1), .O(G582));

  xor2  gate729(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate730(.a(gate166inter0), .b(s_26), .O(gate166inter1));
  and2  gate731(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate732(.a(s_26), .O(gate166inter3));
  inv1  gate733(.a(s_27), .O(gate166inter4));
  nand2 gate734(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate735(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate736(.a(G465), .O(gate166inter7));
  inv1  gate737(.a(G540), .O(gate166inter8));
  nand2 gate738(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate739(.a(s_27), .b(gate166inter3), .O(gate166inter10));
  nor2  gate740(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate741(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate742(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate1821(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate1822(.a(gate172inter0), .b(s_182), .O(gate172inter1));
  and2  gate1823(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate1824(.a(s_182), .O(gate172inter3));
  inv1  gate1825(.a(s_183), .O(gate172inter4));
  nand2 gate1826(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate1827(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate1828(.a(G483), .O(gate172inter7));
  inv1  gate1829(.a(G549), .O(gate172inter8));
  nand2 gate1830(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate1831(.a(s_183), .b(gate172inter3), .O(gate172inter10));
  nor2  gate1832(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate1833(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate1834(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate1485(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate1486(.a(gate185inter0), .b(s_134), .O(gate185inter1));
  and2  gate1487(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate1488(.a(s_134), .O(gate185inter3));
  inv1  gate1489(.a(s_135), .O(gate185inter4));
  nand2 gate1490(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate1491(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate1492(.a(G570), .O(gate185inter7));
  inv1  gate1493(.a(G571), .O(gate185inter8));
  nand2 gate1494(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate1495(.a(s_135), .b(gate185inter3), .O(gate185inter10));
  nor2  gate1496(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate1497(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate1498(.a(gate185inter12), .b(gate185inter1), .O(G602));
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate911(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate912(.a(gate187inter0), .b(s_52), .O(gate187inter1));
  and2  gate913(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate914(.a(s_52), .O(gate187inter3));
  inv1  gate915(.a(s_53), .O(gate187inter4));
  nand2 gate916(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate917(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate918(.a(G574), .O(gate187inter7));
  inv1  gate919(.a(G575), .O(gate187inter8));
  nand2 gate920(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate921(.a(s_53), .b(gate187inter3), .O(gate187inter10));
  nor2  gate922(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate923(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate924(.a(gate187inter12), .b(gate187inter1), .O(G612));
nand2 gate188( .a(G576), .b(G577), .O(G617) );

  xor2  gate631(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate632(.a(gate189inter0), .b(s_12), .O(gate189inter1));
  and2  gate633(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate634(.a(s_12), .O(gate189inter3));
  inv1  gate635(.a(s_13), .O(gate189inter4));
  nand2 gate636(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate637(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate638(.a(G578), .O(gate189inter7));
  inv1  gate639(.a(G579), .O(gate189inter8));
  nand2 gate640(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate641(.a(s_13), .b(gate189inter3), .O(gate189inter10));
  nor2  gate642(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate643(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate644(.a(gate189inter12), .b(gate189inter1), .O(G622));

  xor2  gate1625(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate1626(.a(gate190inter0), .b(s_154), .O(gate190inter1));
  and2  gate1627(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate1628(.a(s_154), .O(gate190inter3));
  inv1  gate1629(.a(s_155), .O(gate190inter4));
  nand2 gate1630(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate1631(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate1632(.a(G580), .O(gate190inter7));
  inv1  gate1633(.a(G581), .O(gate190inter8));
  nand2 gate1634(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate1635(.a(s_155), .b(gate190inter3), .O(gate190inter10));
  nor2  gate1636(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate1637(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate1638(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate1569(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate1570(.a(gate193inter0), .b(s_146), .O(gate193inter1));
  and2  gate1571(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate1572(.a(s_146), .O(gate193inter3));
  inv1  gate1573(.a(s_147), .O(gate193inter4));
  nand2 gate1574(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate1575(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate1576(.a(G586), .O(gate193inter7));
  inv1  gate1577(.a(G587), .O(gate193inter8));
  nand2 gate1578(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate1579(.a(s_147), .b(gate193inter3), .O(gate193inter10));
  nor2  gate1580(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate1581(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate1582(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate1219(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate1220(.a(gate196inter0), .b(s_96), .O(gate196inter1));
  and2  gate1221(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate1222(.a(s_96), .O(gate196inter3));
  inv1  gate1223(.a(s_97), .O(gate196inter4));
  nand2 gate1224(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate1225(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate1226(.a(G592), .O(gate196inter7));
  inv1  gate1227(.a(G593), .O(gate196inter8));
  nand2 gate1228(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate1229(.a(s_97), .b(gate196inter3), .O(gate196inter10));
  nor2  gate1230(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate1231(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate1232(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate1317(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate1318(.a(gate205inter0), .b(s_110), .O(gate205inter1));
  and2  gate1319(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate1320(.a(s_110), .O(gate205inter3));
  inv1  gate1321(.a(s_111), .O(gate205inter4));
  nand2 gate1322(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate1323(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate1324(.a(G622), .O(gate205inter7));
  inv1  gate1325(.a(G627), .O(gate205inter8));
  nand2 gate1326(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate1327(.a(s_111), .b(gate205inter3), .O(gate205inter10));
  nor2  gate1328(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate1329(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate1330(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );

  xor2  gate1093(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate1094(.a(gate208inter0), .b(s_78), .O(gate208inter1));
  and2  gate1095(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate1096(.a(s_78), .O(gate208inter3));
  inv1  gate1097(.a(s_79), .O(gate208inter4));
  nand2 gate1098(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate1099(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate1100(.a(G627), .O(gate208inter7));
  inv1  gate1101(.a(G637), .O(gate208inter8));
  nand2 gate1102(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate1103(.a(s_79), .b(gate208inter3), .O(gate208inter10));
  nor2  gate1104(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate1105(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate1106(.a(gate208inter12), .b(gate208inter1), .O(G687));
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate1373(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate1374(.a(gate214inter0), .b(s_118), .O(gate214inter1));
  and2  gate1375(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate1376(.a(s_118), .O(gate214inter3));
  inv1  gate1377(.a(s_119), .O(gate214inter4));
  nand2 gate1378(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate1379(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate1380(.a(G612), .O(gate214inter7));
  inv1  gate1381(.a(G672), .O(gate214inter8));
  nand2 gate1382(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate1383(.a(s_119), .b(gate214inter3), .O(gate214inter10));
  nor2  gate1384(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate1385(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate1386(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );

  xor2  gate1135(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate1136(.a(gate222inter0), .b(s_84), .O(gate222inter1));
  and2  gate1137(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate1138(.a(s_84), .O(gate222inter3));
  inv1  gate1139(.a(s_85), .O(gate222inter4));
  nand2 gate1140(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate1141(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate1142(.a(G632), .O(gate222inter7));
  inv1  gate1143(.a(G684), .O(gate222inter8));
  nand2 gate1144(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate1145(.a(s_85), .b(gate222inter3), .O(gate222inter10));
  nor2  gate1146(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate1147(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate1148(.a(gate222inter12), .b(gate222inter1), .O(G703));

  xor2  gate1583(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate1584(.a(gate223inter0), .b(s_148), .O(gate223inter1));
  and2  gate1585(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate1586(.a(s_148), .O(gate223inter3));
  inv1  gate1587(.a(s_149), .O(gate223inter4));
  nand2 gate1588(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate1589(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate1590(.a(G627), .O(gate223inter7));
  inv1  gate1591(.a(G687), .O(gate223inter8));
  nand2 gate1592(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate1593(.a(s_149), .b(gate223inter3), .O(gate223inter10));
  nor2  gate1594(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate1595(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate1596(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate771(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate772(.a(gate226inter0), .b(s_32), .O(gate226inter1));
  and2  gate773(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate774(.a(s_32), .O(gate226inter3));
  inv1  gate775(.a(s_33), .O(gate226inter4));
  nand2 gate776(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate777(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate778(.a(G692), .O(gate226inter7));
  inv1  gate779(.a(G693), .O(gate226inter8));
  nand2 gate780(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate781(.a(s_33), .b(gate226inter3), .O(gate226inter10));
  nor2  gate782(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate783(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate784(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate1205(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate1206(.a(gate228inter0), .b(s_94), .O(gate228inter1));
  and2  gate1207(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate1208(.a(s_94), .O(gate228inter3));
  inv1  gate1209(.a(s_95), .O(gate228inter4));
  nand2 gate1210(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate1211(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate1212(.a(G696), .O(gate228inter7));
  inv1  gate1213(.a(G697), .O(gate228inter8));
  nand2 gate1214(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate1215(.a(s_95), .b(gate228inter3), .O(gate228inter10));
  nor2  gate1216(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate1217(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate1218(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate1331(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate1332(.a(gate231inter0), .b(s_112), .O(gate231inter1));
  and2  gate1333(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate1334(.a(s_112), .O(gate231inter3));
  inv1  gate1335(.a(s_113), .O(gate231inter4));
  nand2 gate1336(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate1337(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate1338(.a(G702), .O(gate231inter7));
  inv1  gate1339(.a(G703), .O(gate231inter8));
  nand2 gate1340(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate1341(.a(s_113), .b(gate231inter3), .O(gate231inter10));
  nor2  gate1342(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate1343(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate1344(.a(gate231inter12), .b(gate231inter1), .O(G724));

  xor2  gate1793(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate1794(.a(gate232inter0), .b(s_178), .O(gate232inter1));
  and2  gate1795(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate1796(.a(s_178), .O(gate232inter3));
  inv1  gate1797(.a(s_179), .O(gate232inter4));
  nand2 gate1798(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate1799(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate1800(.a(G704), .O(gate232inter7));
  inv1  gate1801(.a(G705), .O(gate232inter8));
  nand2 gate1802(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate1803(.a(s_179), .b(gate232inter3), .O(gate232inter10));
  nor2  gate1804(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate1805(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate1806(.a(gate232inter12), .b(gate232inter1), .O(G727));
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );

  xor2  gate1401(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate1402(.a(gate235inter0), .b(s_122), .O(gate235inter1));
  and2  gate1403(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate1404(.a(s_122), .O(gate235inter3));
  inv1  gate1405(.a(s_123), .O(gate235inter4));
  nand2 gate1406(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate1407(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate1408(.a(G248), .O(gate235inter7));
  inv1  gate1409(.a(G724), .O(gate235inter8));
  nand2 gate1410(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate1411(.a(s_123), .b(gate235inter3), .O(gate235inter10));
  nor2  gate1412(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate1413(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate1414(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate995(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate996(.a(gate237inter0), .b(s_64), .O(gate237inter1));
  and2  gate997(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate998(.a(s_64), .O(gate237inter3));
  inv1  gate999(.a(s_65), .O(gate237inter4));
  nand2 gate1000(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1001(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1002(.a(G254), .O(gate237inter7));
  inv1  gate1003(.a(G706), .O(gate237inter8));
  nand2 gate1004(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1005(.a(s_65), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1006(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1007(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1008(.a(gate237inter12), .b(gate237inter1), .O(G742));

  xor2  gate645(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate646(.a(gate238inter0), .b(s_14), .O(gate238inter1));
  and2  gate647(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate648(.a(s_14), .O(gate238inter3));
  inv1  gate649(.a(s_15), .O(gate238inter4));
  nand2 gate650(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate651(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate652(.a(G257), .O(gate238inter7));
  inv1  gate653(.a(G709), .O(gate238inter8));
  nand2 gate654(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate655(.a(s_15), .b(gate238inter3), .O(gate238inter10));
  nor2  gate656(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate657(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate658(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate1723(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1724(.a(gate243inter0), .b(s_168), .O(gate243inter1));
  and2  gate1725(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1726(.a(s_168), .O(gate243inter3));
  inv1  gate1727(.a(s_169), .O(gate243inter4));
  nand2 gate1728(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1729(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1730(.a(G245), .O(gate243inter7));
  inv1  gate1731(.a(G733), .O(gate243inter8));
  nand2 gate1732(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1733(.a(s_169), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1734(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1735(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1736(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate869(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate870(.a(gate245inter0), .b(s_46), .O(gate245inter1));
  and2  gate871(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate872(.a(s_46), .O(gate245inter3));
  inv1  gate873(.a(s_47), .O(gate245inter4));
  nand2 gate874(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate875(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate876(.a(G248), .O(gate245inter7));
  inv1  gate877(.a(G736), .O(gate245inter8));
  nand2 gate878(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate879(.a(s_47), .b(gate245inter3), .O(gate245inter10));
  nor2  gate880(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate881(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate882(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate1023(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate1024(.a(gate249inter0), .b(s_68), .O(gate249inter1));
  and2  gate1025(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate1026(.a(s_68), .O(gate249inter3));
  inv1  gate1027(.a(s_69), .O(gate249inter4));
  nand2 gate1028(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate1029(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate1030(.a(G254), .O(gate249inter7));
  inv1  gate1031(.a(G742), .O(gate249inter8));
  nand2 gate1032(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate1033(.a(s_69), .b(gate249inter3), .O(gate249inter10));
  nor2  gate1034(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate1035(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate1036(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate1275(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate1276(.a(gate252inter0), .b(s_104), .O(gate252inter1));
  and2  gate1277(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate1278(.a(s_104), .O(gate252inter3));
  inv1  gate1279(.a(s_105), .O(gate252inter4));
  nand2 gate1280(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate1281(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate1282(.a(G709), .O(gate252inter7));
  inv1  gate1283(.a(G745), .O(gate252inter8));
  nand2 gate1284(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate1285(.a(s_105), .b(gate252inter3), .O(gate252inter10));
  nor2  gate1286(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate1287(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate1288(.a(gate252inter12), .b(gate252inter1), .O(G765));

  xor2  gate1359(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate1360(.a(gate253inter0), .b(s_116), .O(gate253inter1));
  and2  gate1361(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate1362(.a(s_116), .O(gate253inter3));
  inv1  gate1363(.a(s_117), .O(gate253inter4));
  nand2 gate1364(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate1365(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate1366(.a(G260), .O(gate253inter7));
  inv1  gate1367(.a(G748), .O(gate253inter8));
  nand2 gate1368(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate1369(.a(s_117), .b(gate253inter3), .O(gate253inter10));
  nor2  gate1370(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate1371(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate1372(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate1415(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate1416(.a(gate262inter0), .b(s_124), .O(gate262inter1));
  and2  gate1417(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate1418(.a(s_124), .O(gate262inter3));
  inv1  gate1419(.a(s_125), .O(gate262inter4));
  nand2 gate1420(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate1421(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate1422(.a(G764), .O(gate262inter7));
  inv1  gate1423(.a(G765), .O(gate262inter8));
  nand2 gate1424(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate1425(.a(s_125), .b(gate262inter3), .O(gate262inter10));
  nor2  gate1426(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate1427(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate1428(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate1191(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate1192(.a(gate266inter0), .b(s_92), .O(gate266inter1));
  and2  gate1193(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate1194(.a(s_92), .O(gate266inter3));
  inv1  gate1195(.a(s_93), .O(gate266inter4));
  nand2 gate1196(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate1197(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate1198(.a(G645), .O(gate266inter7));
  inv1  gate1199(.a(G773), .O(gate266inter8));
  nand2 gate1200(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate1201(.a(s_93), .b(gate266inter3), .O(gate266inter10));
  nor2  gate1202(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate1203(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate1204(.a(gate266inter12), .b(gate266inter1), .O(G797));

  xor2  gate1471(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate1472(.a(gate267inter0), .b(s_132), .O(gate267inter1));
  and2  gate1473(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate1474(.a(s_132), .O(gate267inter3));
  inv1  gate1475(.a(s_133), .O(gate267inter4));
  nand2 gate1476(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate1477(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate1478(.a(G648), .O(gate267inter7));
  inv1  gate1479(.a(G776), .O(gate267inter8));
  nand2 gate1480(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate1481(.a(s_133), .b(gate267inter3), .O(gate267inter10));
  nor2  gate1482(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate1483(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate1484(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );

  xor2  gate1709(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate1710(.a(gate273inter0), .b(s_166), .O(gate273inter1));
  and2  gate1711(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate1712(.a(s_166), .O(gate273inter3));
  inv1  gate1713(.a(s_167), .O(gate273inter4));
  nand2 gate1714(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate1715(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate1716(.a(G642), .O(gate273inter7));
  inv1  gate1717(.a(G794), .O(gate273inter8));
  nand2 gate1718(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate1719(.a(s_167), .b(gate273inter3), .O(gate273inter10));
  nor2  gate1720(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate1721(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate1722(.a(gate273inter12), .b(gate273inter1), .O(G818));
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate617(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate618(.a(gate278inter0), .b(s_10), .O(gate278inter1));
  and2  gate619(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate620(.a(s_10), .O(gate278inter3));
  inv1  gate621(.a(s_11), .O(gate278inter4));
  nand2 gate622(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate623(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate624(.a(G776), .O(gate278inter7));
  inv1  gate625(.a(G800), .O(gate278inter8));
  nand2 gate626(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate627(.a(s_11), .b(gate278inter3), .O(gate278inter10));
  nor2  gate628(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate629(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate630(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate715(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate716(.a(gate280inter0), .b(s_24), .O(gate280inter1));
  and2  gate717(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate718(.a(s_24), .O(gate280inter3));
  inv1  gate719(.a(s_25), .O(gate280inter4));
  nand2 gate720(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate721(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate722(.a(G779), .O(gate280inter7));
  inv1  gate723(.a(G803), .O(gate280inter8));
  nand2 gate724(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate725(.a(s_25), .b(gate280inter3), .O(gate280inter10));
  nor2  gate726(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate727(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate728(.a(gate280inter12), .b(gate280inter1), .O(G825));
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate757(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate758(.a(gate286inter0), .b(s_30), .O(gate286inter1));
  and2  gate759(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate760(.a(s_30), .O(gate286inter3));
  inv1  gate761(.a(s_31), .O(gate286inter4));
  nand2 gate762(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate763(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate764(.a(G788), .O(gate286inter7));
  inv1  gate765(.a(G812), .O(gate286inter8));
  nand2 gate766(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate767(.a(s_31), .b(gate286inter3), .O(gate286inter10));
  nor2  gate768(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate769(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate770(.a(gate286inter12), .b(gate286inter1), .O(G831));
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate1457(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate1458(.a(gate291inter0), .b(s_130), .O(gate291inter1));
  and2  gate1459(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate1460(.a(s_130), .O(gate291inter3));
  inv1  gate1461(.a(s_131), .O(gate291inter4));
  nand2 gate1462(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate1463(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate1464(.a(G822), .O(gate291inter7));
  inv1  gate1465(.a(G823), .O(gate291inter8));
  nand2 gate1466(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate1467(.a(s_131), .b(gate291inter3), .O(gate291inter10));
  nor2  gate1468(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate1469(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate1470(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate813(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate814(.a(gate293inter0), .b(s_38), .O(gate293inter1));
  and2  gate815(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate816(.a(s_38), .O(gate293inter3));
  inv1  gate817(.a(s_39), .O(gate293inter4));
  nand2 gate818(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate819(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate820(.a(G828), .O(gate293inter7));
  inv1  gate821(.a(G829), .O(gate293inter8));
  nand2 gate822(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate823(.a(s_39), .b(gate293inter3), .O(gate293inter10));
  nor2  gate824(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate825(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate826(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate1261(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate1262(.a(gate388inter0), .b(s_102), .O(gate388inter1));
  and2  gate1263(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate1264(.a(s_102), .O(gate388inter3));
  inv1  gate1265(.a(s_103), .O(gate388inter4));
  nand2 gate1266(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate1267(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate1268(.a(G2), .O(gate388inter7));
  inv1  gate1269(.a(G1039), .O(gate388inter8));
  nand2 gate1270(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate1271(.a(s_103), .b(gate388inter3), .O(gate388inter10));
  nor2  gate1272(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate1273(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate1274(.a(gate388inter12), .b(gate388inter1), .O(G1135));

  xor2  gate1653(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate1654(.a(gate389inter0), .b(s_158), .O(gate389inter1));
  and2  gate1655(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate1656(.a(s_158), .O(gate389inter3));
  inv1  gate1657(.a(s_159), .O(gate389inter4));
  nand2 gate1658(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate1659(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate1660(.a(G3), .O(gate389inter7));
  inv1  gate1661(.a(G1042), .O(gate389inter8));
  nand2 gate1662(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate1663(.a(s_159), .b(gate389inter3), .O(gate389inter10));
  nor2  gate1664(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate1665(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate1666(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate1107(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate1108(.a(gate391inter0), .b(s_80), .O(gate391inter1));
  and2  gate1109(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate1110(.a(s_80), .O(gate391inter3));
  inv1  gate1111(.a(s_81), .O(gate391inter4));
  nand2 gate1112(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate1113(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate1114(.a(G5), .O(gate391inter7));
  inv1  gate1115(.a(G1048), .O(gate391inter8));
  nand2 gate1116(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate1117(.a(s_81), .b(gate391inter3), .O(gate391inter10));
  nor2  gate1118(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate1119(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate1120(.a(gate391inter12), .b(gate391inter1), .O(G1144));

  xor2  gate547(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate548(.a(gate392inter0), .b(s_0), .O(gate392inter1));
  and2  gate549(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate550(.a(s_0), .O(gate392inter3));
  inv1  gate551(.a(s_1), .O(gate392inter4));
  nand2 gate552(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate553(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate554(.a(G6), .O(gate392inter7));
  inv1  gate555(.a(G1051), .O(gate392inter8));
  nand2 gate556(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate557(.a(s_1), .b(gate392inter3), .O(gate392inter10));
  nor2  gate558(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate559(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate560(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate967(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate968(.a(gate394inter0), .b(s_60), .O(gate394inter1));
  and2  gate969(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate970(.a(s_60), .O(gate394inter3));
  inv1  gate971(.a(s_61), .O(gate394inter4));
  nand2 gate972(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate973(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate974(.a(G8), .O(gate394inter7));
  inv1  gate975(.a(G1057), .O(gate394inter8));
  nand2 gate976(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate977(.a(s_61), .b(gate394inter3), .O(gate394inter10));
  nor2  gate978(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate979(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate980(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate1835(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate1836(.a(gate397inter0), .b(s_184), .O(gate397inter1));
  and2  gate1837(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate1838(.a(s_184), .O(gate397inter3));
  inv1  gate1839(.a(s_185), .O(gate397inter4));
  nand2 gate1840(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate1841(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate1842(.a(G11), .O(gate397inter7));
  inv1  gate1843(.a(G1066), .O(gate397inter8));
  nand2 gate1844(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate1845(.a(s_185), .b(gate397inter3), .O(gate397inter10));
  nor2  gate1846(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate1847(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate1848(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate799(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate800(.a(gate399inter0), .b(s_36), .O(gate399inter1));
  and2  gate801(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate802(.a(s_36), .O(gate399inter3));
  inv1  gate803(.a(s_37), .O(gate399inter4));
  nand2 gate804(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate805(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate806(.a(G13), .O(gate399inter7));
  inv1  gate807(.a(G1072), .O(gate399inter8));
  nand2 gate808(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate809(.a(s_37), .b(gate399inter3), .O(gate399inter10));
  nor2  gate810(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate811(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate812(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate1009(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate1010(.a(gate406inter0), .b(s_66), .O(gate406inter1));
  and2  gate1011(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate1012(.a(s_66), .O(gate406inter3));
  inv1  gate1013(.a(s_67), .O(gate406inter4));
  nand2 gate1014(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate1015(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate1016(.a(G20), .O(gate406inter7));
  inv1  gate1017(.a(G1093), .O(gate406inter8));
  nand2 gate1018(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate1019(.a(s_67), .b(gate406inter3), .O(gate406inter10));
  nor2  gate1020(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate1021(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate1022(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate785(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate786(.a(gate410inter0), .b(s_34), .O(gate410inter1));
  and2  gate787(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate788(.a(s_34), .O(gate410inter3));
  inv1  gate789(.a(s_35), .O(gate410inter4));
  nand2 gate790(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate791(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate792(.a(G24), .O(gate410inter7));
  inv1  gate793(.a(G1105), .O(gate410inter8));
  nand2 gate794(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate795(.a(s_35), .b(gate410inter3), .O(gate410inter10));
  nor2  gate796(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate797(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate798(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );

  xor2  gate1639(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate1640(.a(gate414inter0), .b(s_156), .O(gate414inter1));
  and2  gate1641(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate1642(.a(s_156), .O(gate414inter3));
  inv1  gate1643(.a(s_157), .O(gate414inter4));
  nand2 gate1644(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate1645(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate1646(.a(G28), .O(gate414inter7));
  inv1  gate1647(.a(G1117), .O(gate414inter8));
  nand2 gate1648(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate1649(.a(s_157), .b(gate414inter3), .O(gate414inter10));
  nor2  gate1650(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate1651(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate1652(.a(gate414inter12), .b(gate414inter1), .O(G1213));
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );

  xor2  gate1289(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate1290(.a(gate423inter0), .b(s_106), .O(gate423inter1));
  and2  gate1291(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate1292(.a(s_106), .O(gate423inter3));
  inv1  gate1293(.a(s_107), .O(gate423inter4));
  nand2 gate1294(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate1295(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate1296(.a(G3), .O(gate423inter7));
  inv1  gate1297(.a(G1138), .O(gate423inter8));
  nand2 gate1298(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate1299(.a(s_107), .b(gate423inter3), .O(gate423inter10));
  nor2  gate1300(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate1301(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate1302(.a(gate423inter12), .b(gate423inter1), .O(G1232));
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );

  xor2  gate575(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate576(.a(gate429inter0), .b(s_4), .O(gate429inter1));
  and2  gate577(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate578(.a(s_4), .O(gate429inter3));
  inv1  gate579(.a(s_5), .O(gate429inter4));
  nand2 gate580(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate581(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate582(.a(G6), .O(gate429inter7));
  inv1  gate583(.a(G1147), .O(gate429inter8));
  nand2 gate584(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate585(.a(s_5), .b(gate429inter3), .O(gate429inter10));
  nor2  gate586(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate587(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate588(.a(gate429inter12), .b(gate429inter1), .O(G1238));
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate1555(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate1556(.a(gate434inter0), .b(s_144), .O(gate434inter1));
  and2  gate1557(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate1558(.a(s_144), .O(gate434inter3));
  inv1  gate1559(.a(s_145), .O(gate434inter4));
  nand2 gate1560(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate1561(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate1562(.a(G1057), .O(gate434inter7));
  inv1  gate1563(.a(G1153), .O(gate434inter8));
  nand2 gate1564(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate1565(.a(s_145), .b(gate434inter3), .O(gate434inter10));
  nor2  gate1566(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate1567(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate1568(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate1611(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate1612(.a(gate437inter0), .b(s_152), .O(gate437inter1));
  and2  gate1613(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate1614(.a(s_152), .O(gate437inter3));
  inv1  gate1615(.a(s_153), .O(gate437inter4));
  nand2 gate1616(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate1617(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate1618(.a(G10), .O(gate437inter7));
  inv1  gate1619(.a(G1159), .O(gate437inter8));
  nand2 gate1620(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate1621(.a(s_153), .b(gate437inter3), .O(gate437inter10));
  nor2  gate1622(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate1623(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate1624(.a(gate437inter12), .b(gate437inter1), .O(G1246));

  xor2  gate1345(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate1346(.a(gate438inter0), .b(s_114), .O(gate438inter1));
  and2  gate1347(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate1348(.a(s_114), .O(gate438inter3));
  inv1  gate1349(.a(s_115), .O(gate438inter4));
  nand2 gate1350(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate1351(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate1352(.a(G1063), .O(gate438inter7));
  inv1  gate1353(.a(G1159), .O(gate438inter8));
  nand2 gate1354(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate1355(.a(s_115), .b(gate438inter3), .O(gate438inter10));
  nor2  gate1356(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate1357(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate1358(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate981(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate982(.a(gate444inter0), .b(s_62), .O(gate444inter1));
  and2  gate983(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate984(.a(s_62), .O(gate444inter3));
  inv1  gate985(.a(s_63), .O(gate444inter4));
  nand2 gate986(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate987(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate988(.a(G1072), .O(gate444inter7));
  inv1  gate989(.a(G1168), .O(gate444inter8));
  nand2 gate990(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate991(.a(s_63), .b(gate444inter3), .O(gate444inter10));
  nor2  gate992(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate993(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate994(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate603(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate604(.a(gate453inter0), .b(s_8), .O(gate453inter1));
  and2  gate605(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate606(.a(s_8), .O(gate453inter3));
  inv1  gate607(.a(s_9), .O(gate453inter4));
  nand2 gate608(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate609(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate610(.a(G18), .O(gate453inter7));
  inv1  gate611(.a(G1183), .O(gate453inter8));
  nand2 gate612(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate613(.a(s_9), .b(gate453inter3), .O(gate453inter10));
  nor2  gate614(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate615(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate616(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );

  xor2  gate673(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate674(.a(gate455inter0), .b(s_18), .O(gate455inter1));
  and2  gate675(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate676(.a(s_18), .O(gate455inter3));
  inv1  gate677(.a(s_19), .O(gate455inter4));
  nand2 gate678(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate679(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate680(.a(G19), .O(gate455inter7));
  inv1  gate681(.a(G1186), .O(gate455inter8));
  nand2 gate682(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate683(.a(s_19), .b(gate455inter3), .O(gate455inter10));
  nor2  gate684(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate685(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate686(.a(gate455inter12), .b(gate455inter1), .O(G1264));
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate1877(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate1878(.a(gate459inter0), .b(s_190), .O(gate459inter1));
  and2  gate1879(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate1880(.a(s_190), .O(gate459inter3));
  inv1  gate1881(.a(s_191), .O(gate459inter4));
  nand2 gate1882(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate1883(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate1884(.a(G21), .O(gate459inter7));
  inv1  gate1885(.a(G1192), .O(gate459inter8));
  nand2 gate1886(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate1887(.a(s_191), .b(gate459inter3), .O(gate459inter10));
  nor2  gate1888(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate1889(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate1890(.a(gate459inter12), .b(gate459inter1), .O(G1268));

  xor2  gate1849(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate1850(.a(gate460inter0), .b(s_186), .O(gate460inter1));
  and2  gate1851(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate1852(.a(s_186), .O(gate460inter3));
  inv1  gate1853(.a(s_187), .O(gate460inter4));
  nand2 gate1854(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate1855(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate1856(.a(G1096), .O(gate460inter7));
  inv1  gate1857(.a(G1192), .O(gate460inter8));
  nand2 gate1858(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate1859(.a(s_187), .b(gate460inter3), .O(gate460inter10));
  nor2  gate1860(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate1861(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate1862(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );

  xor2  gate897(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate898(.a(gate462inter0), .b(s_50), .O(gate462inter1));
  and2  gate899(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate900(.a(s_50), .O(gate462inter3));
  inv1  gate901(.a(s_51), .O(gate462inter4));
  nand2 gate902(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate903(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate904(.a(G1099), .O(gate462inter7));
  inv1  gate905(.a(G1195), .O(gate462inter8));
  nand2 gate906(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate907(.a(s_51), .b(gate462inter3), .O(gate462inter10));
  nor2  gate908(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate909(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate910(.a(gate462inter12), .b(gate462inter1), .O(G1271));

  xor2  gate925(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate926(.a(gate463inter0), .b(s_54), .O(gate463inter1));
  and2  gate927(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate928(.a(s_54), .O(gate463inter3));
  inv1  gate929(.a(s_55), .O(gate463inter4));
  nand2 gate930(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate931(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate932(.a(G23), .O(gate463inter7));
  inv1  gate933(.a(G1198), .O(gate463inter8));
  nand2 gate934(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate935(.a(s_55), .b(gate463inter3), .O(gate463inter10));
  nor2  gate936(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate937(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate938(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate743(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate744(.a(gate467inter0), .b(s_28), .O(gate467inter1));
  and2  gate745(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate746(.a(s_28), .O(gate467inter3));
  inv1  gate747(.a(s_29), .O(gate467inter4));
  nand2 gate748(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate749(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate750(.a(G25), .O(gate467inter7));
  inv1  gate751(.a(G1204), .O(gate467inter8));
  nand2 gate752(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate753(.a(s_29), .b(gate467inter3), .O(gate467inter10));
  nor2  gate754(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate755(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate756(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );

  xor2  gate1429(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate1430(.a(gate473inter0), .b(s_126), .O(gate473inter1));
  and2  gate1431(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate1432(.a(s_126), .O(gate473inter3));
  inv1  gate1433(.a(s_127), .O(gate473inter4));
  nand2 gate1434(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate1435(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate1436(.a(G28), .O(gate473inter7));
  inv1  gate1437(.a(G1213), .O(gate473inter8));
  nand2 gate1438(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate1439(.a(s_127), .b(gate473inter3), .O(gate473inter10));
  nor2  gate1440(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate1441(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate1442(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate589(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate590(.a(gate480inter0), .b(s_6), .O(gate480inter1));
  and2  gate591(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate592(.a(s_6), .O(gate480inter3));
  inv1  gate593(.a(s_7), .O(gate480inter4));
  nand2 gate594(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate595(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate596(.a(G1126), .O(gate480inter7));
  inv1  gate597(.a(G1222), .O(gate480inter8));
  nand2 gate598(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate599(.a(s_7), .b(gate480inter3), .O(gate480inter10));
  nor2  gate600(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate601(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate602(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );

  xor2  gate1541(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate1542(.a(gate498inter0), .b(s_142), .O(gate498inter1));
  and2  gate1543(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate1544(.a(s_142), .O(gate498inter3));
  inv1  gate1545(.a(s_143), .O(gate498inter4));
  nand2 gate1546(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate1547(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate1548(.a(G1258), .O(gate498inter7));
  inv1  gate1549(.a(G1259), .O(gate498inter8));
  nand2 gate1550(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate1551(.a(s_143), .b(gate498inter3), .O(gate498inter10));
  nor2  gate1552(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate1553(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate1554(.a(gate498inter12), .b(gate498inter1), .O(G1307));
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate1079(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate1080(.a(gate500inter0), .b(s_76), .O(gate500inter1));
  and2  gate1081(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate1082(.a(s_76), .O(gate500inter3));
  inv1  gate1083(.a(s_77), .O(gate500inter4));
  nand2 gate1084(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate1085(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate1086(.a(G1262), .O(gate500inter7));
  inv1  gate1087(.a(G1263), .O(gate500inter8));
  nand2 gate1088(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate1089(.a(s_77), .b(gate500inter3), .O(gate500inter10));
  nor2  gate1090(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate1091(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate1092(.a(gate500inter12), .b(gate500inter1), .O(G1309));
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate1737(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate1738(.a(gate506inter0), .b(s_170), .O(gate506inter1));
  and2  gate1739(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate1740(.a(s_170), .O(gate506inter3));
  inv1  gate1741(.a(s_171), .O(gate506inter4));
  nand2 gate1742(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate1743(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate1744(.a(G1274), .O(gate506inter7));
  inv1  gate1745(.a(G1275), .O(gate506inter8));
  nand2 gate1746(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate1747(.a(s_171), .b(gate506inter3), .O(gate506inter10));
  nor2  gate1748(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate1749(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate1750(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate701(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate702(.a(gate508inter0), .b(s_22), .O(gate508inter1));
  and2  gate703(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate704(.a(s_22), .O(gate508inter3));
  inv1  gate705(.a(s_23), .O(gate508inter4));
  nand2 gate706(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate707(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate708(.a(G1278), .O(gate508inter7));
  inv1  gate709(.a(G1279), .O(gate508inter8));
  nand2 gate710(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate711(.a(s_23), .b(gate508inter3), .O(gate508inter10));
  nor2  gate712(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate713(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate714(.a(gate508inter12), .b(gate508inter1), .O(G1317));

  xor2  gate1233(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate1234(.a(gate509inter0), .b(s_98), .O(gate509inter1));
  and2  gate1235(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate1236(.a(s_98), .O(gate509inter3));
  inv1  gate1237(.a(s_99), .O(gate509inter4));
  nand2 gate1238(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate1239(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate1240(.a(G1280), .O(gate509inter7));
  inv1  gate1241(.a(G1281), .O(gate509inter8));
  nand2 gate1242(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate1243(.a(s_99), .b(gate509inter3), .O(gate509inter10));
  nor2  gate1244(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate1245(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate1246(.a(gate509inter12), .b(gate509inter1), .O(G1318));

  xor2  gate1163(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate1164(.a(gate510inter0), .b(s_88), .O(gate510inter1));
  and2  gate1165(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate1166(.a(s_88), .O(gate510inter3));
  inv1  gate1167(.a(s_89), .O(gate510inter4));
  nand2 gate1168(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate1169(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate1170(.a(G1282), .O(gate510inter7));
  inv1  gate1171(.a(G1283), .O(gate510inter8));
  nand2 gate1172(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate1173(.a(s_89), .b(gate510inter3), .O(gate510inter10));
  nor2  gate1174(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate1175(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate1176(.a(gate510inter12), .b(gate510inter1), .O(G1319));

  xor2  gate1443(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate1444(.a(gate511inter0), .b(s_128), .O(gate511inter1));
  and2  gate1445(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate1446(.a(s_128), .O(gate511inter3));
  inv1  gate1447(.a(s_129), .O(gate511inter4));
  nand2 gate1448(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate1449(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate1450(.a(G1284), .O(gate511inter7));
  inv1  gate1451(.a(G1285), .O(gate511inter8));
  nand2 gate1452(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate1453(.a(s_129), .b(gate511inter3), .O(gate511inter10));
  nor2  gate1454(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate1455(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate1456(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule