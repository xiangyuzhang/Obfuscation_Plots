module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate1429(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate1430(.a(gate9inter0), .b(s_126), .O(gate9inter1));
  and2  gate1431(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate1432(.a(s_126), .O(gate9inter3));
  inv1  gate1433(.a(s_127), .O(gate9inter4));
  nand2 gate1434(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate1435(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate1436(.a(G1), .O(gate9inter7));
  inv1  gate1437(.a(G2), .O(gate9inter8));
  nand2 gate1438(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate1439(.a(s_127), .b(gate9inter3), .O(gate9inter10));
  nor2  gate1440(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate1441(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate1442(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate631(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate632(.a(gate11inter0), .b(s_12), .O(gate11inter1));
  and2  gate633(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate634(.a(s_12), .O(gate11inter3));
  inv1  gate635(.a(s_13), .O(gate11inter4));
  nand2 gate636(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate637(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate638(.a(G5), .O(gate11inter7));
  inv1  gate639(.a(G6), .O(gate11inter8));
  nand2 gate640(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate641(.a(s_13), .b(gate11inter3), .O(gate11inter10));
  nor2  gate642(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate643(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate644(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );

  xor2  gate1135(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate1136(.a(gate14inter0), .b(s_84), .O(gate14inter1));
  and2  gate1137(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate1138(.a(s_84), .O(gate14inter3));
  inv1  gate1139(.a(s_85), .O(gate14inter4));
  nand2 gate1140(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate1141(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate1142(.a(G11), .O(gate14inter7));
  inv1  gate1143(.a(G12), .O(gate14inter8));
  nand2 gate1144(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate1145(.a(s_85), .b(gate14inter3), .O(gate14inter10));
  nor2  gate1146(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate1147(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate1148(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate1653(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate1654(.a(gate20inter0), .b(s_158), .O(gate20inter1));
  and2  gate1655(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate1656(.a(s_158), .O(gate20inter3));
  inv1  gate1657(.a(s_159), .O(gate20inter4));
  nand2 gate1658(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate1659(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate1660(.a(G23), .O(gate20inter7));
  inv1  gate1661(.a(G24), .O(gate20inter8));
  nand2 gate1662(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate1663(.a(s_159), .b(gate20inter3), .O(gate20inter10));
  nor2  gate1664(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate1665(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate1666(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate1079(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate1080(.a(gate26inter0), .b(s_76), .O(gate26inter1));
  and2  gate1081(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate1082(.a(s_76), .O(gate26inter3));
  inv1  gate1083(.a(s_77), .O(gate26inter4));
  nand2 gate1084(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate1085(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate1086(.a(G9), .O(gate26inter7));
  inv1  gate1087(.a(G13), .O(gate26inter8));
  nand2 gate1088(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate1089(.a(s_77), .b(gate26inter3), .O(gate26inter10));
  nor2  gate1090(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate1091(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate1092(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate1485(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate1486(.a(gate33inter0), .b(s_134), .O(gate33inter1));
  and2  gate1487(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate1488(.a(s_134), .O(gate33inter3));
  inv1  gate1489(.a(s_135), .O(gate33inter4));
  nand2 gate1490(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate1491(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate1492(.a(G17), .O(gate33inter7));
  inv1  gate1493(.a(G21), .O(gate33inter8));
  nand2 gate1494(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate1495(.a(s_135), .b(gate33inter3), .O(gate33inter10));
  nor2  gate1496(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate1497(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate1498(.a(gate33inter12), .b(gate33inter1), .O(G338));
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );

  xor2  gate1037(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate1038(.a(gate42inter0), .b(s_70), .O(gate42inter1));
  and2  gate1039(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate1040(.a(s_70), .O(gate42inter3));
  inv1  gate1041(.a(s_71), .O(gate42inter4));
  nand2 gate1042(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate1043(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate1044(.a(G2), .O(gate42inter7));
  inv1  gate1045(.a(G266), .O(gate42inter8));
  nand2 gate1046(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate1047(.a(s_71), .b(gate42inter3), .O(gate42inter10));
  nor2  gate1048(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate1049(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate1050(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate967(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate968(.a(gate44inter0), .b(s_60), .O(gate44inter1));
  and2  gate969(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate970(.a(s_60), .O(gate44inter3));
  inv1  gate971(.a(s_61), .O(gate44inter4));
  nand2 gate972(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate973(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate974(.a(G4), .O(gate44inter7));
  inv1  gate975(.a(G269), .O(gate44inter8));
  nand2 gate976(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate977(.a(s_61), .b(gate44inter3), .O(gate44inter10));
  nor2  gate978(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate979(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate980(.a(gate44inter12), .b(gate44inter1), .O(G365));

  xor2  gate799(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate800(.a(gate45inter0), .b(s_36), .O(gate45inter1));
  and2  gate801(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate802(.a(s_36), .O(gate45inter3));
  inv1  gate803(.a(s_37), .O(gate45inter4));
  nand2 gate804(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate805(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate806(.a(G5), .O(gate45inter7));
  inv1  gate807(.a(G272), .O(gate45inter8));
  nand2 gate808(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate809(.a(s_37), .b(gate45inter3), .O(gate45inter10));
  nor2  gate810(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate811(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate812(.a(gate45inter12), .b(gate45inter1), .O(G366));
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate1569(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate1570(.a(gate52inter0), .b(s_146), .O(gate52inter1));
  and2  gate1571(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate1572(.a(s_146), .O(gate52inter3));
  inv1  gate1573(.a(s_147), .O(gate52inter4));
  nand2 gate1574(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate1575(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate1576(.a(G12), .O(gate52inter7));
  inv1  gate1577(.a(G281), .O(gate52inter8));
  nand2 gate1578(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate1579(.a(s_147), .b(gate52inter3), .O(gate52inter10));
  nor2  gate1580(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate1581(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate1582(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );

  xor2  gate1807(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate1808(.a(gate56inter0), .b(s_180), .O(gate56inter1));
  and2  gate1809(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate1810(.a(s_180), .O(gate56inter3));
  inv1  gate1811(.a(s_181), .O(gate56inter4));
  nand2 gate1812(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate1813(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate1814(.a(G16), .O(gate56inter7));
  inv1  gate1815(.a(G287), .O(gate56inter8));
  nand2 gate1816(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate1817(.a(s_181), .b(gate56inter3), .O(gate56inter10));
  nor2  gate1818(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate1819(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate1820(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate1401(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate1402(.a(gate62inter0), .b(s_122), .O(gate62inter1));
  and2  gate1403(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate1404(.a(s_122), .O(gate62inter3));
  inv1  gate1405(.a(s_123), .O(gate62inter4));
  nand2 gate1406(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate1407(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate1408(.a(G22), .O(gate62inter7));
  inv1  gate1409(.a(G296), .O(gate62inter8));
  nand2 gate1410(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate1411(.a(s_123), .b(gate62inter3), .O(gate62inter10));
  nor2  gate1412(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate1413(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate1414(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate1275(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate1276(.a(gate70inter0), .b(s_104), .O(gate70inter1));
  and2  gate1277(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate1278(.a(s_104), .O(gate70inter3));
  inv1  gate1279(.a(s_105), .O(gate70inter4));
  nand2 gate1280(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate1281(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate1282(.a(G30), .O(gate70inter7));
  inv1  gate1283(.a(G308), .O(gate70inter8));
  nand2 gate1284(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate1285(.a(s_105), .b(gate70inter3), .O(gate70inter10));
  nor2  gate1286(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate1287(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate1288(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate743(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate744(.a(gate75inter0), .b(s_28), .O(gate75inter1));
  and2  gate745(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate746(.a(s_28), .O(gate75inter3));
  inv1  gate747(.a(s_29), .O(gate75inter4));
  nand2 gate748(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate749(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate750(.a(G9), .O(gate75inter7));
  inv1  gate751(.a(G317), .O(gate75inter8));
  nand2 gate752(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate753(.a(s_29), .b(gate75inter3), .O(gate75inter10));
  nor2  gate754(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate755(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate756(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate1611(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate1612(.a(gate80inter0), .b(s_152), .O(gate80inter1));
  and2  gate1613(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate1614(.a(s_152), .O(gate80inter3));
  inv1  gate1615(.a(s_153), .O(gate80inter4));
  nand2 gate1616(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate1617(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate1618(.a(G14), .O(gate80inter7));
  inv1  gate1619(.a(G323), .O(gate80inter8));
  nand2 gate1620(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate1621(.a(s_153), .b(gate80inter3), .O(gate80inter10));
  nor2  gate1622(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate1623(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate1624(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate925(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate926(.a(gate90inter0), .b(s_54), .O(gate90inter1));
  and2  gate927(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate928(.a(s_54), .O(gate90inter3));
  inv1  gate929(.a(s_55), .O(gate90inter4));
  nand2 gate930(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate931(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate932(.a(G21), .O(gate90inter7));
  inv1  gate933(.a(G338), .O(gate90inter8));
  nand2 gate934(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate935(.a(s_55), .b(gate90inter3), .O(gate90inter10));
  nor2  gate936(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate937(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate938(.a(gate90inter12), .b(gate90inter1), .O(G411));
nand2 gate91( .a(G25), .b(G341), .O(G412) );

  xor2  gate673(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate674(.a(gate92inter0), .b(s_18), .O(gate92inter1));
  and2  gate675(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate676(.a(s_18), .O(gate92inter3));
  inv1  gate677(.a(s_19), .O(gate92inter4));
  nand2 gate678(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate679(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate680(.a(G29), .O(gate92inter7));
  inv1  gate681(.a(G341), .O(gate92inter8));
  nand2 gate682(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate683(.a(s_19), .b(gate92inter3), .O(gate92inter10));
  nor2  gate684(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate685(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate686(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate813(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate814(.a(gate112inter0), .b(s_38), .O(gate112inter1));
  and2  gate815(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate816(.a(s_38), .O(gate112inter3));
  inv1  gate817(.a(s_39), .O(gate112inter4));
  nand2 gate818(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate819(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate820(.a(G376), .O(gate112inter7));
  inv1  gate821(.a(G377), .O(gate112inter8));
  nand2 gate822(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate823(.a(s_39), .b(gate112inter3), .O(gate112inter10));
  nor2  gate824(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate825(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate826(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate1205(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate1206(.a(gate116inter0), .b(s_94), .O(gate116inter1));
  and2  gate1207(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate1208(.a(s_94), .O(gate116inter3));
  inv1  gate1209(.a(s_95), .O(gate116inter4));
  nand2 gate1210(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate1211(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate1212(.a(G384), .O(gate116inter7));
  inv1  gate1213(.a(G385), .O(gate116inter8));
  nand2 gate1214(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate1215(.a(s_95), .b(gate116inter3), .O(gate116inter10));
  nor2  gate1216(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate1217(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate1218(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate1709(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate1710(.a(gate124inter0), .b(s_166), .O(gate124inter1));
  and2  gate1711(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate1712(.a(s_166), .O(gate124inter3));
  inv1  gate1713(.a(s_167), .O(gate124inter4));
  nand2 gate1714(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate1715(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate1716(.a(G400), .O(gate124inter7));
  inv1  gate1717(.a(G401), .O(gate124inter8));
  nand2 gate1718(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate1719(.a(s_167), .b(gate124inter3), .O(gate124inter10));
  nor2  gate1720(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate1721(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate1722(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );

  xor2  gate1597(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate1598(.a(gate140inter0), .b(s_150), .O(gate140inter1));
  and2  gate1599(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate1600(.a(s_150), .O(gate140inter3));
  inv1  gate1601(.a(s_151), .O(gate140inter4));
  nand2 gate1602(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate1603(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate1604(.a(G444), .O(gate140inter7));
  inv1  gate1605(.a(G447), .O(gate140inter8));
  nand2 gate1606(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate1607(.a(s_151), .b(gate140inter3), .O(gate140inter10));
  nor2  gate1608(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate1609(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate1610(.a(gate140inter12), .b(gate140inter1), .O(G531));
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );

  xor2  gate1583(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate1584(.a(gate146inter0), .b(s_148), .O(gate146inter1));
  and2  gate1585(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate1586(.a(s_148), .O(gate146inter3));
  inv1  gate1587(.a(s_149), .O(gate146inter4));
  nand2 gate1588(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate1589(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate1590(.a(G480), .O(gate146inter7));
  inv1  gate1591(.a(G483), .O(gate146inter8));
  nand2 gate1592(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate1593(.a(s_149), .b(gate146inter3), .O(gate146inter10));
  nor2  gate1594(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate1595(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate1596(.a(gate146inter12), .b(gate146inter1), .O(G549));
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate1317(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate1318(.a(gate150inter0), .b(s_110), .O(gate150inter1));
  and2  gate1319(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate1320(.a(s_110), .O(gate150inter3));
  inv1  gate1321(.a(s_111), .O(gate150inter4));
  nand2 gate1322(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate1323(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate1324(.a(G504), .O(gate150inter7));
  inv1  gate1325(.a(G507), .O(gate150inter8));
  nand2 gate1326(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate1327(.a(s_111), .b(gate150inter3), .O(gate150inter10));
  nor2  gate1328(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate1329(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate1330(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate939(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate940(.a(gate155inter0), .b(s_56), .O(gate155inter1));
  and2  gate941(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate942(.a(s_56), .O(gate155inter3));
  inv1  gate943(.a(s_57), .O(gate155inter4));
  nand2 gate944(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate945(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate946(.a(G432), .O(gate155inter7));
  inv1  gate947(.a(G525), .O(gate155inter8));
  nand2 gate948(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate949(.a(s_57), .b(gate155inter3), .O(gate155inter10));
  nor2  gate950(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate951(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate952(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate1695(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate1696(.a(gate160inter0), .b(s_164), .O(gate160inter1));
  and2  gate1697(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate1698(.a(s_164), .O(gate160inter3));
  inv1  gate1699(.a(s_165), .O(gate160inter4));
  nand2 gate1700(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate1701(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate1702(.a(G447), .O(gate160inter7));
  inv1  gate1703(.a(G531), .O(gate160inter8));
  nand2 gate1704(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate1705(.a(s_165), .b(gate160inter3), .O(gate160inter10));
  nor2  gate1706(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate1707(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate1708(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );

  xor2  gate561(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate562(.a(gate169inter0), .b(s_2), .O(gate169inter1));
  and2  gate563(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate564(.a(s_2), .O(gate169inter3));
  inv1  gate565(.a(s_3), .O(gate169inter4));
  nand2 gate566(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate567(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate568(.a(G474), .O(gate169inter7));
  inv1  gate569(.a(G546), .O(gate169inter8));
  nand2 gate570(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate571(.a(s_3), .b(gate169inter3), .O(gate169inter10));
  nor2  gate572(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate573(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate574(.a(gate169inter12), .b(gate169inter1), .O(G586));
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate1261(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate1262(.a(gate174inter0), .b(s_102), .O(gate174inter1));
  and2  gate1263(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate1264(.a(s_102), .O(gate174inter3));
  inv1  gate1265(.a(s_103), .O(gate174inter4));
  nand2 gate1266(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate1267(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate1268(.a(G489), .O(gate174inter7));
  inv1  gate1269(.a(G552), .O(gate174inter8));
  nand2 gate1270(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate1271(.a(s_103), .b(gate174inter3), .O(gate174inter10));
  nor2  gate1272(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate1273(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate1274(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate603(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate604(.a(gate178inter0), .b(s_8), .O(gate178inter1));
  and2  gate605(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate606(.a(s_8), .O(gate178inter3));
  inv1  gate607(.a(s_9), .O(gate178inter4));
  nand2 gate608(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate609(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate610(.a(G501), .O(gate178inter7));
  inv1  gate611(.a(G558), .O(gate178inter8));
  nand2 gate612(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate613(.a(s_9), .b(gate178inter3), .O(gate178inter10));
  nor2  gate614(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate615(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate616(.a(gate178inter12), .b(gate178inter1), .O(G595));
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate1359(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate1360(.a(gate187inter0), .b(s_116), .O(gate187inter1));
  and2  gate1361(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate1362(.a(s_116), .O(gate187inter3));
  inv1  gate1363(.a(s_117), .O(gate187inter4));
  nand2 gate1364(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate1365(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate1366(.a(G574), .O(gate187inter7));
  inv1  gate1367(.a(G575), .O(gate187inter8));
  nand2 gate1368(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate1369(.a(s_117), .b(gate187inter3), .O(gate187inter10));
  nor2  gate1370(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate1371(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate1372(.a(gate187inter12), .b(gate187inter1), .O(G612));

  xor2  gate1177(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate1178(.a(gate188inter0), .b(s_90), .O(gate188inter1));
  and2  gate1179(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate1180(.a(s_90), .O(gate188inter3));
  inv1  gate1181(.a(s_91), .O(gate188inter4));
  nand2 gate1182(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate1183(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate1184(.a(G576), .O(gate188inter7));
  inv1  gate1185(.a(G577), .O(gate188inter8));
  nand2 gate1186(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate1187(.a(s_91), .b(gate188inter3), .O(gate188inter10));
  nor2  gate1188(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate1189(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate1190(.a(gate188inter12), .b(gate188inter1), .O(G617));

  xor2  gate1373(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate1374(.a(gate189inter0), .b(s_118), .O(gate189inter1));
  and2  gate1375(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate1376(.a(s_118), .O(gate189inter3));
  inv1  gate1377(.a(s_119), .O(gate189inter4));
  nand2 gate1378(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate1379(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate1380(.a(G578), .O(gate189inter7));
  inv1  gate1381(.a(G579), .O(gate189inter8));
  nand2 gate1382(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate1383(.a(s_119), .b(gate189inter3), .O(gate189inter10));
  nor2  gate1384(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate1385(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate1386(.a(gate189inter12), .b(gate189inter1), .O(G622));
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate1023(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate1024(.a(gate193inter0), .b(s_68), .O(gate193inter1));
  and2  gate1025(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate1026(.a(s_68), .O(gate193inter3));
  inv1  gate1027(.a(s_69), .O(gate193inter4));
  nand2 gate1028(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate1029(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate1030(.a(G586), .O(gate193inter7));
  inv1  gate1031(.a(G587), .O(gate193inter8));
  nand2 gate1032(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate1033(.a(s_69), .b(gate193inter3), .O(gate193inter10));
  nor2  gate1034(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate1035(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate1036(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate1555(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate1556(.a(gate197inter0), .b(s_144), .O(gate197inter1));
  and2  gate1557(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate1558(.a(s_144), .O(gate197inter3));
  inv1  gate1559(.a(s_145), .O(gate197inter4));
  nand2 gate1560(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate1561(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate1562(.a(G594), .O(gate197inter7));
  inv1  gate1563(.a(G595), .O(gate197inter8));
  nand2 gate1564(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate1565(.a(s_145), .b(gate197inter3), .O(gate197inter10));
  nor2  gate1566(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate1567(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate1568(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );

  xor2  gate981(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate982(.a(gate202inter0), .b(s_62), .O(gate202inter1));
  and2  gate983(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate984(.a(s_62), .O(gate202inter3));
  inv1  gate985(.a(s_63), .O(gate202inter4));
  nand2 gate986(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate987(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate988(.a(G612), .O(gate202inter7));
  inv1  gate989(.a(G617), .O(gate202inter8));
  nand2 gate990(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate991(.a(s_63), .b(gate202inter3), .O(gate202inter10));
  nor2  gate992(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate993(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate994(.a(gate202inter12), .b(gate202inter1), .O(G669));

  xor2  gate1387(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate1388(.a(gate203inter0), .b(s_120), .O(gate203inter1));
  and2  gate1389(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate1390(.a(s_120), .O(gate203inter3));
  inv1  gate1391(.a(s_121), .O(gate203inter4));
  nand2 gate1392(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate1393(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate1394(.a(G602), .O(gate203inter7));
  inv1  gate1395(.a(G612), .O(gate203inter8));
  nand2 gate1396(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate1397(.a(s_121), .b(gate203inter3), .O(gate203inter10));
  nor2  gate1398(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate1399(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate1400(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );

  xor2  gate855(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate856(.a(gate209inter0), .b(s_44), .O(gate209inter1));
  and2  gate857(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate858(.a(s_44), .O(gate209inter3));
  inv1  gate859(.a(s_45), .O(gate209inter4));
  nand2 gate860(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate861(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate862(.a(G602), .O(gate209inter7));
  inv1  gate863(.a(G666), .O(gate209inter8));
  nand2 gate864(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate865(.a(s_45), .b(gate209inter3), .O(gate209inter10));
  nor2  gate866(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate867(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate868(.a(gate209inter12), .b(gate209inter1), .O(G690));

  xor2  gate1107(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate1108(.a(gate210inter0), .b(s_80), .O(gate210inter1));
  and2  gate1109(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate1110(.a(s_80), .O(gate210inter3));
  inv1  gate1111(.a(s_81), .O(gate210inter4));
  nand2 gate1112(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate1113(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate1114(.a(G607), .O(gate210inter7));
  inv1  gate1115(.a(G666), .O(gate210inter8));
  nand2 gate1116(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate1117(.a(s_81), .b(gate210inter3), .O(gate210inter10));
  nor2  gate1118(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate1119(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate1120(.a(gate210inter12), .b(gate210inter1), .O(G691));

  xor2  gate547(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate548(.a(gate211inter0), .b(s_0), .O(gate211inter1));
  and2  gate549(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate550(.a(s_0), .O(gate211inter3));
  inv1  gate551(.a(s_1), .O(gate211inter4));
  nand2 gate552(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate553(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate554(.a(G612), .O(gate211inter7));
  inv1  gate555(.a(G669), .O(gate211inter8));
  nand2 gate556(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate557(.a(s_1), .b(gate211inter3), .O(gate211inter10));
  nor2  gate558(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate559(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate560(.a(gate211inter12), .b(gate211inter1), .O(G692));

  xor2  gate1765(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate1766(.a(gate212inter0), .b(s_174), .O(gate212inter1));
  and2  gate1767(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate1768(.a(s_174), .O(gate212inter3));
  inv1  gate1769(.a(s_175), .O(gate212inter4));
  nand2 gate1770(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate1771(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate1772(.a(G617), .O(gate212inter7));
  inv1  gate1773(.a(G669), .O(gate212inter8));
  nand2 gate1774(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate1775(.a(s_175), .b(gate212inter3), .O(gate212inter10));
  nor2  gate1776(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate1777(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate1778(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );

  xor2  gate869(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate870(.a(gate221inter0), .b(s_46), .O(gate221inter1));
  and2  gate871(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate872(.a(s_46), .O(gate221inter3));
  inv1  gate873(.a(s_47), .O(gate221inter4));
  nand2 gate874(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate875(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate876(.a(G622), .O(gate221inter7));
  inv1  gate877(.a(G684), .O(gate221inter8));
  nand2 gate878(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate879(.a(s_47), .b(gate221inter3), .O(gate221inter10));
  nor2  gate880(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate881(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate882(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );

  xor2  gate1737(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate1738(.a(gate225inter0), .b(s_170), .O(gate225inter1));
  and2  gate1739(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate1740(.a(s_170), .O(gate225inter3));
  inv1  gate1741(.a(s_171), .O(gate225inter4));
  nand2 gate1742(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate1743(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate1744(.a(G690), .O(gate225inter7));
  inv1  gate1745(.a(G691), .O(gate225inter8));
  nand2 gate1746(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate1747(.a(s_171), .b(gate225inter3), .O(gate225inter10));
  nor2  gate1748(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate1749(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate1750(.a(gate225inter12), .b(gate225inter1), .O(G706));
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate841(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate842(.a(gate227inter0), .b(s_42), .O(gate227inter1));
  and2  gate843(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate844(.a(s_42), .O(gate227inter3));
  inv1  gate845(.a(s_43), .O(gate227inter4));
  nand2 gate846(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate847(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate848(.a(G694), .O(gate227inter7));
  inv1  gate849(.a(G695), .O(gate227inter8));
  nand2 gate850(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate851(.a(s_43), .b(gate227inter3), .O(gate227inter10));
  nor2  gate852(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate853(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate854(.a(gate227inter12), .b(gate227inter1), .O(G712));
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate1009(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate1010(.a(gate237inter0), .b(s_66), .O(gate237inter1));
  and2  gate1011(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate1012(.a(s_66), .O(gate237inter3));
  inv1  gate1013(.a(s_67), .O(gate237inter4));
  nand2 gate1014(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1015(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1016(.a(G254), .O(gate237inter7));
  inv1  gate1017(.a(G706), .O(gate237inter8));
  nand2 gate1018(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1019(.a(s_67), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1020(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1021(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1022(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );

  xor2  gate785(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate786(.a(gate242inter0), .b(s_34), .O(gate242inter1));
  and2  gate787(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate788(.a(s_34), .O(gate242inter3));
  inv1  gate789(.a(s_35), .O(gate242inter4));
  nand2 gate790(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate791(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate792(.a(G718), .O(gate242inter7));
  inv1  gate793(.a(G730), .O(gate242inter8));
  nand2 gate794(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate795(.a(s_35), .b(gate242inter3), .O(gate242inter10));
  nor2  gate796(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate797(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate798(.a(gate242inter12), .b(gate242inter1), .O(G755));
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate1149(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate1150(.a(gate245inter0), .b(s_86), .O(gate245inter1));
  and2  gate1151(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate1152(.a(s_86), .O(gate245inter3));
  inv1  gate1153(.a(s_87), .O(gate245inter4));
  nand2 gate1154(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate1155(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate1156(.a(G248), .O(gate245inter7));
  inv1  gate1157(.a(G736), .O(gate245inter8));
  nand2 gate1158(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate1159(.a(s_87), .b(gate245inter3), .O(gate245inter10));
  nor2  gate1160(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate1161(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate1162(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate1289(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate1290(.a(gate249inter0), .b(s_106), .O(gate249inter1));
  and2  gate1291(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate1292(.a(s_106), .O(gate249inter3));
  inv1  gate1293(.a(s_107), .O(gate249inter4));
  nand2 gate1294(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate1295(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate1296(.a(G254), .O(gate249inter7));
  inv1  gate1297(.a(G742), .O(gate249inter8));
  nand2 gate1298(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate1299(.a(s_107), .b(gate249inter3), .O(gate249inter10));
  nor2  gate1300(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate1301(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate1302(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );

  xor2  gate1345(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate1346(.a(gate251inter0), .b(s_114), .O(gate251inter1));
  and2  gate1347(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate1348(.a(s_114), .O(gate251inter3));
  inv1  gate1349(.a(s_115), .O(gate251inter4));
  nand2 gate1350(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate1351(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate1352(.a(G257), .O(gate251inter7));
  inv1  gate1353(.a(G745), .O(gate251inter8));
  nand2 gate1354(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate1355(.a(s_115), .b(gate251inter3), .O(gate251inter10));
  nor2  gate1356(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate1357(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate1358(.a(gate251inter12), .b(gate251inter1), .O(G764));
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate1779(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate1780(.a(gate253inter0), .b(s_176), .O(gate253inter1));
  and2  gate1781(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate1782(.a(s_176), .O(gate253inter3));
  inv1  gate1783(.a(s_177), .O(gate253inter4));
  nand2 gate1784(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate1785(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate1786(.a(G260), .O(gate253inter7));
  inv1  gate1787(.a(G748), .O(gate253inter8));
  nand2 gate1788(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate1789(.a(s_177), .b(gate253inter3), .O(gate253inter10));
  nor2  gate1790(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate1791(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate1792(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );

  xor2  gate897(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate898(.a(gate259inter0), .b(s_50), .O(gate259inter1));
  and2  gate899(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate900(.a(s_50), .O(gate259inter3));
  inv1  gate901(.a(s_51), .O(gate259inter4));
  nand2 gate902(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate903(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate904(.a(G758), .O(gate259inter7));
  inv1  gate905(.a(G759), .O(gate259inter8));
  nand2 gate906(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate907(.a(s_51), .b(gate259inter3), .O(gate259inter10));
  nor2  gate908(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate909(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate910(.a(gate259inter12), .b(gate259inter1), .O(G776));

  xor2  gate827(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate828(.a(gate260inter0), .b(s_40), .O(gate260inter1));
  and2  gate829(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate830(.a(s_40), .O(gate260inter3));
  inv1  gate831(.a(s_41), .O(gate260inter4));
  nand2 gate832(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate833(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate834(.a(G760), .O(gate260inter7));
  inv1  gate835(.a(G761), .O(gate260inter8));
  nand2 gate836(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate837(.a(s_41), .b(gate260inter3), .O(gate260inter10));
  nor2  gate838(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate839(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate840(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );

  xor2  gate911(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate912(.a(gate264inter0), .b(s_52), .O(gate264inter1));
  and2  gate913(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate914(.a(s_52), .O(gate264inter3));
  inv1  gate915(.a(s_53), .O(gate264inter4));
  nand2 gate916(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate917(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate918(.a(G768), .O(gate264inter7));
  inv1  gate919(.a(G769), .O(gate264inter8));
  nand2 gate920(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate921(.a(s_53), .b(gate264inter3), .O(gate264inter10));
  nor2  gate922(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate923(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate924(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate1065(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate1066(.a(gate267inter0), .b(s_74), .O(gate267inter1));
  and2  gate1067(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate1068(.a(s_74), .O(gate267inter3));
  inv1  gate1069(.a(s_75), .O(gate267inter4));
  nand2 gate1070(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate1071(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate1072(.a(G648), .O(gate267inter7));
  inv1  gate1073(.a(G776), .O(gate267inter8));
  nand2 gate1074(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate1075(.a(s_75), .b(gate267inter3), .O(gate267inter10));
  nor2  gate1076(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate1077(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate1078(.a(gate267inter12), .b(gate267inter1), .O(G800));

  xor2  gate1163(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate1164(.a(gate268inter0), .b(s_88), .O(gate268inter1));
  and2  gate1165(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate1166(.a(s_88), .O(gate268inter3));
  inv1  gate1167(.a(s_89), .O(gate268inter4));
  nand2 gate1168(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1169(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1170(.a(G651), .O(gate268inter7));
  inv1  gate1171(.a(G779), .O(gate268inter8));
  nand2 gate1172(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1173(.a(s_89), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1174(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1175(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1176(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate659(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate660(.a(gate271inter0), .b(s_16), .O(gate271inter1));
  and2  gate661(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate662(.a(s_16), .O(gate271inter3));
  inv1  gate663(.a(s_17), .O(gate271inter4));
  nand2 gate664(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate665(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate666(.a(G660), .O(gate271inter7));
  inv1  gate667(.a(G788), .O(gate271inter8));
  nand2 gate668(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate669(.a(s_17), .b(gate271inter3), .O(gate271inter10));
  nor2  gate670(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate671(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate672(.a(gate271inter12), .b(gate271inter1), .O(G812));

  xor2  gate575(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate576(.a(gate272inter0), .b(s_4), .O(gate272inter1));
  and2  gate577(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate578(.a(s_4), .O(gate272inter3));
  inv1  gate579(.a(s_5), .O(gate272inter4));
  nand2 gate580(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate581(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate582(.a(G663), .O(gate272inter7));
  inv1  gate583(.a(G791), .O(gate272inter8));
  nand2 gate584(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate585(.a(s_5), .b(gate272inter3), .O(gate272inter10));
  nor2  gate586(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate587(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate588(.a(gate272inter12), .b(gate272inter1), .O(G815));

  xor2  gate1051(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate1052(.a(gate273inter0), .b(s_72), .O(gate273inter1));
  and2  gate1053(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate1054(.a(s_72), .O(gate273inter3));
  inv1  gate1055(.a(s_73), .O(gate273inter4));
  nand2 gate1056(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate1057(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate1058(.a(G642), .O(gate273inter7));
  inv1  gate1059(.a(G794), .O(gate273inter8));
  nand2 gate1060(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate1061(.a(s_73), .b(gate273inter3), .O(gate273inter10));
  nor2  gate1062(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate1063(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate1064(.a(gate273inter12), .b(gate273inter1), .O(G818));
nand2 gate274( .a(G770), .b(G794), .O(G819) );

  xor2  gate701(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate702(.a(gate275inter0), .b(s_22), .O(gate275inter1));
  and2  gate703(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate704(.a(s_22), .O(gate275inter3));
  inv1  gate705(.a(s_23), .O(gate275inter4));
  nand2 gate706(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate707(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate708(.a(G645), .O(gate275inter7));
  inv1  gate709(.a(G797), .O(gate275inter8));
  nand2 gate710(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate711(.a(s_23), .b(gate275inter3), .O(gate275inter10));
  nor2  gate712(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate713(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate714(.a(gate275inter12), .b(gate275inter1), .O(G820));
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate1191(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate1192(.a(gate280inter0), .b(s_92), .O(gate280inter1));
  and2  gate1193(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate1194(.a(s_92), .O(gate280inter3));
  inv1  gate1195(.a(s_93), .O(gate280inter4));
  nand2 gate1196(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate1197(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate1198(.a(G779), .O(gate280inter7));
  inv1  gate1199(.a(G803), .O(gate280inter8));
  nand2 gate1200(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate1201(.a(s_93), .b(gate280inter3), .O(gate280inter10));
  nor2  gate1202(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate1203(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate1204(.a(gate280inter12), .b(gate280inter1), .O(G825));
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );

  xor2  gate1527(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate1528(.a(gate284inter0), .b(s_140), .O(gate284inter1));
  and2  gate1529(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate1530(.a(s_140), .O(gate284inter3));
  inv1  gate1531(.a(s_141), .O(gate284inter4));
  nand2 gate1532(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate1533(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate1534(.a(G785), .O(gate284inter7));
  inv1  gate1535(.a(G809), .O(gate284inter8));
  nand2 gate1536(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate1537(.a(s_141), .b(gate284inter3), .O(gate284inter10));
  nor2  gate1538(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate1539(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate1540(.a(gate284inter12), .b(gate284inter1), .O(G829));
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate645(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate646(.a(gate288inter0), .b(s_14), .O(gate288inter1));
  and2  gate647(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate648(.a(s_14), .O(gate288inter3));
  inv1  gate649(.a(s_15), .O(gate288inter4));
  nand2 gate650(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate651(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate652(.a(G791), .O(gate288inter7));
  inv1  gate653(.a(G815), .O(gate288inter8));
  nand2 gate654(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate655(.a(s_15), .b(gate288inter3), .O(gate288inter10));
  nor2  gate656(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate657(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate658(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate729(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate730(.a(gate290inter0), .b(s_26), .O(gate290inter1));
  and2  gate731(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate732(.a(s_26), .O(gate290inter3));
  inv1  gate733(.a(s_27), .O(gate290inter4));
  nand2 gate734(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate735(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate736(.a(G820), .O(gate290inter7));
  inv1  gate737(.a(G821), .O(gate290inter8));
  nand2 gate738(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate739(.a(s_27), .b(gate290inter3), .O(gate290inter10));
  nor2  gate740(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate741(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate742(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate617(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate618(.a(gate292inter0), .b(s_10), .O(gate292inter1));
  and2  gate619(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate620(.a(s_10), .O(gate292inter3));
  inv1  gate621(.a(s_11), .O(gate292inter4));
  nand2 gate622(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate623(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate624(.a(G824), .O(gate292inter7));
  inv1  gate625(.a(G825), .O(gate292inter8));
  nand2 gate626(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate627(.a(s_11), .b(gate292inter3), .O(gate292inter10));
  nor2  gate628(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate629(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate630(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate1443(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate1444(.a(gate295inter0), .b(s_128), .O(gate295inter1));
  and2  gate1445(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate1446(.a(s_128), .O(gate295inter3));
  inv1  gate1447(.a(s_129), .O(gate295inter4));
  nand2 gate1448(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate1449(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate1450(.a(G830), .O(gate295inter7));
  inv1  gate1451(.a(G831), .O(gate295inter8));
  nand2 gate1452(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate1453(.a(s_129), .b(gate295inter3), .O(gate295inter10));
  nor2  gate1454(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate1455(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate1456(.a(gate295inter12), .b(gate295inter1), .O(G912));

  xor2  gate1513(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate1514(.a(gate296inter0), .b(s_138), .O(gate296inter1));
  and2  gate1515(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate1516(.a(s_138), .O(gate296inter3));
  inv1  gate1517(.a(s_139), .O(gate296inter4));
  nand2 gate1518(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate1519(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate1520(.a(G826), .O(gate296inter7));
  inv1  gate1521(.a(G827), .O(gate296inter8));
  nand2 gate1522(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate1523(.a(s_139), .b(gate296inter3), .O(gate296inter10));
  nor2  gate1524(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate1525(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate1526(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate687(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate688(.a(gate395inter0), .b(s_20), .O(gate395inter1));
  and2  gate689(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate690(.a(s_20), .O(gate395inter3));
  inv1  gate691(.a(s_21), .O(gate395inter4));
  nand2 gate692(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate693(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate694(.a(G9), .O(gate395inter7));
  inv1  gate695(.a(G1060), .O(gate395inter8));
  nand2 gate696(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate697(.a(s_21), .b(gate395inter3), .O(gate395inter10));
  nor2  gate698(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate699(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate700(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate1415(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate1416(.a(gate400inter0), .b(s_124), .O(gate400inter1));
  and2  gate1417(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate1418(.a(s_124), .O(gate400inter3));
  inv1  gate1419(.a(s_125), .O(gate400inter4));
  nand2 gate1420(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate1421(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate1422(.a(G14), .O(gate400inter7));
  inv1  gate1423(.a(G1075), .O(gate400inter8));
  nand2 gate1424(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate1425(.a(s_125), .b(gate400inter3), .O(gate400inter10));
  nor2  gate1426(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate1427(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate1428(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate1793(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate1794(.a(gate403inter0), .b(s_178), .O(gate403inter1));
  and2  gate1795(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate1796(.a(s_178), .O(gate403inter3));
  inv1  gate1797(.a(s_179), .O(gate403inter4));
  nand2 gate1798(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate1799(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate1800(.a(G17), .O(gate403inter7));
  inv1  gate1801(.a(G1084), .O(gate403inter8));
  nand2 gate1802(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate1803(.a(s_179), .b(gate403inter3), .O(gate403inter10));
  nor2  gate1804(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate1805(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate1806(.a(gate403inter12), .b(gate403inter1), .O(G1180));
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate1247(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate1248(.a(gate407inter0), .b(s_100), .O(gate407inter1));
  and2  gate1249(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate1250(.a(s_100), .O(gate407inter3));
  inv1  gate1251(.a(s_101), .O(gate407inter4));
  nand2 gate1252(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate1253(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate1254(.a(G21), .O(gate407inter7));
  inv1  gate1255(.a(G1096), .O(gate407inter8));
  nand2 gate1256(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate1257(.a(s_101), .b(gate407inter3), .O(gate407inter10));
  nor2  gate1258(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate1259(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate1260(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate1667(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate1668(.a(gate411inter0), .b(s_160), .O(gate411inter1));
  and2  gate1669(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate1670(.a(s_160), .O(gate411inter3));
  inv1  gate1671(.a(s_161), .O(gate411inter4));
  nand2 gate1672(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate1673(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate1674(.a(G25), .O(gate411inter7));
  inv1  gate1675(.a(G1108), .O(gate411inter8));
  nand2 gate1676(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate1677(.a(s_161), .b(gate411inter3), .O(gate411inter10));
  nor2  gate1678(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate1679(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate1680(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate1751(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1752(.a(gate420inter0), .b(s_172), .O(gate420inter1));
  and2  gate1753(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1754(.a(s_172), .O(gate420inter3));
  inv1  gate1755(.a(s_173), .O(gate420inter4));
  nand2 gate1756(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1757(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1758(.a(G1036), .O(gate420inter7));
  inv1  gate1759(.a(G1132), .O(gate420inter8));
  nand2 gate1760(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1761(.a(s_173), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1762(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1763(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1764(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );

  xor2  gate883(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate884(.a(gate429inter0), .b(s_48), .O(gate429inter1));
  and2  gate885(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate886(.a(s_48), .O(gate429inter3));
  inv1  gate887(.a(s_49), .O(gate429inter4));
  nand2 gate888(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate889(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate890(.a(G6), .O(gate429inter7));
  inv1  gate891(.a(G1147), .O(gate429inter8));
  nand2 gate892(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate893(.a(s_49), .b(gate429inter3), .O(gate429inter10));
  nor2  gate894(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate895(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate896(.a(gate429inter12), .b(gate429inter1), .O(G1238));

  xor2  gate995(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate996(.a(gate430inter0), .b(s_64), .O(gate430inter1));
  and2  gate997(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate998(.a(s_64), .O(gate430inter3));
  inv1  gate999(.a(s_65), .O(gate430inter4));
  nand2 gate1000(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate1001(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate1002(.a(G1051), .O(gate430inter7));
  inv1  gate1003(.a(G1147), .O(gate430inter8));
  nand2 gate1004(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate1005(.a(s_65), .b(gate430inter3), .O(gate430inter10));
  nor2  gate1006(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate1007(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate1008(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );

  xor2  gate757(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate758(.a(gate436inter0), .b(s_30), .O(gate436inter1));
  and2  gate759(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate760(.a(s_30), .O(gate436inter3));
  inv1  gate761(.a(s_31), .O(gate436inter4));
  nand2 gate762(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate763(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate764(.a(G1060), .O(gate436inter7));
  inv1  gate765(.a(G1156), .O(gate436inter8));
  nand2 gate766(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate767(.a(s_31), .b(gate436inter3), .O(gate436inter10));
  nor2  gate768(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate769(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate770(.a(gate436inter12), .b(gate436inter1), .O(G1245));
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate1499(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate1500(.a(gate443inter0), .b(s_136), .O(gate443inter1));
  and2  gate1501(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate1502(.a(s_136), .O(gate443inter3));
  inv1  gate1503(.a(s_137), .O(gate443inter4));
  nand2 gate1504(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate1505(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate1506(.a(G13), .O(gate443inter7));
  inv1  gate1507(.a(G1168), .O(gate443inter8));
  nand2 gate1508(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate1509(.a(s_137), .b(gate443inter3), .O(gate443inter10));
  nor2  gate1510(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate1511(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate1512(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );

  xor2  gate1639(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate1640(.a(gate450inter0), .b(s_156), .O(gate450inter1));
  and2  gate1641(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate1642(.a(s_156), .O(gate450inter3));
  inv1  gate1643(.a(s_157), .O(gate450inter4));
  nand2 gate1644(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate1645(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate1646(.a(G1081), .O(gate450inter7));
  inv1  gate1647(.a(G1177), .O(gate450inter8));
  nand2 gate1648(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate1649(.a(s_157), .b(gate450inter3), .O(gate450inter10));
  nor2  gate1650(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate1651(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate1652(.a(gate450inter12), .b(gate450inter1), .O(G1259));
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );

  xor2  gate715(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate716(.a(gate452inter0), .b(s_24), .O(gate452inter1));
  and2  gate717(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate718(.a(s_24), .O(gate452inter3));
  inv1  gate719(.a(s_25), .O(gate452inter4));
  nand2 gate720(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate721(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate722(.a(G1084), .O(gate452inter7));
  inv1  gate723(.a(G1180), .O(gate452inter8));
  nand2 gate724(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate725(.a(s_25), .b(gate452inter3), .O(gate452inter10));
  nor2  gate726(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate727(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate728(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );

  xor2  gate1723(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate1724(.a(gate454inter0), .b(s_168), .O(gate454inter1));
  and2  gate1725(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate1726(.a(s_168), .O(gate454inter3));
  inv1  gate1727(.a(s_169), .O(gate454inter4));
  nand2 gate1728(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate1729(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate1730(.a(G1087), .O(gate454inter7));
  inv1  gate1731(.a(G1183), .O(gate454inter8));
  nand2 gate1732(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate1733(.a(s_169), .b(gate454inter3), .O(gate454inter10));
  nor2  gate1734(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate1735(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate1736(.a(gate454inter12), .b(gate454inter1), .O(G1263));
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate1093(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate1094(.a(gate465inter0), .b(s_78), .O(gate465inter1));
  and2  gate1095(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate1096(.a(s_78), .O(gate465inter3));
  inv1  gate1097(.a(s_79), .O(gate465inter4));
  nand2 gate1098(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate1099(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate1100(.a(G24), .O(gate465inter7));
  inv1  gate1101(.a(G1201), .O(gate465inter8));
  nand2 gate1102(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate1103(.a(s_79), .b(gate465inter3), .O(gate465inter10));
  nor2  gate1104(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate1105(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate1106(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate1121(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate1122(.a(gate467inter0), .b(s_82), .O(gate467inter1));
  and2  gate1123(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate1124(.a(s_82), .O(gate467inter3));
  inv1  gate1125(.a(s_83), .O(gate467inter4));
  nand2 gate1126(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate1127(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate1128(.a(G25), .O(gate467inter7));
  inv1  gate1129(.a(G1204), .O(gate467inter8));
  nand2 gate1130(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate1131(.a(s_83), .b(gate467inter3), .O(gate467inter10));
  nor2  gate1132(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate1133(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate1134(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );

  xor2  gate1471(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate1472(.a(gate469inter0), .b(s_132), .O(gate469inter1));
  and2  gate1473(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate1474(.a(s_132), .O(gate469inter3));
  inv1  gate1475(.a(s_133), .O(gate469inter4));
  nand2 gate1476(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate1477(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate1478(.a(G26), .O(gate469inter7));
  inv1  gate1479(.a(G1207), .O(gate469inter8));
  nand2 gate1480(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate1481(.a(s_133), .b(gate469inter3), .O(gate469inter10));
  nor2  gate1482(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate1483(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate1484(.a(gate469inter12), .b(gate469inter1), .O(G1278));
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );

  xor2  gate1625(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate1626(.a(gate473inter0), .b(s_154), .O(gate473inter1));
  and2  gate1627(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate1628(.a(s_154), .O(gate473inter3));
  inv1  gate1629(.a(s_155), .O(gate473inter4));
  nand2 gate1630(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate1631(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate1632(.a(G28), .O(gate473inter7));
  inv1  gate1633(.a(G1213), .O(gate473inter8));
  nand2 gate1634(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate1635(.a(s_155), .b(gate473inter3), .O(gate473inter10));
  nor2  gate1636(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate1637(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate1638(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate1303(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate1304(.a(gate475inter0), .b(s_108), .O(gate475inter1));
  and2  gate1305(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate1306(.a(s_108), .O(gate475inter3));
  inv1  gate1307(.a(s_109), .O(gate475inter4));
  nand2 gate1308(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate1309(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate1310(.a(G29), .O(gate475inter7));
  inv1  gate1311(.a(G1216), .O(gate475inter8));
  nand2 gate1312(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate1313(.a(s_109), .b(gate475inter3), .O(gate475inter10));
  nor2  gate1314(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate1315(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate1316(.a(gate475inter12), .b(gate475inter1), .O(G1284));
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate953(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate954(.a(gate481inter0), .b(s_58), .O(gate481inter1));
  and2  gate955(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate956(.a(s_58), .O(gate481inter3));
  inv1  gate957(.a(s_59), .O(gate481inter4));
  nand2 gate958(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate959(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate960(.a(G32), .O(gate481inter7));
  inv1  gate961(.a(G1225), .O(gate481inter8));
  nand2 gate962(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate963(.a(s_59), .b(gate481inter3), .O(gate481inter10));
  nor2  gate964(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate965(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate966(.a(gate481inter12), .b(gate481inter1), .O(G1290));
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );

  xor2  gate1219(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate1220(.a(gate483inter0), .b(s_96), .O(gate483inter1));
  and2  gate1221(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate1222(.a(s_96), .O(gate483inter3));
  inv1  gate1223(.a(s_97), .O(gate483inter4));
  nand2 gate1224(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate1225(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate1226(.a(G1228), .O(gate483inter7));
  inv1  gate1227(.a(G1229), .O(gate483inter8));
  nand2 gate1228(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate1229(.a(s_97), .b(gate483inter3), .O(gate483inter10));
  nor2  gate1230(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate1231(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate1232(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate1681(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate1682(.a(gate487inter0), .b(s_162), .O(gate487inter1));
  and2  gate1683(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate1684(.a(s_162), .O(gate487inter3));
  inv1  gate1685(.a(s_163), .O(gate487inter4));
  nand2 gate1686(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate1687(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate1688(.a(G1236), .O(gate487inter7));
  inv1  gate1689(.a(G1237), .O(gate487inter8));
  nand2 gate1690(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate1691(.a(s_163), .b(gate487inter3), .O(gate487inter10));
  nor2  gate1692(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate1693(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate1694(.a(gate487inter12), .b(gate487inter1), .O(G1296));

  xor2  gate1457(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate1458(.a(gate488inter0), .b(s_130), .O(gate488inter1));
  and2  gate1459(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate1460(.a(s_130), .O(gate488inter3));
  inv1  gate1461(.a(s_131), .O(gate488inter4));
  nand2 gate1462(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate1463(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate1464(.a(G1238), .O(gate488inter7));
  inv1  gate1465(.a(G1239), .O(gate488inter8));
  nand2 gate1466(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate1467(.a(s_131), .b(gate488inter3), .O(gate488inter10));
  nor2  gate1468(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate1469(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate1470(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate1233(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate1234(.a(gate490inter0), .b(s_98), .O(gate490inter1));
  and2  gate1235(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate1236(.a(s_98), .O(gate490inter3));
  inv1  gate1237(.a(s_99), .O(gate490inter4));
  nand2 gate1238(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate1239(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate1240(.a(G1242), .O(gate490inter7));
  inv1  gate1241(.a(G1243), .O(gate490inter8));
  nand2 gate1242(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate1243(.a(s_99), .b(gate490inter3), .O(gate490inter10));
  nor2  gate1244(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate1245(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate1246(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate771(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate772(.a(gate504inter0), .b(s_32), .O(gate504inter1));
  and2  gate773(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate774(.a(s_32), .O(gate504inter3));
  inv1  gate775(.a(s_33), .O(gate504inter4));
  nand2 gate776(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate777(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate778(.a(G1270), .O(gate504inter7));
  inv1  gate779(.a(G1271), .O(gate504inter8));
  nand2 gate780(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate781(.a(s_33), .b(gate504inter3), .O(gate504inter10));
  nor2  gate782(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate783(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate784(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate1541(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate1542(.a(gate510inter0), .b(s_142), .O(gate510inter1));
  and2  gate1543(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate1544(.a(s_142), .O(gate510inter3));
  inv1  gate1545(.a(s_143), .O(gate510inter4));
  nand2 gate1546(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate1547(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate1548(.a(G1282), .O(gate510inter7));
  inv1  gate1549(.a(G1283), .O(gate510inter8));
  nand2 gate1550(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate1551(.a(s_143), .b(gate510inter3), .O(gate510inter10));
  nor2  gate1552(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate1553(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate1554(.a(gate510inter12), .b(gate510inter1), .O(G1319));

  xor2  gate589(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate590(.a(gate511inter0), .b(s_6), .O(gate511inter1));
  and2  gate591(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate592(.a(s_6), .O(gate511inter3));
  inv1  gate593(.a(s_7), .O(gate511inter4));
  nand2 gate594(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate595(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate596(.a(G1284), .O(gate511inter7));
  inv1  gate597(.a(G1285), .O(gate511inter8));
  nand2 gate598(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate599(.a(s_7), .b(gate511inter3), .O(gate511inter10));
  nor2  gate600(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate601(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate602(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate1331(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate1332(.a(gate514inter0), .b(s_112), .O(gate514inter1));
  and2  gate1333(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate1334(.a(s_112), .O(gate514inter3));
  inv1  gate1335(.a(s_113), .O(gate514inter4));
  nand2 gate1336(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate1337(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate1338(.a(G1290), .O(gate514inter7));
  inv1  gate1339(.a(G1291), .O(gate514inter8));
  nand2 gate1340(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate1341(.a(s_113), .b(gate514inter3), .O(gate514inter10));
  nor2  gate1342(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate1343(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate1344(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule