module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate1401(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate1402(.a(gate15inter0), .b(s_122), .O(gate15inter1));
  and2  gate1403(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate1404(.a(s_122), .O(gate15inter3));
  inv1  gate1405(.a(s_123), .O(gate15inter4));
  nand2 gate1406(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate1407(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate1408(.a(G13), .O(gate15inter7));
  inv1  gate1409(.a(G14), .O(gate15inter8));
  nand2 gate1410(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate1411(.a(s_123), .b(gate15inter3), .O(gate15inter10));
  nor2  gate1412(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate1413(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate1414(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate925(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate926(.a(gate27inter0), .b(s_54), .O(gate27inter1));
  and2  gate927(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate928(.a(s_54), .O(gate27inter3));
  inv1  gate929(.a(s_55), .O(gate27inter4));
  nand2 gate930(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate931(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate932(.a(G2), .O(gate27inter7));
  inv1  gate933(.a(G6), .O(gate27inter8));
  nand2 gate934(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate935(.a(s_55), .b(gate27inter3), .O(gate27inter10));
  nor2  gate936(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate937(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate938(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );

  xor2  gate1079(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate1080(.a(gate30inter0), .b(s_76), .O(gate30inter1));
  and2  gate1081(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate1082(.a(s_76), .O(gate30inter3));
  inv1  gate1083(.a(s_77), .O(gate30inter4));
  nand2 gate1084(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate1085(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate1086(.a(G11), .O(gate30inter7));
  inv1  gate1087(.a(G15), .O(gate30inter8));
  nand2 gate1088(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate1089(.a(s_77), .b(gate30inter3), .O(gate30inter10));
  nor2  gate1090(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate1091(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate1092(.a(gate30inter12), .b(gate30inter1), .O(G329));
nand2 gate31( .a(G4), .b(G8), .O(G332) );

  xor2  gate1457(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate1458(.a(gate32inter0), .b(s_130), .O(gate32inter1));
  and2  gate1459(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate1460(.a(s_130), .O(gate32inter3));
  inv1  gate1461(.a(s_131), .O(gate32inter4));
  nand2 gate1462(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate1463(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate1464(.a(G12), .O(gate32inter7));
  inv1  gate1465(.a(G16), .O(gate32inter8));
  nand2 gate1466(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate1467(.a(s_131), .b(gate32inter3), .O(gate32inter10));
  nor2  gate1468(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate1469(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate1470(.a(gate32inter12), .b(gate32inter1), .O(G335));
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );

  xor2  gate799(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate800(.a(gate35inter0), .b(s_36), .O(gate35inter1));
  and2  gate801(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate802(.a(s_36), .O(gate35inter3));
  inv1  gate803(.a(s_37), .O(gate35inter4));
  nand2 gate804(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate805(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate806(.a(G18), .O(gate35inter7));
  inv1  gate807(.a(G22), .O(gate35inter8));
  nand2 gate808(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate809(.a(s_37), .b(gate35inter3), .O(gate35inter10));
  nor2  gate810(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate811(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate812(.a(gate35inter12), .b(gate35inter1), .O(G344));
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );

  xor2  gate911(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate912(.a(gate48inter0), .b(s_52), .O(gate48inter1));
  and2  gate913(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate914(.a(s_52), .O(gate48inter3));
  inv1  gate915(.a(s_53), .O(gate48inter4));
  nand2 gate916(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate917(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate918(.a(G8), .O(gate48inter7));
  inv1  gate919(.a(G275), .O(gate48inter8));
  nand2 gate920(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate921(.a(s_53), .b(gate48inter3), .O(gate48inter10));
  nor2  gate922(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate923(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate924(.a(gate48inter12), .b(gate48inter1), .O(G369));
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate1163(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate1164(.a(gate51inter0), .b(s_88), .O(gate51inter1));
  and2  gate1165(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate1166(.a(s_88), .O(gate51inter3));
  inv1  gate1167(.a(s_89), .O(gate51inter4));
  nand2 gate1168(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate1169(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate1170(.a(G11), .O(gate51inter7));
  inv1  gate1171(.a(G281), .O(gate51inter8));
  nand2 gate1172(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate1173(.a(s_89), .b(gate51inter3), .O(gate51inter10));
  nor2  gate1174(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate1175(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate1176(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );

  xor2  gate771(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate772(.a(gate56inter0), .b(s_32), .O(gate56inter1));
  and2  gate773(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate774(.a(s_32), .O(gate56inter3));
  inv1  gate775(.a(s_33), .O(gate56inter4));
  nand2 gate776(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate777(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate778(.a(G16), .O(gate56inter7));
  inv1  gate779(.a(G287), .O(gate56inter8));
  nand2 gate780(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate781(.a(s_33), .b(gate56inter3), .O(gate56inter10));
  nor2  gate782(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate783(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate784(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate701(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate702(.a(gate60inter0), .b(s_22), .O(gate60inter1));
  and2  gate703(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate704(.a(s_22), .O(gate60inter3));
  inv1  gate705(.a(s_23), .O(gate60inter4));
  nand2 gate706(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate707(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate708(.a(G20), .O(gate60inter7));
  inv1  gate709(.a(G293), .O(gate60inter8));
  nand2 gate710(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate711(.a(s_23), .b(gate60inter3), .O(gate60inter10));
  nor2  gate712(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate713(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate714(.a(gate60inter12), .b(gate60inter1), .O(G381));

  xor2  gate855(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate856(.a(gate61inter0), .b(s_44), .O(gate61inter1));
  and2  gate857(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate858(.a(s_44), .O(gate61inter3));
  inv1  gate859(.a(s_45), .O(gate61inter4));
  nand2 gate860(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate861(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate862(.a(G21), .O(gate61inter7));
  inv1  gate863(.a(G296), .O(gate61inter8));
  nand2 gate864(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate865(.a(s_45), .b(gate61inter3), .O(gate61inter10));
  nor2  gate866(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate867(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate868(.a(gate61inter12), .b(gate61inter1), .O(G382));
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate1331(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate1332(.a(gate66inter0), .b(s_112), .O(gate66inter1));
  and2  gate1333(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate1334(.a(s_112), .O(gate66inter3));
  inv1  gate1335(.a(s_113), .O(gate66inter4));
  nand2 gate1336(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate1337(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate1338(.a(G26), .O(gate66inter7));
  inv1  gate1339(.a(G302), .O(gate66inter8));
  nand2 gate1340(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate1341(.a(s_113), .b(gate66inter3), .O(gate66inter10));
  nor2  gate1342(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate1343(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate1344(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate953(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate954(.a(gate69inter0), .b(s_58), .O(gate69inter1));
  and2  gate955(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate956(.a(s_58), .O(gate69inter3));
  inv1  gate957(.a(s_59), .O(gate69inter4));
  nand2 gate958(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate959(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate960(.a(G29), .O(gate69inter7));
  inv1  gate961(.a(G308), .O(gate69inter8));
  nand2 gate962(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate963(.a(s_59), .b(gate69inter3), .O(gate69inter10));
  nor2  gate964(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate965(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate966(.a(gate69inter12), .b(gate69inter1), .O(G390));
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate757(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate758(.a(gate85inter0), .b(s_30), .O(gate85inter1));
  and2  gate759(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate760(.a(s_30), .O(gate85inter3));
  inv1  gate761(.a(s_31), .O(gate85inter4));
  nand2 gate762(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate763(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate764(.a(G4), .O(gate85inter7));
  inv1  gate765(.a(G332), .O(gate85inter8));
  nand2 gate766(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate767(.a(s_31), .b(gate85inter3), .O(gate85inter10));
  nor2  gate768(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate769(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate770(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );

  xor2  gate673(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate674(.a(gate87inter0), .b(s_18), .O(gate87inter1));
  and2  gate675(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate676(.a(s_18), .O(gate87inter3));
  inv1  gate677(.a(s_19), .O(gate87inter4));
  nand2 gate678(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate679(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate680(.a(G12), .O(gate87inter7));
  inv1  gate681(.a(G335), .O(gate87inter8));
  nand2 gate682(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate683(.a(s_19), .b(gate87inter3), .O(gate87inter10));
  nor2  gate684(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate685(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate686(.a(gate87inter12), .b(gate87inter1), .O(G408));

  xor2  gate575(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate576(.a(gate88inter0), .b(s_4), .O(gate88inter1));
  and2  gate577(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate578(.a(s_4), .O(gate88inter3));
  inv1  gate579(.a(s_5), .O(gate88inter4));
  nand2 gate580(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate581(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate582(.a(G16), .O(gate88inter7));
  inv1  gate583(.a(G335), .O(gate88inter8));
  nand2 gate584(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate585(.a(s_5), .b(gate88inter3), .O(gate88inter10));
  nor2  gate586(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate587(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate588(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate1065(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate1066(.a(gate96inter0), .b(s_74), .O(gate96inter1));
  and2  gate1067(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate1068(.a(s_74), .O(gate96inter3));
  inv1  gate1069(.a(s_75), .O(gate96inter4));
  nand2 gate1070(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate1071(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate1072(.a(G30), .O(gate96inter7));
  inv1  gate1073(.a(G347), .O(gate96inter8));
  nand2 gate1074(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate1075(.a(s_75), .b(gate96inter3), .O(gate96inter10));
  nor2  gate1076(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate1077(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate1078(.a(gate96inter12), .b(gate96inter1), .O(G417));
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate1135(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate1136(.a(gate98inter0), .b(s_84), .O(gate98inter1));
  and2  gate1137(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate1138(.a(s_84), .O(gate98inter3));
  inv1  gate1139(.a(s_85), .O(gate98inter4));
  nand2 gate1140(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1141(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1142(.a(G23), .O(gate98inter7));
  inv1  gate1143(.a(G350), .O(gate98inter8));
  nand2 gate1144(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1145(.a(s_85), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1146(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1147(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1148(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate827(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate828(.a(gate106inter0), .b(s_40), .O(gate106inter1));
  and2  gate829(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate830(.a(s_40), .O(gate106inter3));
  inv1  gate831(.a(s_41), .O(gate106inter4));
  nand2 gate832(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate833(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate834(.a(G364), .O(gate106inter7));
  inv1  gate835(.a(G365), .O(gate106inter8));
  nand2 gate836(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate837(.a(s_41), .b(gate106inter3), .O(gate106inter10));
  nor2  gate838(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate839(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate840(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate1485(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate1486(.a(gate116inter0), .b(s_134), .O(gate116inter1));
  and2  gate1487(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate1488(.a(s_134), .O(gate116inter3));
  inv1  gate1489(.a(s_135), .O(gate116inter4));
  nand2 gate1490(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate1491(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate1492(.a(G384), .O(gate116inter7));
  inv1  gate1493(.a(G385), .O(gate116inter8));
  nand2 gate1494(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate1495(.a(s_135), .b(gate116inter3), .O(gate116inter10));
  nor2  gate1496(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate1497(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate1498(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate1219(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate1220(.a(gate121inter0), .b(s_96), .O(gate121inter1));
  and2  gate1221(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate1222(.a(s_96), .O(gate121inter3));
  inv1  gate1223(.a(s_97), .O(gate121inter4));
  nand2 gate1224(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate1225(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate1226(.a(G394), .O(gate121inter7));
  inv1  gate1227(.a(G395), .O(gate121inter8));
  nand2 gate1228(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate1229(.a(s_97), .b(gate121inter3), .O(gate121inter10));
  nor2  gate1230(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate1231(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate1232(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate547(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate548(.a(gate124inter0), .b(s_0), .O(gate124inter1));
  and2  gate549(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate550(.a(s_0), .O(gate124inter3));
  inv1  gate551(.a(s_1), .O(gate124inter4));
  nand2 gate552(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate553(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate554(.a(G400), .O(gate124inter7));
  inv1  gate555(.a(G401), .O(gate124inter8));
  nand2 gate556(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate557(.a(s_1), .b(gate124inter3), .O(gate124inter10));
  nor2  gate558(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate559(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate560(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate1023(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate1024(.a(gate128inter0), .b(s_68), .O(gate128inter1));
  and2  gate1025(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate1026(.a(s_68), .O(gate128inter3));
  inv1  gate1027(.a(s_69), .O(gate128inter4));
  nand2 gate1028(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate1029(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate1030(.a(G408), .O(gate128inter7));
  inv1  gate1031(.a(G409), .O(gate128inter8));
  nand2 gate1032(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate1033(.a(s_69), .b(gate128inter3), .O(gate128inter10));
  nor2  gate1034(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate1035(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate1036(.a(gate128inter12), .b(gate128inter1), .O(G495));
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate1415(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate1416(.a(gate130inter0), .b(s_124), .O(gate130inter1));
  and2  gate1417(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate1418(.a(s_124), .O(gate130inter3));
  inv1  gate1419(.a(s_125), .O(gate130inter4));
  nand2 gate1420(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate1421(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate1422(.a(G412), .O(gate130inter7));
  inv1  gate1423(.a(G413), .O(gate130inter8));
  nand2 gate1424(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate1425(.a(s_125), .b(gate130inter3), .O(gate130inter10));
  nor2  gate1426(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate1427(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate1428(.a(gate130inter12), .b(gate130inter1), .O(G501));
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate841(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate842(.a(gate138inter0), .b(s_42), .O(gate138inter1));
  and2  gate843(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate844(.a(s_42), .O(gate138inter3));
  inv1  gate845(.a(s_43), .O(gate138inter4));
  nand2 gate846(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate847(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate848(.a(G432), .O(gate138inter7));
  inv1  gate849(.a(G435), .O(gate138inter8));
  nand2 gate850(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate851(.a(s_43), .b(gate138inter3), .O(gate138inter10));
  nor2  gate852(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate853(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate854(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate883(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate884(.a(gate143inter0), .b(s_48), .O(gate143inter1));
  and2  gate885(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate886(.a(s_48), .O(gate143inter3));
  inv1  gate887(.a(s_49), .O(gate143inter4));
  nand2 gate888(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate889(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate890(.a(G462), .O(gate143inter7));
  inv1  gate891(.a(G465), .O(gate143inter8));
  nand2 gate892(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate893(.a(s_49), .b(gate143inter3), .O(gate143inter10));
  nor2  gate894(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate895(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate896(.a(gate143inter12), .b(gate143inter1), .O(G540));
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate1499(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1500(.a(gate148inter0), .b(s_136), .O(gate148inter1));
  and2  gate1501(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1502(.a(s_136), .O(gate148inter3));
  inv1  gate1503(.a(s_137), .O(gate148inter4));
  nand2 gate1504(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1505(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1506(.a(G492), .O(gate148inter7));
  inv1  gate1507(.a(G495), .O(gate148inter8));
  nand2 gate1508(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1509(.a(s_137), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1510(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1511(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1512(.a(gate148inter12), .b(gate148inter1), .O(G555));

  xor2  gate897(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate898(.a(gate149inter0), .b(s_50), .O(gate149inter1));
  and2  gate899(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate900(.a(s_50), .O(gate149inter3));
  inv1  gate901(.a(s_51), .O(gate149inter4));
  nand2 gate902(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate903(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate904(.a(G498), .O(gate149inter7));
  inv1  gate905(.a(G501), .O(gate149inter8));
  nand2 gate906(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate907(.a(s_51), .b(gate149inter3), .O(gate149inter10));
  nor2  gate908(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate909(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate910(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate659(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate660(.a(gate164inter0), .b(s_16), .O(gate164inter1));
  and2  gate661(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate662(.a(s_16), .O(gate164inter3));
  inv1  gate663(.a(s_17), .O(gate164inter4));
  nand2 gate664(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate665(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate666(.a(G459), .O(gate164inter7));
  inv1  gate667(.a(G537), .O(gate164inter8));
  nand2 gate668(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate669(.a(s_17), .b(gate164inter3), .O(gate164inter10));
  nor2  gate670(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate671(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate672(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );

  xor2  gate1345(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate1346(.a(gate166inter0), .b(s_114), .O(gate166inter1));
  and2  gate1347(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate1348(.a(s_114), .O(gate166inter3));
  inv1  gate1349(.a(s_115), .O(gate166inter4));
  nand2 gate1350(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate1351(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate1352(.a(G465), .O(gate166inter7));
  inv1  gate1353(.a(G540), .O(gate166inter8));
  nand2 gate1354(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate1355(.a(s_115), .b(gate166inter3), .O(gate166inter10));
  nor2  gate1356(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate1357(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate1358(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate1107(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate1108(.a(gate178inter0), .b(s_80), .O(gate178inter1));
  and2  gate1109(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate1110(.a(s_80), .O(gate178inter3));
  inv1  gate1111(.a(s_81), .O(gate178inter4));
  nand2 gate1112(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate1113(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate1114(.a(G501), .O(gate178inter7));
  inv1  gate1115(.a(G558), .O(gate178inter8));
  nand2 gate1116(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate1117(.a(s_81), .b(gate178inter3), .O(gate178inter10));
  nor2  gate1118(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate1119(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate1120(.a(gate178inter12), .b(gate178inter1), .O(G595));
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate1471(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1472(.a(gate186inter0), .b(s_132), .O(gate186inter1));
  and2  gate1473(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1474(.a(s_132), .O(gate186inter3));
  inv1  gate1475(.a(s_133), .O(gate186inter4));
  nand2 gate1476(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1477(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1478(.a(G572), .O(gate186inter7));
  inv1  gate1479(.a(G573), .O(gate186inter8));
  nand2 gate1480(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1481(.a(s_133), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1482(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1483(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1484(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );

  xor2  gate869(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate870(.a(gate194inter0), .b(s_46), .O(gate194inter1));
  and2  gate871(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate872(.a(s_46), .O(gate194inter3));
  inv1  gate873(.a(s_47), .O(gate194inter4));
  nand2 gate874(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate875(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate876(.a(G588), .O(gate194inter7));
  inv1  gate877(.a(G589), .O(gate194inter8));
  nand2 gate878(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate879(.a(s_47), .b(gate194inter3), .O(gate194inter10));
  nor2  gate880(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate881(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate882(.a(gate194inter12), .b(gate194inter1), .O(G645));

  xor2  gate687(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate688(.a(gate195inter0), .b(s_20), .O(gate195inter1));
  and2  gate689(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate690(.a(s_20), .O(gate195inter3));
  inv1  gate691(.a(s_21), .O(gate195inter4));
  nand2 gate692(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate693(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate694(.a(G590), .O(gate195inter7));
  inv1  gate695(.a(G591), .O(gate195inter8));
  nand2 gate696(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate697(.a(s_21), .b(gate195inter3), .O(gate195inter10));
  nor2  gate698(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate699(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate700(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate1513(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate1514(.a(gate198inter0), .b(s_138), .O(gate198inter1));
  and2  gate1515(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate1516(.a(s_138), .O(gate198inter3));
  inv1  gate1517(.a(s_139), .O(gate198inter4));
  nand2 gate1518(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate1519(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate1520(.a(G596), .O(gate198inter7));
  inv1  gate1521(.a(G597), .O(gate198inter8));
  nand2 gate1522(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate1523(.a(s_139), .b(gate198inter3), .O(gate198inter10));
  nor2  gate1524(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate1525(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate1526(.a(gate198inter12), .b(gate198inter1), .O(G657));

  xor2  gate1149(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate1150(.a(gate199inter0), .b(s_86), .O(gate199inter1));
  and2  gate1151(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate1152(.a(s_86), .O(gate199inter3));
  inv1  gate1153(.a(s_87), .O(gate199inter4));
  nand2 gate1154(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate1155(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate1156(.a(G598), .O(gate199inter7));
  inv1  gate1157(.a(G599), .O(gate199inter8));
  nand2 gate1158(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate1159(.a(s_87), .b(gate199inter3), .O(gate199inter10));
  nor2  gate1160(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate1161(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate1162(.a(gate199inter12), .b(gate199inter1), .O(G660));

  xor2  gate715(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate716(.a(gate200inter0), .b(s_24), .O(gate200inter1));
  and2  gate717(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate718(.a(s_24), .O(gate200inter3));
  inv1  gate719(.a(s_25), .O(gate200inter4));
  nand2 gate720(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate721(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate722(.a(G600), .O(gate200inter7));
  inv1  gate723(.a(G601), .O(gate200inter8));
  nand2 gate724(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate725(.a(s_25), .b(gate200inter3), .O(gate200inter10));
  nor2  gate726(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate727(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate728(.a(gate200inter12), .b(gate200inter1), .O(G663));
nand2 gate201( .a(G602), .b(G607), .O(G666) );

  xor2  gate1009(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate1010(.a(gate202inter0), .b(s_66), .O(gate202inter1));
  and2  gate1011(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate1012(.a(s_66), .O(gate202inter3));
  inv1  gate1013(.a(s_67), .O(gate202inter4));
  nand2 gate1014(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate1015(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate1016(.a(G612), .O(gate202inter7));
  inv1  gate1017(.a(G617), .O(gate202inter8));
  nand2 gate1018(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate1019(.a(s_67), .b(gate202inter3), .O(gate202inter10));
  nor2  gate1020(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate1021(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate1022(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate1303(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate1304(.a(gate205inter0), .b(s_108), .O(gate205inter1));
  and2  gate1305(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate1306(.a(s_108), .O(gate205inter3));
  inv1  gate1307(.a(s_109), .O(gate205inter4));
  nand2 gate1308(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate1309(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate1310(.a(G622), .O(gate205inter7));
  inv1  gate1311(.a(G627), .O(gate205inter8));
  nand2 gate1312(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate1313(.a(s_109), .b(gate205inter3), .O(gate205inter10));
  nor2  gate1314(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate1315(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate1316(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );

  xor2  gate1359(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate1360(.a(gate210inter0), .b(s_116), .O(gate210inter1));
  and2  gate1361(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate1362(.a(s_116), .O(gate210inter3));
  inv1  gate1363(.a(s_117), .O(gate210inter4));
  nand2 gate1364(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate1365(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate1366(.a(G607), .O(gate210inter7));
  inv1  gate1367(.a(G666), .O(gate210inter8));
  nand2 gate1368(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate1369(.a(s_117), .b(gate210inter3), .O(gate210inter10));
  nor2  gate1370(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate1371(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate1372(.a(gate210inter12), .b(gate210inter1), .O(G691));
nand2 gate211( .a(G612), .b(G669), .O(G692) );

  xor2  gate785(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate786(.a(gate212inter0), .b(s_34), .O(gate212inter1));
  and2  gate787(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate788(.a(s_34), .O(gate212inter3));
  inv1  gate789(.a(s_35), .O(gate212inter4));
  nand2 gate790(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate791(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate792(.a(G617), .O(gate212inter7));
  inv1  gate793(.a(G669), .O(gate212inter8));
  nand2 gate794(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate795(.a(s_35), .b(gate212inter3), .O(gate212inter10));
  nor2  gate796(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate797(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate798(.a(gate212inter12), .b(gate212inter1), .O(G693));

  xor2  gate603(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate604(.a(gate213inter0), .b(s_8), .O(gate213inter1));
  and2  gate605(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate606(.a(s_8), .O(gate213inter3));
  inv1  gate607(.a(s_9), .O(gate213inter4));
  nand2 gate608(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate609(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate610(.a(G602), .O(gate213inter7));
  inv1  gate611(.a(G672), .O(gate213inter8));
  nand2 gate612(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate613(.a(s_9), .b(gate213inter3), .O(gate213inter10));
  nor2  gate614(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate615(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate616(.a(gate213inter12), .b(gate213inter1), .O(G694));

  xor2  gate645(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate646(.a(gate214inter0), .b(s_14), .O(gate214inter1));
  and2  gate647(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate648(.a(s_14), .O(gate214inter3));
  inv1  gate649(.a(s_15), .O(gate214inter4));
  nand2 gate650(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate651(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate652(.a(G612), .O(gate214inter7));
  inv1  gate653(.a(G672), .O(gate214inter8));
  nand2 gate654(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate655(.a(s_15), .b(gate214inter3), .O(gate214inter10));
  nor2  gate656(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate657(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate658(.a(gate214inter12), .b(gate214inter1), .O(G695));

  xor2  gate1289(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate1290(.a(gate215inter0), .b(s_106), .O(gate215inter1));
  and2  gate1291(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate1292(.a(s_106), .O(gate215inter3));
  inv1  gate1293(.a(s_107), .O(gate215inter4));
  nand2 gate1294(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate1295(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate1296(.a(G607), .O(gate215inter7));
  inv1  gate1297(.a(G675), .O(gate215inter8));
  nand2 gate1298(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate1299(.a(s_107), .b(gate215inter3), .O(gate215inter10));
  nor2  gate1300(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate1301(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate1302(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate1191(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate1192(.a(gate228inter0), .b(s_92), .O(gate228inter1));
  and2  gate1193(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate1194(.a(s_92), .O(gate228inter3));
  inv1  gate1195(.a(s_93), .O(gate228inter4));
  nand2 gate1196(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate1197(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate1198(.a(G696), .O(gate228inter7));
  inv1  gate1199(.a(G697), .O(gate228inter8));
  nand2 gate1200(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate1201(.a(s_93), .b(gate228inter3), .O(gate228inter10));
  nor2  gate1202(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate1203(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate1204(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate1233(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate1234(.a(gate231inter0), .b(s_98), .O(gate231inter1));
  and2  gate1235(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate1236(.a(s_98), .O(gate231inter3));
  inv1  gate1237(.a(s_99), .O(gate231inter4));
  nand2 gate1238(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate1239(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate1240(.a(G702), .O(gate231inter7));
  inv1  gate1241(.a(G703), .O(gate231inter8));
  nand2 gate1242(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate1243(.a(s_99), .b(gate231inter3), .O(gate231inter10));
  nor2  gate1244(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate1245(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate1246(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate1527(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate1528(.a(gate234inter0), .b(s_140), .O(gate234inter1));
  and2  gate1529(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate1530(.a(s_140), .O(gate234inter3));
  inv1  gate1531(.a(s_141), .O(gate234inter4));
  nand2 gate1532(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1533(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1534(.a(G245), .O(gate234inter7));
  inv1  gate1535(.a(G721), .O(gate234inter8));
  nand2 gate1536(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1537(.a(s_141), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1538(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1539(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1540(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate1429(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate1430(.a(gate249inter0), .b(s_126), .O(gate249inter1));
  and2  gate1431(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate1432(.a(s_126), .O(gate249inter3));
  inv1  gate1433(.a(s_127), .O(gate249inter4));
  nand2 gate1434(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate1435(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate1436(.a(G254), .O(gate249inter7));
  inv1  gate1437(.a(G742), .O(gate249inter8));
  nand2 gate1438(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate1439(.a(s_127), .b(gate249inter3), .O(gate249inter10));
  nor2  gate1440(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate1441(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate1442(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate1121(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate1122(.a(gate252inter0), .b(s_82), .O(gate252inter1));
  and2  gate1123(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate1124(.a(s_82), .O(gate252inter3));
  inv1  gate1125(.a(s_83), .O(gate252inter4));
  nand2 gate1126(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate1127(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate1128(.a(G709), .O(gate252inter7));
  inv1  gate1129(.a(G745), .O(gate252inter8));
  nand2 gate1130(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate1131(.a(s_83), .b(gate252inter3), .O(gate252inter10));
  nor2  gate1132(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate1133(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate1134(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate1387(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate1388(.a(gate262inter0), .b(s_120), .O(gate262inter1));
  and2  gate1389(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate1390(.a(s_120), .O(gate262inter3));
  inv1  gate1391(.a(s_121), .O(gate262inter4));
  nand2 gate1392(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate1393(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate1394(.a(G764), .O(gate262inter7));
  inv1  gate1395(.a(G765), .O(gate262inter8));
  nand2 gate1396(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate1397(.a(s_121), .b(gate262inter3), .O(gate262inter10));
  nor2  gate1398(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate1399(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate1400(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate729(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate730(.a(gate269inter0), .b(s_26), .O(gate269inter1));
  and2  gate731(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate732(.a(s_26), .O(gate269inter3));
  inv1  gate733(.a(s_27), .O(gate269inter4));
  nand2 gate734(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate735(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate736(.a(G654), .O(gate269inter7));
  inv1  gate737(.a(G782), .O(gate269inter8));
  nand2 gate738(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate739(.a(s_27), .b(gate269inter3), .O(gate269inter10));
  nor2  gate740(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate741(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate742(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate1051(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate1052(.a(gate276inter0), .b(s_72), .O(gate276inter1));
  and2  gate1053(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate1054(.a(s_72), .O(gate276inter3));
  inv1  gate1055(.a(s_73), .O(gate276inter4));
  nand2 gate1056(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate1057(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate1058(.a(G773), .O(gate276inter7));
  inv1  gate1059(.a(G797), .O(gate276inter8));
  nand2 gate1060(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate1061(.a(s_73), .b(gate276inter3), .O(gate276inter10));
  nor2  gate1062(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate1063(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate1064(.a(gate276inter12), .b(gate276inter1), .O(G821));

  xor2  gate1177(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate1178(.a(gate277inter0), .b(s_90), .O(gate277inter1));
  and2  gate1179(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate1180(.a(s_90), .O(gate277inter3));
  inv1  gate1181(.a(s_91), .O(gate277inter4));
  nand2 gate1182(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate1183(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate1184(.a(G648), .O(gate277inter7));
  inv1  gate1185(.a(G800), .O(gate277inter8));
  nand2 gate1186(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate1187(.a(s_91), .b(gate277inter3), .O(gate277inter10));
  nor2  gate1188(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate1189(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate1190(.a(gate277inter12), .b(gate277inter1), .O(G822));
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );

  xor2  gate743(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate744(.a(gate284inter0), .b(s_28), .O(gate284inter1));
  and2  gate745(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate746(.a(s_28), .O(gate284inter3));
  inv1  gate747(.a(s_29), .O(gate284inter4));
  nand2 gate748(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate749(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate750(.a(G785), .O(gate284inter7));
  inv1  gate751(.a(G809), .O(gate284inter8));
  nand2 gate752(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate753(.a(s_29), .b(gate284inter3), .O(gate284inter10));
  nor2  gate754(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate755(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate756(.a(gate284inter12), .b(gate284inter1), .O(G829));
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate1037(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate1038(.a(gate288inter0), .b(s_70), .O(gate288inter1));
  and2  gate1039(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate1040(.a(s_70), .O(gate288inter3));
  inv1  gate1041(.a(s_71), .O(gate288inter4));
  nand2 gate1042(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate1043(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate1044(.a(G791), .O(gate288inter7));
  inv1  gate1045(.a(G815), .O(gate288inter8));
  nand2 gate1046(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate1047(.a(s_71), .b(gate288inter3), .O(gate288inter10));
  nor2  gate1048(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate1049(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate1050(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate995(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate996(.a(gate292inter0), .b(s_64), .O(gate292inter1));
  and2  gate997(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate998(.a(s_64), .O(gate292inter3));
  inv1  gate999(.a(s_65), .O(gate292inter4));
  nand2 gate1000(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate1001(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate1002(.a(G824), .O(gate292inter7));
  inv1  gate1003(.a(G825), .O(gate292inter8));
  nand2 gate1004(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate1005(.a(s_65), .b(gate292inter3), .O(gate292inter10));
  nor2  gate1006(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate1007(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate1008(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate813(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate814(.a(gate296inter0), .b(s_38), .O(gate296inter1));
  and2  gate815(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate816(.a(s_38), .O(gate296inter3));
  inv1  gate817(.a(s_39), .O(gate296inter4));
  nand2 gate818(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate819(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate820(.a(G826), .O(gate296inter7));
  inv1  gate821(.a(G827), .O(gate296inter8));
  nand2 gate822(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate823(.a(s_39), .b(gate296inter3), .O(gate296inter10));
  nor2  gate824(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate825(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate826(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );

  xor2  gate1205(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate1206(.a(gate412inter0), .b(s_94), .O(gate412inter1));
  and2  gate1207(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate1208(.a(s_94), .O(gate412inter3));
  inv1  gate1209(.a(s_95), .O(gate412inter4));
  nand2 gate1210(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate1211(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate1212(.a(G26), .O(gate412inter7));
  inv1  gate1213(.a(G1111), .O(gate412inter8));
  nand2 gate1214(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate1215(.a(s_95), .b(gate412inter3), .O(gate412inter10));
  nor2  gate1216(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate1217(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate1218(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate561(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate562(.a(gate425inter0), .b(s_2), .O(gate425inter1));
  and2  gate563(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate564(.a(s_2), .O(gate425inter3));
  inv1  gate565(.a(s_3), .O(gate425inter4));
  nand2 gate566(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate567(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate568(.a(G4), .O(gate425inter7));
  inv1  gate569(.a(G1141), .O(gate425inter8));
  nand2 gate570(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate571(.a(s_3), .b(gate425inter3), .O(gate425inter10));
  nor2  gate572(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate573(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate574(.a(gate425inter12), .b(gate425inter1), .O(G1234));
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate1275(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate1276(.a(gate428inter0), .b(s_104), .O(gate428inter1));
  and2  gate1277(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate1278(.a(s_104), .O(gate428inter3));
  inv1  gate1279(.a(s_105), .O(gate428inter4));
  nand2 gate1280(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate1281(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate1282(.a(G1048), .O(gate428inter7));
  inv1  gate1283(.a(G1144), .O(gate428inter8));
  nand2 gate1284(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate1285(.a(s_105), .b(gate428inter3), .O(gate428inter10));
  nor2  gate1286(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate1287(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate1288(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate939(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate940(.a(gate432inter0), .b(s_56), .O(gate432inter1));
  and2  gate941(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate942(.a(s_56), .O(gate432inter3));
  inv1  gate943(.a(s_57), .O(gate432inter4));
  nand2 gate944(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate945(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate946(.a(G1054), .O(gate432inter7));
  inv1  gate947(.a(G1150), .O(gate432inter8));
  nand2 gate948(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate949(.a(s_57), .b(gate432inter3), .O(gate432inter10));
  nor2  gate950(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate951(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate952(.a(gate432inter12), .b(gate432inter1), .O(G1241));

  xor2  gate631(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate632(.a(gate433inter0), .b(s_12), .O(gate433inter1));
  and2  gate633(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate634(.a(s_12), .O(gate433inter3));
  inv1  gate635(.a(s_13), .O(gate433inter4));
  nand2 gate636(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate637(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate638(.a(G8), .O(gate433inter7));
  inv1  gate639(.a(G1153), .O(gate433inter8));
  nand2 gate640(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate641(.a(s_13), .b(gate433inter3), .O(gate433inter10));
  nor2  gate642(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate643(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate644(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate1317(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate1318(.a(gate438inter0), .b(s_110), .O(gate438inter1));
  and2  gate1319(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate1320(.a(s_110), .O(gate438inter3));
  inv1  gate1321(.a(s_111), .O(gate438inter4));
  nand2 gate1322(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate1323(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate1324(.a(G1063), .O(gate438inter7));
  inv1  gate1325(.a(G1159), .O(gate438inter8));
  nand2 gate1326(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate1327(.a(s_111), .b(gate438inter3), .O(gate438inter10));
  nor2  gate1328(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate1329(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate1330(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate1443(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate1444(.a(gate445inter0), .b(s_128), .O(gate445inter1));
  and2  gate1445(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate1446(.a(s_128), .O(gate445inter3));
  inv1  gate1447(.a(s_129), .O(gate445inter4));
  nand2 gate1448(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate1449(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate1450(.a(G14), .O(gate445inter7));
  inv1  gate1451(.a(G1171), .O(gate445inter8));
  nand2 gate1452(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate1453(.a(s_129), .b(gate445inter3), .O(gate445inter10));
  nor2  gate1454(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate1455(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate1456(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );

  xor2  gate1261(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate1262(.a(gate451inter0), .b(s_102), .O(gate451inter1));
  and2  gate1263(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate1264(.a(s_102), .O(gate451inter3));
  inv1  gate1265(.a(s_103), .O(gate451inter4));
  nand2 gate1266(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate1267(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate1268(.a(G17), .O(gate451inter7));
  inv1  gate1269(.a(G1180), .O(gate451inter8));
  nand2 gate1270(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate1271(.a(s_103), .b(gate451inter3), .O(gate451inter10));
  nor2  gate1272(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate1273(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate1274(.a(gate451inter12), .b(gate451inter1), .O(G1260));
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );

  xor2  gate981(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate982(.a(gate454inter0), .b(s_62), .O(gate454inter1));
  and2  gate983(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate984(.a(s_62), .O(gate454inter3));
  inv1  gate985(.a(s_63), .O(gate454inter4));
  nand2 gate986(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate987(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate988(.a(G1087), .O(gate454inter7));
  inv1  gate989(.a(G1183), .O(gate454inter8));
  nand2 gate990(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate991(.a(s_63), .b(gate454inter3), .O(gate454inter10));
  nor2  gate992(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate993(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate994(.a(gate454inter12), .b(gate454inter1), .O(G1263));
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate1247(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate1248(.a(gate459inter0), .b(s_100), .O(gate459inter1));
  and2  gate1249(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate1250(.a(s_100), .O(gate459inter3));
  inv1  gate1251(.a(s_101), .O(gate459inter4));
  nand2 gate1252(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate1253(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate1254(.a(G21), .O(gate459inter7));
  inv1  gate1255(.a(G1192), .O(gate459inter8));
  nand2 gate1256(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate1257(.a(s_101), .b(gate459inter3), .O(gate459inter10));
  nor2  gate1258(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate1259(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate1260(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate1373(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate1374(.a(gate472inter0), .b(s_118), .O(gate472inter1));
  and2  gate1375(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate1376(.a(s_118), .O(gate472inter3));
  inv1  gate1377(.a(s_119), .O(gate472inter4));
  nand2 gate1378(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate1379(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate1380(.a(G1114), .O(gate472inter7));
  inv1  gate1381(.a(G1210), .O(gate472inter8));
  nand2 gate1382(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate1383(.a(s_119), .b(gate472inter3), .O(gate472inter10));
  nor2  gate1384(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate1385(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate1386(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate617(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate618(.a(gate485inter0), .b(s_10), .O(gate485inter1));
  and2  gate619(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate620(.a(s_10), .O(gate485inter3));
  inv1  gate621(.a(s_11), .O(gate485inter4));
  nand2 gate622(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate623(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate624(.a(G1232), .O(gate485inter7));
  inv1  gate625(.a(G1233), .O(gate485inter8));
  nand2 gate626(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate627(.a(s_11), .b(gate485inter3), .O(gate485inter10));
  nor2  gate628(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate629(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate630(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate1093(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate1094(.a(gate487inter0), .b(s_78), .O(gate487inter1));
  and2  gate1095(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate1096(.a(s_78), .O(gate487inter3));
  inv1  gate1097(.a(s_79), .O(gate487inter4));
  nand2 gate1098(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate1099(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate1100(.a(G1236), .O(gate487inter7));
  inv1  gate1101(.a(G1237), .O(gate487inter8));
  nand2 gate1102(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate1103(.a(s_79), .b(gate487inter3), .O(gate487inter10));
  nor2  gate1104(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate1105(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate1106(.a(gate487inter12), .b(gate487inter1), .O(G1296));
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate589(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate590(.a(gate489inter0), .b(s_6), .O(gate489inter1));
  and2  gate591(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate592(.a(s_6), .O(gate489inter3));
  inv1  gate593(.a(s_7), .O(gate489inter4));
  nand2 gate594(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate595(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate596(.a(G1240), .O(gate489inter7));
  inv1  gate597(.a(G1241), .O(gate489inter8));
  nand2 gate598(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate599(.a(s_7), .b(gate489inter3), .O(gate489inter10));
  nor2  gate600(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate601(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate602(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate967(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate968(.a(gate504inter0), .b(s_60), .O(gate504inter1));
  and2  gate969(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate970(.a(s_60), .O(gate504inter3));
  inv1  gate971(.a(s_61), .O(gate504inter4));
  nand2 gate972(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate973(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate974(.a(G1270), .O(gate504inter7));
  inv1  gate975(.a(G1271), .O(gate504inter8));
  nand2 gate976(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate977(.a(s_61), .b(gate504inter3), .O(gate504inter10));
  nor2  gate978(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate979(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate980(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule