module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );

  xor2  gate547(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate548(.a(gate10inter0), .b(s_0), .O(gate10inter1));
  and2  gate549(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate550(.a(s_0), .O(gate10inter3));
  inv1  gate551(.a(s_1), .O(gate10inter4));
  nand2 gate552(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate553(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate554(.a(G3), .O(gate10inter7));
  inv1  gate555(.a(G4), .O(gate10inter8));
  nand2 gate556(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate557(.a(s_1), .b(gate10inter3), .O(gate10inter10));
  nor2  gate558(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate559(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate560(.a(gate10inter12), .b(gate10inter1), .O(G269));
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );

  xor2  gate953(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate954(.a(gate14inter0), .b(s_58), .O(gate14inter1));
  and2  gate955(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate956(.a(s_58), .O(gate14inter3));
  inv1  gate957(.a(s_59), .O(gate14inter4));
  nand2 gate958(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate959(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate960(.a(G11), .O(gate14inter7));
  inv1  gate961(.a(G12), .O(gate14inter8));
  nand2 gate962(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate963(.a(s_59), .b(gate14inter3), .O(gate14inter10));
  nor2  gate964(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate965(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate966(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate1513(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate1514(.a(gate18inter0), .b(s_138), .O(gate18inter1));
  and2  gate1515(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate1516(.a(s_138), .O(gate18inter3));
  inv1  gate1517(.a(s_139), .O(gate18inter4));
  nand2 gate1518(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate1519(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate1520(.a(G19), .O(gate18inter7));
  inv1  gate1521(.a(G20), .O(gate18inter8));
  nand2 gate1522(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate1523(.a(s_139), .b(gate18inter3), .O(gate18inter10));
  nor2  gate1524(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate1525(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate1526(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate1527(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate1528(.a(gate27inter0), .b(s_140), .O(gate27inter1));
  and2  gate1529(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate1530(.a(s_140), .O(gate27inter3));
  inv1  gate1531(.a(s_141), .O(gate27inter4));
  nand2 gate1532(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate1533(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate1534(.a(G2), .O(gate27inter7));
  inv1  gate1535(.a(G6), .O(gate27inter8));
  nand2 gate1536(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate1537(.a(s_141), .b(gate27inter3), .O(gate27inter10));
  nor2  gate1538(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate1539(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate1540(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate1149(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate1150(.a(gate29inter0), .b(s_86), .O(gate29inter1));
  and2  gate1151(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate1152(.a(s_86), .O(gate29inter3));
  inv1  gate1153(.a(s_87), .O(gate29inter4));
  nand2 gate1154(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate1155(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate1156(.a(G3), .O(gate29inter7));
  inv1  gate1157(.a(G7), .O(gate29inter8));
  nand2 gate1158(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate1159(.a(s_87), .b(gate29inter3), .O(gate29inter10));
  nor2  gate1160(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate1161(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate1162(.a(gate29inter12), .b(gate29inter1), .O(G326));

  xor2  gate1303(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate1304(.a(gate30inter0), .b(s_108), .O(gate30inter1));
  and2  gate1305(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate1306(.a(s_108), .O(gate30inter3));
  inv1  gate1307(.a(s_109), .O(gate30inter4));
  nand2 gate1308(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate1309(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate1310(.a(G11), .O(gate30inter7));
  inv1  gate1311(.a(G15), .O(gate30inter8));
  nand2 gate1312(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate1313(.a(s_109), .b(gate30inter3), .O(gate30inter10));
  nor2  gate1314(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate1315(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate1316(.a(gate30inter12), .b(gate30inter1), .O(G329));
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate1415(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate1416(.a(gate38inter0), .b(s_124), .O(gate38inter1));
  and2  gate1417(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate1418(.a(s_124), .O(gate38inter3));
  inv1  gate1419(.a(s_125), .O(gate38inter4));
  nand2 gate1420(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate1421(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate1422(.a(G27), .O(gate38inter7));
  inv1  gate1423(.a(G31), .O(gate38inter8));
  nand2 gate1424(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate1425(.a(s_125), .b(gate38inter3), .O(gate38inter10));
  nor2  gate1426(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate1427(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate1428(.a(gate38inter12), .b(gate38inter1), .O(G353));
nand2 gate39( .a(G20), .b(G24), .O(G356) );

  xor2  gate925(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate926(.a(gate40inter0), .b(s_54), .O(gate40inter1));
  and2  gate927(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate928(.a(s_54), .O(gate40inter3));
  inv1  gate929(.a(s_55), .O(gate40inter4));
  nand2 gate930(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate931(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate932(.a(G28), .O(gate40inter7));
  inv1  gate933(.a(G32), .O(gate40inter8));
  nand2 gate934(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate935(.a(s_55), .b(gate40inter3), .O(gate40inter10));
  nor2  gate936(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate937(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate938(.a(gate40inter12), .b(gate40inter1), .O(G359));
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate603(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate604(.a(gate44inter0), .b(s_8), .O(gate44inter1));
  and2  gate605(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate606(.a(s_8), .O(gate44inter3));
  inv1  gate607(.a(s_9), .O(gate44inter4));
  nand2 gate608(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate609(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate610(.a(G4), .O(gate44inter7));
  inv1  gate611(.a(G269), .O(gate44inter8));
  nand2 gate612(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate613(.a(s_9), .b(gate44inter3), .O(gate44inter10));
  nor2  gate614(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate615(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate616(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate939(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate940(.a(gate58inter0), .b(s_56), .O(gate58inter1));
  and2  gate941(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate942(.a(s_56), .O(gate58inter3));
  inv1  gate943(.a(s_57), .O(gate58inter4));
  nand2 gate944(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate945(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate946(.a(G18), .O(gate58inter7));
  inv1  gate947(.a(G290), .O(gate58inter8));
  nand2 gate948(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate949(.a(s_57), .b(gate58inter3), .O(gate58inter10));
  nor2  gate950(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate951(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate952(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate1107(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate1108(.a(gate63inter0), .b(s_80), .O(gate63inter1));
  and2  gate1109(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate1110(.a(s_80), .O(gate63inter3));
  inv1  gate1111(.a(s_81), .O(gate63inter4));
  nand2 gate1112(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate1113(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate1114(.a(G23), .O(gate63inter7));
  inv1  gate1115(.a(G299), .O(gate63inter8));
  nand2 gate1116(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate1117(.a(s_81), .b(gate63inter3), .O(gate63inter10));
  nor2  gate1118(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate1119(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate1120(.a(gate63inter12), .b(gate63inter1), .O(G384));

  xor2  gate1009(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate1010(.a(gate64inter0), .b(s_66), .O(gate64inter1));
  and2  gate1011(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate1012(.a(s_66), .O(gate64inter3));
  inv1  gate1013(.a(s_67), .O(gate64inter4));
  nand2 gate1014(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate1015(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate1016(.a(G24), .O(gate64inter7));
  inv1  gate1017(.a(G299), .O(gate64inter8));
  nand2 gate1018(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate1019(.a(s_67), .b(gate64inter3), .O(gate64inter10));
  nor2  gate1020(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate1021(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate1022(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate1401(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate1402(.a(gate71inter0), .b(s_122), .O(gate71inter1));
  and2  gate1403(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate1404(.a(s_122), .O(gate71inter3));
  inv1  gate1405(.a(s_123), .O(gate71inter4));
  nand2 gate1406(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate1407(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate1408(.a(G31), .O(gate71inter7));
  inv1  gate1409(.a(G311), .O(gate71inter8));
  nand2 gate1410(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate1411(.a(s_123), .b(gate71inter3), .O(gate71inter10));
  nor2  gate1412(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate1413(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate1414(.a(gate71inter12), .b(gate71inter1), .O(G392));

  xor2  gate687(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate688(.a(gate72inter0), .b(s_20), .O(gate72inter1));
  and2  gate689(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate690(.a(s_20), .O(gate72inter3));
  inv1  gate691(.a(s_21), .O(gate72inter4));
  nand2 gate692(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate693(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate694(.a(G32), .O(gate72inter7));
  inv1  gate695(.a(G311), .O(gate72inter8));
  nand2 gate696(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate697(.a(s_21), .b(gate72inter3), .O(gate72inter10));
  nor2  gate698(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate699(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate700(.a(gate72inter12), .b(gate72inter1), .O(G393));
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate967(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate968(.a(gate78inter0), .b(s_60), .O(gate78inter1));
  and2  gate969(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate970(.a(s_60), .O(gate78inter3));
  inv1  gate971(.a(s_61), .O(gate78inter4));
  nand2 gate972(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate973(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate974(.a(G6), .O(gate78inter7));
  inv1  gate975(.a(G320), .O(gate78inter8));
  nand2 gate976(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate977(.a(s_61), .b(gate78inter3), .O(gate78inter10));
  nor2  gate978(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate979(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate980(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate1191(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate1192(.a(gate80inter0), .b(s_92), .O(gate80inter1));
  and2  gate1193(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate1194(.a(s_92), .O(gate80inter3));
  inv1  gate1195(.a(s_93), .O(gate80inter4));
  nand2 gate1196(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate1197(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate1198(.a(G14), .O(gate80inter7));
  inv1  gate1199(.a(G323), .O(gate80inter8));
  nand2 gate1200(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate1201(.a(s_93), .b(gate80inter3), .O(gate80inter10));
  nor2  gate1202(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate1203(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate1204(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate1317(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate1318(.a(gate94inter0), .b(s_110), .O(gate94inter1));
  and2  gate1319(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate1320(.a(s_110), .O(gate94inter3));
  inv1  gate1321(.a(s_111), .O(gate94inter4));
  nand2 gate1322(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate1323(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate1324(.a(G22), .O(gate94inter7));
  inv1  gate1325(.a(G344), .O(gate94inter8));
  nand2 gate1326(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate1327(.a(s_111), .b(gate94inter3), .O(gate94inter10));
  nor2  gate1328(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate1329(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate1330(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate1429(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate1430(.a(gate109inter0), .b(s_126), .O(gate109inter1));
  and2  gate1431(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate1432(.a(s_126), .O(gate109inter3));
  inv1  gate1433(.a(s_127), .O(gate109inter4));
  nand2 gate1434(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate1435(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate1436(.a(G370), .O(gate109inter7));
  inv1  gate1437(.a(G371), .O(gate109inter8));
  nand2 gate1438(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate1439(.a(s_127), .b(gate109inter3), .O(gate109inter10));
  nor2  gate1440(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate1441(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate1442(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate631(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate632(.a(gate112inter0), .b(s_12), .O(gate112inter1));
  and2  gate633(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate634(.a(s_12), .O(gate112inter3));
  inv1  gate635(.a(s_13), .O(gate112inter4));
  nand2 gate636(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate637(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate638(.a(G376), .O(gate112inter7));
  inv1  gate639(.a(G377), .O(gate112inter8));
  nand2 gate640(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate641(.a(s_13), .b(gate112inter3), .O(gate112inter10));
  nor2  gate642(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate643(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate644(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );

  xor2  gate827(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate828(.a(gate114inter0), .b(s_40), .O(gate114inter1));
  and2  gate829(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate830(.a(s_40), .O(gate114inter3));
  inv1  gate831(.a(s_41), .O(gate114inter4));
  nand2 gate832(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate833(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate834(.a(G380), .O(gate114inter7));
  inv1  gate835(.a(G381), .O(gate114inter8));
  nand2 gate836(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate837(.a(s_41), .b(gate114inter3), .O(gate114inter10));
  nor2  gate838(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate839(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate840(.a(gate114inter12), .b(gate114inter1), .O(G453));

  xor2  gate1569(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate1570(.a(gate115inter0), .b(s_146), .O(gate115inter1));
  and2  gate1571(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate1572(.a(s_146), .O(gate115inter3));
  inv1  gate1573(.a(s_147), .O(gate115inter4));
  nand2 gate1574(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate1575(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate1576(.a(G382), .O(gate115inter7));
  inv1  gate1577(.a(G383), .O(gate115inter8));
  nand2 gate1578(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate1579(.a(s_147), .b(gate115inter3), .O(gate115inter10));
  nor2  gate1580(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate1581(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate1582(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate1219(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate1220(.a(gate119inter0), .b(s_96), .O(gate119inter1));
  and2  gate1221(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate1222(.a(s_96), .O(gate119inter3));
  inv1  gate1223(.a(s_97), .O(gate119inter4));
  nand2 gate1224(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate1225(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate1226(.a(G390), .O(gate119inter7));
  inv1  gate1227(.a(G391), .O(gate119inter8));
  nand2 gate1228(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate1229(.a(s_97), .b(gate119inter3), .O(gate119inter10));
  nor2  gate1230(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate1231(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate1232(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate1065(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate1066(.a(gate123inter0), .b(s_74), .O(gate123inter1));
  and2  gate1067(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate1068(.a(s_74), .O(gate123inter3));
  inv1  gate1069(.a(s_75), .O(gate123inter4));
  nand2 gate1070(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate1071(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate1072(.a(G398), .O(gate123inter7));
  inv1  gate1073(.a(G399), .O(gate123inter8));
  nand2 gate1074(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate1075(.a(s_75), .b(gate123inter3), .O(gate123inter10));
  nor2  gate1076(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate1077(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate1078(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate1289(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate1290(.a(gate126inter0), .b(s_106), .O(gate126inter1));
  and2  gate1291(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate1292(.a(s_106), .O(gate126inter3));
  inv1  gate1293(.a(s_107), .O(gate126inter4));
  nand2 gate1294(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate1295(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate1296(.a(G404), .O(gate126inter7));
  inv1  gate1297(.a(G405), .O(gate126inter8));
  nand2 gate1298(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate1299(.a(s_107), .b(gate126inter3), .O(gate126inter10));
  nor2  gate1300(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate1301(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate1302(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate1457(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate1458(.a(gate130inter0), .b(s_130), .O(gate130inter1));
  and2  gate1459(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate1460(.a(s_130), .O(gate130inter3));
  inv1  gate1461(.a(s_131), .O(gate130inter4));
  nand2 gate1462(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate1463(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate1464(.a(G412), .O(gate130inter7));
  inv1  gate1465(.a(G413), .O(gate130inter8));
  nand2 gate1466(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate1467(.a(s_131), .b(gate130inter3), .O(gate130inter10));
  nor2  gate1468(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate1469(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate1470(.a(gate130inter12), .b(gate130inter1), .O(G501));
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate1373(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate1374(.a(gate132inter0), .b(s_118), .O(gate132inter1));
  and2  gate1375(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate1376(.a(s_118), .O(gate132inter3));
  inv1  gate1377(.a(s_119), .O(gate132inter4));
  nand2 gate1378(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate1379(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate1380(.a(G416), .O(gate132inter7));
  inv1  gate1381(.a(G417), .O(gate132inter8));
  nand2 gate1382(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate1383(.a(s_119), .b(gate132inter3), .O(gate132inter10));
  nor2  gate1384(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate1385(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate1386(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate1583(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate1584(.a(gate135inter0), .b(s_148), .O(gate135inter1));
  and2  gate1585(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate1586(.a(s_148), .O(gate135inter3));
  inv1  gate1587(.a(s_149), .O(gate135inter4));
  nand2 gate1588(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate1589(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate1590(.a(G422), .O(gate135inter7));
  inv1  gate1591(.a(G423), .O(gate135inter8));
  nand2 gate1592(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate1593(.a(s_149), .b(gate135inter3), .O(gate135inter10));
  nor2  gate1594(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate1595(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate1596(.a(gate135inter12), .b(gate135inter1), .O(G516));
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate1205(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate1206(.a(gate142inter0), .b(s_94), .O(gate142inter1));
  and2  gate1207(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate1208(.a(s_94), .O(gate142inter3));
  inv1  gate1209(.a(s_95), .O(gate142inter4));
  nand2 gate1210(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate1211(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate1212(.a(G456), .O(gate142inter7));
  inv1  gate1213(.a(G459), .O(gate142inter8));
  nand2 gate1214(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate1215(.a(s_95), .b(gate142inter3), .O(gate142inter10));
  nor2  gate1216(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate1217(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate1218(.a(gate142inter12), .b(gate142inter1), .O(G537));
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate869(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate870(.a(gate147inter0), .b(s_46), .O(gate147inter1));
  and2  gate871(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate872(.a(s_46), .O(gate147inter3));
  inv1  gate873(.a(s_47), .O(gate147inter4));
  nand2 gate874(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate875(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate876(.a(G486), .O(gate147inter7));
  inv1  gate877(.a(G489), .O(gate147inter8));
  nand2 gate878(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate879(.a(s_47), .b(gate147inter3), .O(gate147inter10));
  nor2  gate880(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate881(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate882(.a(gate147inter12), .b(gate147inter1), .O(G552));

  xor2  gate645(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate646(.a(gate148inter0), .b(s_14), .O(gate148inter1));
  and2  gate647(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate648(.a(s_14), .O(gate148inter3));
  inv1  gate649(.a(s_15), .O(gate148inter4));
  nand2 gate650(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate651(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate652(.a(G492), .O(gate148inter7));
  inv1  gate653(.a(G495), .O(gate148inter8));
  nand2 gate654(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate655(.a(s_15), .b(gate148inter3), .O(gate148inter10));
  nor2  gate656(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate657(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate658(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate617(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate618(.a(gate155inter0), .b(s_10), .O(gate155inter1));
  and2  gate619(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate620(.a(s_10), .O(gate155inter3));
  inv1  gate621(.a(s_11), .O(gate155inter4));
  nand2 gate622(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate623(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate624(.a(G432), .O(gate155inter7));
  inv1  gate625(.a(G525), .O(gate155inter8));
  nand2 gate626(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate627(.a(s_11), .b(gate155inter3), .O(gate155inter10));
  nor2  gate628(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate629(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate630(.a(gate155inter12), .b(gate155inter1), .O(G572));

  xor2  gate1555(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate1556(.a(gate156inter0), .b(s_144), .O(gate156inter1));
  and2  gate1557(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate1558(.a(s_144), .O(gate156inter3));
  inv1  gate1559(.a(s_145), .O(gate156inter4));
  nand2 gate1560(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate1561(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate1562(.a(G435), .O(gate156inter7));
  inv1  gate1563(.a(G525), .O(gate156inter8));
  nand2 gate1564(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate1565(.a(s_145), .b(gate156inter3), .O(gate156inter10));
  nor2  gate1566(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate1567(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate1568(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate743(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate744(.a(gate162inter0), .b(s_28), .O(gate162inter1));
  and2  gate745(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate746(.a(s_28), .O(gate162inter3));
  inv1  gate747(.a(s_29), .O(gate162inter4));
  nand2 gate748(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate749(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate750(.a(G453), .O(gate162inter7));
  inv1  gate751(.a(G534), .O(gate162inter8));
  nand2 gate752(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate753(.a(s_29), .b(gate162inter3), .O(gate162inter10));
  nor2  gate754(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate755(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate756(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate729(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate730(.a(gate170inter0), .b(s_26), .O(gate170inter1));
  and2  gate731(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate732(.a(s_26), .O(gate170inter3));
  inv1  gate733(.a(s_27), .O(gate170inter4));
  nand2 gate734(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate735(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate736(.a(G477), .O(gate170inter7));
  inv1  gate737(.a(G546), .O(gate170inter8));
  nand2 gate738(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate739(.a(s_27), .b(gate170inter3), .O(gate170inter10));
  nor2  gate740(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate741(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate742(.a(gate170inter12), .b(gate170inter1), .O(G587));

  xor2  gate883(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate884(.a(gate171inter0), .b(s_48), .O(gate171inter1));
  and2  gate885(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate886(.a(s_48), .O(gate171inter3));
  inv1  gate887(.a(s_49), .O(gate171inter4));
  nand2 gate888(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate889(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate890(.a(G480), .O(gate171inter7));
  inv1  gate891(.a(G549), .O(gate171inter8));
  nand2 gate892(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate893(.a(s_49), .b(gate171inter3), .O(gate171inter10));
  nor2  gate894(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate895(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate896(.a(gate171inter12), .b(gate171inter1), .O(G588));
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate1485(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate1486(.a(gate181inter0), .b(s_134), .O(gate181inter1));
  and2  gate1487(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate1488(.a(s_134), .O(gate181inter3));
  inv1  gate1489(.a(s_135), .O(gate181inter4));
  nand2 gate1490(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate1491(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate1492(.a(G510), .O(gate181inter7));
  inv1  gate1493(.a(G564), .O(gate181inter8));
  nand2 gate1494(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate1495(.a(s_135), .b(gate181inter3), .O(gate181inter10));
  nor2  gate1496(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate1497(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate1498(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate1331(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate1332(.a(gate188inter0), .b(s_112), .O(gate188inter1));
  and2  gate1333(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate1334(.a(s_112), .O(gate188inter3));
  inv1  gate1335(.a(s_113), .O(gate188inter4));
  nand2 gate1336(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate1337(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate1338(.a(G576), .O(gate188inter7));
  inv1  gate1339(.a(G577), .O(gate188inter8));
  nand2 gate1340(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate1341(.a(s_113), .b(gate188inter3), .O(gate188inter10));
  nor2  gate1342(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate1343(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate1344(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate1079(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate1080(.a(gate190inter0), .b(s_76), .O(gate190inter1));
  and2  gate1081(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate1082(.a(s_76), .O(gate190inter3));
  inv1  gate1083(.a(s_77), .O(gate190inter4));
  nand2 gate1084(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate1085(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate1086(.a(G580), .O(gate190inter7));
  inv1  gate1087(.a(G581), .O(gate190inter8));
  nand2 gate1088(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate1089(.a(s_77), .b(gate190inter3), .O(gate190inter10));
  nor2  gate1090(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate1091(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate1092(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate1541(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate1542(.a(gate196inter0), .b(s_142), .O(gate196inter1));
  and2  gate1543(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate1544(.a(s_142), .O(gate196inter3));
  inv1  gate1545(.a(s_143), .O(gate196inter4));
  nand2 gate1546(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate1547(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate1548(.a(G592), .O(gate196inter7));
  inv1  gate1549(.a(G593), .O(gate196inter8));
  nand2 gate1550(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate1551(.a(s_143), .b(gate196inter3), .O(gate196inter10));
  nor2  gate1552(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate1553(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate1554(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate981(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate982(.a(gate200inter0), .b(s_62), .O(gate200inter1));
  and2  gate983(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate984(.a(s_62), .O(gate200inter3));
  inv1  gate985(.a(s_63), .O(gate200inter4));
  nand2 gate986(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate987(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate988(.a(G600), .O(gate200inter7));
  inv1  gate989(.a(G601), .O(gate200inter8));
  nand2 gate990(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate991(.a(s_63), .b(gate200inter3), .O(gate200inter10));
  nor2  gate992(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate993(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate994(.a(gate200inter12), .b(gate200inter1), .O(G663));
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );

  xor2  gate1499(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate1500(.a(gate217inter0), .b(s_136), .O(gate217inter1));
  and2  gate1501(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate1502(.a(s_136), .O(gate217inter3));
  inv1  gate1503(.a(s_137), .O(gate217inter4));
  nand2 gate1504(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate1505(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate1506(.a(G622), .O(gate217inter7));
  inv1  gate1507(.a(G678), .O(gate217inter8));
  nand2 gate1508(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate1509(.a(s_137), .b(gate217inter3), .O(gate217inter10));
  nor2  gate1510(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate1511(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate1512(.a(gate217inter12), .b(gate217inter1), .O(G698));
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate673(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate674(.a(gate219inter0), .b(s_18), .O(gate219inter1));
  and2  gate675(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate676(.a(s_18), .O(gate219inter3));
  inv1  gate677(.a(s_19), .O(gate219inter4));
  nand2 gate678(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate679(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate680(.a(G632), .O(gate219inter7));
  inv1  gate681(.a(G681), .O(gate219inter8));
  nand2 gate682(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate683(.a(s_19), .b(gate219inter3), .O(gate219inter10));
  nor2  gate684(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate685(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate686(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate757(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate758(.a(gate241inter0), .b(s_30), .O(gate241inter1));
  and2  gate759(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate760(.a(s_30), .O(gate241inter3));
  inv1  gate761(.a(s_31), .O(gate241inter4));
  nand2 gate762(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate763(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate764(.a(G242), .O(gate241inter7));
  inv1  gate765(.a(G730), .O(gate241inter8));
  nand2 gate766(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate767(.a(s_31), .b(gate241inter3), .O(gate241inter10));
  nor2  gate768(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate769(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate770(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );

  xor2  gate841(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate842(.a(gate247inter0), .b(s_42), .O(gate247inter1));
  and2  gate843(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate844(.a(s_42), .O(gate247inter3));
  inv1  gate845(.a(s_43), .O(gate247inter4));
  nand2 gate846(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate847(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate848(.a(G251), .O(gate247inter7));
  inv1  gate849(.a(G739), .O(gate247inter8));
  nand2 gate850(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate851(.a(s_43), .b(gate247inter3), .O(gate247inter10));
  nor2  gate852(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate853(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate854(.a(gate247inter12), .b(gate247inter1), .O(G760));
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate715(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate716(.a(gate252inter0), .b(s_24), .O(gate252inter1));
  and2  gate717(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate718(.a(s_24), .O(gate252inter3));
  inv1  gate719(.a(s_25), .O(gate252inter4));
  nand2 gate720(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate721(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate722(.a(G709), .O(gate252inter7));
  inv1  gate723(.a(G745), .O(gate252inter8));
  nand2 gate724(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate725(.a(s_25), .b(gate252inter3), .O(gate252inter10));
  nor2  gate726(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate727(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate728(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate1177(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate1178(.a(gate255inter0), .b(s_90), .O(gate255inter1));
  and2  gate1179(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate1180(.a(s_90), .O(gate255inter3));
  inv1  gate1181(.a(s_91), .O(gate255inter4));
  nand2 gate1182(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate1183(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate1184(.a(G263), .O(gate255inter7));
  inv1  gate1185(.a(G751), .O(gate255inter8));
  nand2 gate1186(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate1187(.a(s_91), .b(gate255inter3), .O(gate255inter10));
  nor2  gate1188(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate1189(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate1190(.a(gate255inter12), .b(gate255inter1), .O(G768));

  xor2  gate911(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate912(.a(gate256inter0), .b(s_52), .O(gate256inter1));
  and2  gate913(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate914(.a(s_52), .O(gate256inter3));
  inv1  gate915(.a(s_53), .O(gate256inter4));
  nand2 gate916(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate917(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate918(.a(G715), .O(gate256inter7));
  inv1  gate919(.a(G751), .O(gate256inter8));
  nand2 gate920(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate921(.a(s_53), .b(gate256inter3), .O(gate256inter10));
  nor2  gate922(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate923(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate924(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate1261(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate1262(.a(gate263inter0), .b(s_102), .O(gate263inter1));
  and2  gate1263(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate1264(.a(s_102), .O(gate263inter3));
  inv1  gate1265(.a(s_103), .O(gate263inter4));
  nand2 gate1266(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate1267(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate1268(.a(G766), .O(gate263inter7));
  inv1  gate1269(.a(G767), .O(gate263inter8));
  nand2 gate1270(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate1271(.a(s_103), .b(gate263inter3), .O(gate263inter10));
  nor2  gate1272(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate1273(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate1274(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );

  xor2  gate1121(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate1122(.a(gate284inter0), .b(s_82), .O(gate284inter1));
  and2  gate1123(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate1124(.a(s_82), .O(gate284inter3));
  inv1  gate1125(.a(s_83), .O(gate284inter4));
  nand2 gate1126(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate1127(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate1128(.a(G785), .O(gate284inter7));
  inv1  gate1129(.a(G809), .O(gate284inter8));
  nand2 gate1130(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate1131(.a(s_83), .b(gate284inter3), .O(gate284inter10));
  nor2  gate1132(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate1133(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate1134(.a(gate284inter12), .b(gate284inter1), .O(G829));
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate575(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate576(.a(gate289inter0), .b(s_4), .O(gate289inter1));
  and2  gate577(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate578(.a(s_4), .O(gate289inter3));
  inv1  gate579(.a(s_5), .O(gate289inter4));
  nand2 gate580(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate581(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate582(.a(G818), .O(gate289inter7));
  inv1  gate583(.a(G819), .O(gate289inter8));
  nand2 gate584(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate585(.a(s_5), .b(gate289inter3), .O(gate289inter10));
  nor2  gate586(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate587(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate588(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate589(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate590(.a(gate293inter0), .b(s_6), .O(gate293inter1));
  and2  gate591(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate592(.a(s_6), .O(gate293inter3));
  inv1  gate593(.a(s_7), .O(gate293inter4));
  nand2 gate594(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate595(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate596(.a(G828), .O(gate293inter7));
  inv1  gate597(.a(G829), .O(gate293inter8));
  nand2 gate598(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate599(.a(s_7), .b(gate293inter3), .O(gate293inter10));
  nor2  gate600(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate601(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate602(.a(gate293inter12), .b(gate293inter1), .O(G886));

  xor2  gate897(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate898(.a(gate294inter0), .b(s_50), .O(gate294inter1));
  and2  gate899(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate900(.a(s_50), .O(gate294inter3));
  inv1  gate901(.a(s_51), .O(gate294inter4));
  nand2 gate902(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate903(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate904(.a(G832), .O(gate294inter7));
  inv1  gate905(.a(G833), .O(gate294inter8));
  nand2 gate906(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate907(.a(s_51), .b(gate294inter3), .O(gate294inter10));
  nor2  gate908(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate909(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate910(.a(gate294inter12), .b(gate294inter1), .O(G899));

  xor2  gate1345(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate1346(.a(gate295inter0), .b(s_114), .O(gate295inter1));
  and2  gate1347(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate1348(.a(s_114), .O(gate295inter3));
  inv1  gate1349(.a(s_115), .O(gate295inter4));
  nand2 gate1350(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate1351(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate1352(.a(G830), .O(gate295inter7));
  inv1  gate1353(.a(G831), .O(gate295inter8));
  nand2 gate1354(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate1355(.a(s_115), .b(gate295inter3), .O(gate295inter10));
  nor2  gate1356(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate1357(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate1358(.a(gate295inter12), .b(gate295inter1), .O(G912));

  xor2  gate659(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate660(.a(gate296inter0), .b(s_16), .O(gate296inter1));
  and2  gate661(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate662(.a(s_16), .O(gate296inter3));
  inv1  gate663(.a(s_17), .O(gate296inter4));
  nand2 gate664(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate665(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate666(.a(G826), .O(gate296inter7));
  inv1  gate667(.a(G827), .O(gate296inter8));
  nand2 gate668(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate669(.a(s_17), .b(gate296inter3), .O(gate296inter10));
  nor2  gate670(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate671(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate672(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate785(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate786(.a(gate389inter0), .b(s_34), .O(gate389inter1));
  and2  gate787(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate788(.a(s_34), .O(gate389inter3));
  inv1  gate789(.a(s_35), .O(gate389inter4));
  nand2 gate790(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate791(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate792(.a(G3), .O(gate389inter7));
  inv1  gate793(.a(G1042), .O(gate389inter8));
  nand2 gate794(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate795(.a(s_35), .b(gate389inter3), .O(gate389inter10));
  nor2  gate796(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate797(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate798(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate799(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate800(.a(gate398inter0), .b(s_36), .O(gate398inter1));
  and2  gate801(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate802(.a(s_36), .O(gate398inter3));
  inv1  gate803(.a(s_37), .O(gate398inter4));
  nand2 gate804(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate805(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate806(.a(G12), .O(gate398inter7));
  inv1  gate807(.a(G1069), .O(gate398inter8));
  nand2 gate808(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate809(.a(s_37), .b(gate398inter3), .O(gate398inter10));
  nor2  gate810(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate811(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate812(.a(gate398inter12), .b(gate398inter1), .O(G1165));

  xor2  gate1247(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate1248(.a(gate399inter0), .b(s_100), .O(gate399inter1));
  and2  gate1249(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate1250(.a(s_100), .O(gate399inter3));
  inv1  gate1251(.a(s_101), .O(gate399inter4));
  nand2 gate1252(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate1253(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate1254(.a(G13), .O(gate399inter7));
  inv1  gate1255(.a(G1072), .O(gate399inter8));
  nand2 gate1256(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate1257(.a(s_101), .b(gate399inter3), .O(gate399inter10));
  nor2  gate1258(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate1259(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate1260(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate1051(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate1052(.a(gate407inter0), .b(s_72), .O(gate407inter1));
  and2  gate1053(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate1054(.a(s_72), .O(gate407inter3));
  inv1  gate1055(.a(s_73), .O(gate407inter4));
  nand2 gate1056(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate1057(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate1058(.a(G21), .O(gate407inter7));
  inv1  gate1059(.a(G1096), .O(gate407inter8));
  nand2 gate1060(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate1061(.a(s_73), .b(gate407inter3), .O(gate407inter10));
  nor2  gate1062(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate1063(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate1064(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );

  xor2  gate1163(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate1164(.a(gate412inter0), .b(s_88), .O(gate412inter1));
  and2  gate1165(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate1166(.a(s_88), .O(gate412inter3));
  inv1  gate1167(.a(s_89), .O(gate412inter4));
  nand2 gate1168(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate1169(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate1170(.a(G26), .O(gate412inter7));
  inv1  gate1171(.a(G1111), .O(gate412inter8));
  nand2 gate1172(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate1173(.a(s_89), .b(gate412inter3), .O(gate412inter10));
  nor2  gate1174(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate1175(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate1176(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate1597(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1598(.a(gate420inter0), .b(s_150), .O(gate420inter1));
  and2  gate1599(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1600(.a(s_150), .O(gate420inter3));
  inv1  gate1601(.a(s_151), .O(gate420inter4));
  nand2 gate1602(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1603(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1604(.a(G1036), .O(gate420inter7));
  inv1  gate1605(.a(G1132), .O(gate420inter8));
  nand2 gate1606(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1607(.a(s_151), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1608(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1609(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1610(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate1037(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate1038(.a(gate425inter0), .b(s_70), .O(gate425inter1));
  and2  gate1039(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate1040(.a(s_70), .O(gate425inter3));
  inv1  gate1041(.a(s_71), .O(gate425inter4));
  nand2 gate1042(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1043(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1044(.a(G4), .O(gate425inter7));
  inv1  gate1045(.a(G1141), .O(gate425inter8));
  nand2 gate1046(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1047(.a(s_71), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1048(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1049(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1050(.a(gate425inter12), .b(gate425inter1), .O(G1234));
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate1135(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate1136(.a(gate441inter0), .b(s_84), .O(gate441inter1));
  and2  gate1137(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate1138(.a(s_84), .O(gate441inter3));
  inv1  gate1139(.a(s_85), .O(gate441inter4));
  nand2 gate1140(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate1141(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate1142(.a(G12), .O(gate441inter7));
  inv1  gate1143(.a(G1165), .O(gate441inter8));
  nand2 gate1144(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate1145(.a(s_85), .b(gate441inter3), .O(gate441inter10));
  nor2  gate1146(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate1147(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate1148(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate1233(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate1234(.a(gate444inter0), .b(s_98), .O(gate444inter1));
  and2  gate1235(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate1236(.a(s_98), .O(gate444inter3));
  inv1  gate1237(.a(s_99), .O(gate444inter4));
  nand2 gate1238(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate1239(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate1240(.a(G1072), .O(gate444inter7));
  inv1  gate1241(.a(G1168), .O(gate444inter8));
  nand2 gate1242(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate1243(.a(s_99), .b(gate444inter3), .O(gate444inter10));
  nor2  gate1244(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate1245(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate1246(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );

  xor2  gate1443(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate1444(.a(gate447inter0), .b(s_128), .O(gate447inter1));
  and2  gate1445(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate1446(.a(s_128), .O(gate447inter3));
  inv1  gate1447(.a(s_129), .O(gate447inter4));
  nand2 gate1448(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate1449(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate1450(.a(G15), .O(gate447inter7));
  inv1  gate1451(.a(G1174), .O(gate447inter8));
  nand2 gate1452(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate1453(.a(s_129), .b(gate447inter3), .O(gate447inter10));
  nor2  gate1454(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate1455(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate1456(.a(gate447inter12), .b(gate447inter1), .O(G1256));

  xor2  gate1471(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate1472(.a(gate448inter0), .b(s_132), .O(gate448inter1));
  and2  gate1473(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate1474(.a(s_132), .O(gate448inter3));
  inv1  gate1475(.a(s_133), .O(gate448inter4));
  nand2 gate1476(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate1477(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate1478(.a(G1078), .O(gate448inter7));
  inv1  gate1479(.a(G1174), .O(gate448inter8));
  nand2 gate1480(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate1481(.a(s_133), .b(gate448inter3), .O(gate448inter10));
  nor2  gate1482(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate1483(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate1484(.a(gate448inter12), .b(gate448inter1), .O(G1257));
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );

  xor2  gate561(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate562(.a(gate454inter0), .b(s_2), .O(gate454inter1));
  and2  gate563(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate564(.a(s_2), .O(gate454inter3));
  inv1  gate565(.a(s_3), .O(gate454inter4));
  nand2 gate566(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate567(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate568(.a(G1087), .O(gate454inter7));
  inv1  gate569(.a(G1183), .O(gate454inter8));
  nand2 gate570(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate571(.a(s_3), .b(gate454inter3), .O(gate454inter10));
  nor2  gate572(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate573(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate574(.a(gate454inter12), .b(gate454inter1), .O(G1263));

  xor2  gate1275(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate1276(.a(gate455inter0), .b(s_104), .O(gate455inter1));
  and2  gate1277(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate1278(.a(s_104), .O(gate455inter3));
  inv1  gate1279(.a(s_105), .O(gate455inter4));
  nand2 gate1280(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate1281(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate1282(.a(G19), .O(gate455inter7));
  inv1  gate1283(.a(G1186), .O(gate455inter8));
  nand2 gate1284(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate1285(.a(s_105), .b(gate455inter3), .O(gate455inter10));
  nor2  gate1286(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate1287(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate1288(.a(gate455inter12), .b(gate455inter1), .O(G1264));
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate855(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate856(.a(gate461inter0), .b(s_44), .O(gate461inter1));
  and2  gate857(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate858(.a(s_44), .O(gate461inter3));
  inv1  gate859(.a(s_45), .O(gate461inter4));
  nand2 gate860(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate861(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate862(.a(G22), .O(gate461inter7));
  inv1  gate863(.a(G1195), .O(gate461inter8));
  nand2 gate864(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate865(.a(s_45), .b(gate461inter3), .O(gate461inter10));
  nor2  gate866(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate867(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate868(.a(gate461inter12), .b(gate461inter1), .O(G1270));
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate1023(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate1024(.a(gate465inter0), .b(s_68), .O(gate465inter1));
  and2  gate1025(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate1026(.a(s_68), .O(gate465inter3));
  inv1  gate1027(.a(s_69), .O(gate465inter4));
  nand2 gate1028(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate1029(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate1030(.a(G24), .O(gate465inter7));
  inv1  gate1031(.a(G1201), .O(gate465inter8));
  nand2 gate1032(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate1033(.a(s_69), .b(gate465inter3), .O(gate465inter10));
  nor2  gate1034(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate1035(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate1036(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate1359(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate1360(.a(gate480inter0), .b(s_116), .O(gate480inter1));
  and2  gate1361(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate1362(.a(s_116), .O(gate480inter3));
  inv1  gate1363(.a(s_117), .O(gate480inter4));
  nand2 gate1364(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate1365(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate1366(.a(G1126), .O(gate480inter7));
  inv1  gate1367(.a(G1222), .O(gate480inter8));
  nand2 gate1368(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate1369(.a(s_117), .b(gate480inter3), .O(gate480inter10));
  nor2  gate1370(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate1371(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate1372(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate813(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate814(.a(gate487inter0), .b(s_38), .O(gate487inter1));
  and2  gate815(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate816(.a(s_38), .O(gate487inter3));
  inv1  gate817(.a(s_39), .O(gate487inter4));
  nand2 gate818(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate819(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate820(.a(G1236), .O(gate487inter7));
  inv1  gate821(.a(G1237), .O(gate487inter8));
  nand2 gate822(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate823(.a(s_39), .b(gate487inter3), .O(gate487inter10));
  nor2  gate824(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate825(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate826(.a(gate487inter12), .b(gate487inter1), .O(G1296));

  xor2  gate701(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate702(.a(gate488inter0), .b(s_22), .O(gate488inter1));
  and2  gate703(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate704(.a(s_22), .O(gate488inter3));
  inv1  gate705(.a(s_23), .O(gate488inter4));
  nand2 gate706(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate707(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate708(.a(G1238), .O(gate488inter7));
  inv1  gate709(.a(G1239), .O(gate488inter8));
  nand2 gate710(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate711(.a(s_23), .b(gate488inter3), .O(gate488inter10));
  nor2  gate712(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate713(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate714(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );

  xor2  gate1093(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate1094(.a(gate495inter0), .b(s_78), .O(gate495inter1));
  and2  gate1095(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate1096(.a(s_78), .O(gate495inter3));
  inv1  gate1097(.a(s_79), .O(gate495inter4));
  nand2 gate1098(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate1099(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate1100(.a(G1252), .O(gate495inter7));
  inv1  gate1101(.a(G1253), .O(gate495inter8));
  nand2 gate1102(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate1103(.a(s_79), .b(gate495inter3), .O(gate495inter10));
  nor2  gate1104(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate1105(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate1106(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate995(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate996(.a(gate504inter0), .b(s_64), .O(gate504inter1));
  and2  gate997(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate998(.a(s_64), .O(gate504inter3));
  inv1  gate999(.a(s_65), .O(gate504inter4));
  nand2 gate1000(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate1001(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate1002(.a(G1270), .O(gate504inter7));
  inv1  gate1003(.a(G1271), .O(gate504inter8));
  nand2 gate1004(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate1005(.a(s_65), .b(gate504inter3), .O(gate504inter10));
  nor2  gate1006(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate1007(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate1008(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate1387(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate1388(.a(gate510inter0), .b(s_120), .O(gate510inter1));
  and2  gate1389(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate1390(.a(s_120), .O(gate510inter3));
  inv1  gate1391(.a(s_121), .O(gate510inter4));
  nand2 gate1392(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate1393(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate1394(.a(G1282), .O(gate510inter7));
  inv1  gate1395(.a(G1283), .O(gate510inter8));
  nand2 gate1396(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate1397(.a(s_121), .b(gate510inter3), .O(gate510inter10));
  nor2  gate1398(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate1399(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate1400(.a(gate510inter12), .b(gate510inter1), .O(G1319));

  xor2  gate771(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate772(.a(gate511inter0), .b(s_32), .O(gate511inter1));
  and2  gate773(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate774(.a(s_32), .O(gate511inter3));
  inv1  gate775(.a(s_33), .O(gate511inter4));
  nand2 gate776(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate777(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate778(.a(G1284), .O(gate511inter7));
  inv1  gate779(.a(G1285), .O(gate511inter8));
  nand2 gate780(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate781(.a(s_33), .b(gate511inter3), .O(gate511inter10));
  nor2  gate782(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate783(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate784(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule