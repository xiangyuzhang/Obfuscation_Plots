module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate603(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate604(.a(gate15inter0), .b(s_8), .O(gate15inter1));
  and2  gate605(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate606(.a(s_8), .O(gate15inter3));
  inv1  gate607(.a(s_9), .O(gate15inter4));
  nand2 gate608(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate609(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate610(.a(G13), .O(gate15inter7));
  inv1  gate611(.a(G14), .O(gate15inter8));
  nand2 gate612(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate613(.a(s_9), .b(gate15inter3), .O(gate15inter10));
  nor2  gate614(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate615(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate616(.a(gate15inter12), .b(gate15inter1), .O(G284));

  xor2  gate1807(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate1808(.a(gate16inter0), .b(s_180), .O(gate16inter1));
  and2  gate1809(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate1810(.a(s_180), .O(gate16inter3));
  inv1  gate1811(.a(s_181), .O(gate16inter4));
  nand2 gate1812(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate1813(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate1814(.a(G15), .O(gate16inter7));
  inv1  gate1815(.a(G16), .O(gate16inter8));
  nand2 gate1816(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate1817(.a(s_181), .b(gate16inter3), .O(gate16inter10));
  nor2  gate1818(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate1819(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate1820(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate2493(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate2494(.a(gate20inter0), .b(s_278), .O(gate20inter1));
  and2  gate2495(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate2496(.a(s_278), .O(gate20inter3));
  inv1  gate2497(.a(s_279), .O(gate20inter4));
  nand2 gate2498(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate2499(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate2500(.a(G23), .O(gate20inter7));
  inv1  gate2501(.a(G24), .O(gate20inter8));
  nand2 gate2502(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate2503(.a(s_279), .b(gate20inter3), .O(gate20inter10));
  nor2  gate2504(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate2505(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate2506(.a(gate20inter12), .b(gate20inter1), .O(G299));

  xor2  gate2199(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate2200(.a(gate21inter0), .b(s_236), .O(gate21inter1));
  and2  gate2201(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate2202(.a(s_236), .O(gate21inter3));
  inv1  gate2203(.a(s_237), .O(gate21inter4));
  nand2 gate2204(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate2205(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate2206(.a(G25), .O(gate21inter7));
  inv1  gate2207(.a(G26), .O(gate21inter8));
  nand2 gate2208(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate2209(.a(s_237), .b(gate21inter3), .O(gate21inter10));
  nor2  gate2210(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate2211(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate2212(.a(gate21inter12), .b(gate21inter1), .O(G302));

  xor2  gate1345(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate1346(.a(gate22inter0), .b(s_114), .O(gate22inter1));
  and2  gate1347(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate1348(.a(s_114), .O(gate22inter3));
  inv1  gate1349(.a(s_115), .O(gate22inter4));
  nand2 gate1350(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate1351(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate1352(.a(G27), .O(gate22inter7));
  inv1  gate1353(.a(G28), .O(gate22inter8));
  nand2 gate1354(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate1355(.a(s_115), .b(gate22inter3), .O(gate22inter10));
  nor2  gate1356(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate1357(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate1358(.a(gate22inter12), .b(gate22inter1), .O(G305));
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate785(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate786(.a(gate24inter0), .b(s_34), .O(gate24inter1));
  and2  gate787(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate788(.a(s_34), .O(gate24inter3));
  inv1  gate789(.a(s_35), .O(gate24inter4));
  nand2 gate790(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate791(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate792(.a(G31), .O(gate24inter7));
  inv1  gate793(.a(G32), .O(gate24inter8));
  nand2 gate794(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate795(.a(s_35), .b(gate24inter3), .O(gate24inter10));
  nor2  gate796(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate797(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate798(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate2311(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate2312(.a(gate28inter0), .b(s_252), .O(gate28inter1));
  and2  gate2313(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate2314(.a(s_252), .O(gate28inter3));
  inv1  gate2315(.a(s_253), .O(gate28inter4));
  nand2 gate2316(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate2317(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate2318(.a(G10), .O(gate28inter7));
  inv1  gate2319(.a(G14), .O(gate28inter8));
  nand2 gate2320(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate2321(.a(s_253), .b(gate28inter3), .O(gate28inter10));
  nor2  gate2322(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate2323(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate2324(.a(gate28inter12), .b(gate28inter1), .O(G323));
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate743(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate744(.a(gate37inter0), .b(s_28), .O(gate37inter1));
  and2  gate745(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate746(.a(s_28), .O(gate37inter3));
  inv1  gate747(.a(s_29), .O(gate37inter4));
  nand2 gate748(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate749(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate750(.a(G19), .O(gate37inter7));
  inv1  gate751(.a(G23), .O(gate37inter8));
  nand2 gate752(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate753(.a(s_29), .b(gate37inter3), .O(gate37inter10));
  nor2  gate754(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate755(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate756(.a(gate37inter12), .b(gate37inter1), .O(G350));

  xor2  gate1107(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate1108(.a(gate38inter0), .b(s_80), .O(gate38inter1));
  and2  gate1109(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate1110(.a(s_80), .O(gate38inter3));
  inv1  gate1111(.a(s_81), .O(gate38inter4));
  nand2 gate1112(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate1113(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate1114(.a(G27), .O(gate38inter7));
  inv1  gate1115(.a(G31), .O(gate38inter8));
  nand2 gate1116(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate1117(.a(s_81), .b(gate38inter3), .O(gate38inter10));
  nor2  gate1118(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate1119(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate1120(.a(gate38inter12), .b(gate38inter1), .O(G353));
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );

  xor2  gate2395(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate2396(.a(gate42inter0), .b(s_264), .O(gate42inter1));
  and2  gate2397(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate2398(.a(s_264), .O(gate42inter3));
  inv1  gate2399(.a(s_265), .O(gate42inter4));
  nand2 gate2400(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate2401(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate2402(.a(G2), .O(gate42inter7));
  inv1  gate2403(.a(G266), .O(gate42inter8));
  nand2 gate2404(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate2405(.a(s_265), .b(gate42inter3), .O(gate42inter10));
  nor2  gate2406(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate2407(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate2408(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate1121(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate1122(.a(gate46inter0), .b(s_82), .O(gate46inter1));
  and2  gate1123(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate1124(.a(s_82), .O(gate46inter3));
  inv1  gate1125(.a(s_83), .O(gate46inter4));
  nand2 gate1126(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate1127(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate1128(.a(G6), .O(gate46inter7));
  inv1  gate1129(.a(G272), .O(gate46inter8));
  nand2 gate1130(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate1131(.a(s_83), .b(gate46inter3), .O(gate46inter10));
  nor2  gate1132(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate1133(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate1134(.a(gate46inter12), .b(gate46inter1), .O(G367));

  xor2  gate897(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate898(.a(gate47inter0), .b(s_50), .O(gate47inter1));
  and2  gate899(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate900(.a(s_50), .O(gate47inter3));
  inv1  gate901(.a(s_51), .O(gate47inter4));
  nand2 gate902(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate903(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate904(.a(G7), .O(gate47inter7));
  inv1  gate905(.a(G275), .O(gate47inter8));
  nand2 gate906(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate907(.a(s_51), .b(gate47inter3), .O(gate47inter10));
  nor2  gate908(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate909(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate910(.a(gate47inter12), .b(gate47inter1), .O(G368));
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate981(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate982(.a(gate55inter0), .b(s_62), .O(gate55inter1));
  and2  gate983(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate984(.a(s_62), .O(gate55inter3));
  inv1  gate985(.a(s_63), .O(gate55inter4));
  nand2 gate986(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate987(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate988(.a(G15), .O(gate55inter7));
  inv1  gate989(.a(G287), .O(gate55inter8));
  nand2 gate990(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate991(.a(s_63), .b(gate55inter3), .O(gate55inter10));
  nor2  gate992(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate993(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate994(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate1499(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate1500(.a(gate59inter0), .b(s_136), .O(gate59inter1));
  and2  gate1501(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate1502(.a(s_136), .O(gate59inter3));
  inv1  gate1503(.a(s_137), .O(gate59inter4));
  nand2 gate1504(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate1505(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate1506(.a(G19), .O(gate59inter7));
  inv1  gate1507(.a(G293), .O(gate59inter8));
  nand2 gate1508(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate1509(.a(s_137), .b(gate59inter3), .O(gate59inter10));
  nor2  gate1510(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate1511(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate1512(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate1555(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate1556(.a(gate62inter0), .b(s_144), .O(gate62inter1));
  and2  gate1557(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate1558(.a(s_144), .O(gate62inter3));
  inv1  gate1559(.a(s_145), .O(gate62inter4));
  nand2 gate1560(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate1561(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate1562(.a(G22), .O(gate62inter7));
  inv1  gate1563(.a(G296), .O(gate62inter8));
  nand2 gate1564(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate1565(.a(s_145), .b(gate62inter3), .O(gate62inter10));
  nor2  gate1566(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate1567(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate1568(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate1051(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate1052(.a(gate65inter0), .b(s_72), .O(gate65inter1));
  and2  gate1053(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate1054(.a(s_72), .O(gate65inter3));
  inv1  gate1055(.a(s_73), .O(gate65inter4));
  nand2 gate1056(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate1057(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate1058(.a(G25), .O(gate65inter7));
  inv1  gate1059(.a(G302), .O(gate65inter8));
  nand2 gate1060(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate1061(.a(s_73), .b(gate65inter3), .O(gate65inter10));
  nor2  gate1062(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate1063(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate1064(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate2157(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate2158(.a(gate69inter0), .b(s_230), .O(gate69inter1));
  and2  gate2159(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate2160(.a(s_230), .O(gate69inter3));
  inv1  gate2161(.a(s_231), .O(gate69inter4));
  nand2 gate2162(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate2163(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate2164(.a(G29), .O(gate69inter7));
  inv1  gate2165(.a(G308), .O(gate69inter8));
  nand2 gate2166(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate2167(.a(s_231), .b(gate69inter3), .O(gate69inter10));
  nor2  gate2168(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate2169(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate2170(.a(gate69inter12), .b(gate69inter1), .O(G390));

  xor2  gate1037(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate1038(.a(gate70inter0), .b(s_70), .O(gate70inter1));
  and2  gate1039(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate1040(.a(s_70), .O(gate70inter3));
  inv1  gate1041(.a(s_71), .O(gate70inter4));
  nand2 gate1042(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate1043(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate1044(.a(G30), .O(gate70inter7));
  inv1  gate1045(.a(G308), .O(gate70inter8));
  nand2 gate1046(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate1047(.a(s_71), .b(gate70inter3), .O(gate70inter10));
  nor2  gate1048(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate1049(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate1050(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );

  xor2  gate2269(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate2270(.a(gate72inter0), .b(s_246), .O(gate72inter1));
  and2  gate2271(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate2272(.a(s_246), .O(gate72inter3));
  inv1  gate2273(.a(s_247), .O(gate72inter4));
  nand2 gate2274(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate2275(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate2276(.a(G32), .O(gate72inter7));
  inv1  gate2277(.a(G311), .O(gate72inter8));
  nand2 gate2278(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate2279(.a(s_247), .b(gate72inter3), .O(gate72inter10));
  nor2  gate2280(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate2281(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate2282(.a(gate72inter12), .b(gate72inter1), .O(G393));

  xor2  gate617(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate618(.a(gate73inter0), .b(s_10), .O(gate73inter1));
  and2  gate619(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate620(.a(s_10), .O(gate73inter3));
  inv1  gate621(.a(s_11), .O(gate73inter4));
  nand2 gate622(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate623(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate624(.a(G1), .O(gate73inter7));
  inv1  gate625(.a(G314), .O(gate73inter8));
  nand2 gate626(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate627(.a(s_11), .b(gate73inter3), .O(gate73inter10));
  nor2  gate628(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate629(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate630(.a(gate73inter12), .b(gate73inter1), .O(G394));

  xor2  gate813(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate814(.a(gate74inter0), .b(s_38), .O(gate74inter1));
  and2  gate815(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate816(.a(s_38), .O(gate74inter3));
  inv1  gate817(.a(s_39), .O(gate74inter4));
  nand2 gate818(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate819(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate820(.a(G5), .O(gate74inter7));
  inv1  gate821(.a(G314), .O(gate74inter8));
  nand2 gate822(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate823(.a(s_39), .b(gate74inter3), .O(gate74inter10));
  nor2  gate824(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate825(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate826(.a(gate74inter12), .b(gate74inter1), .O(G395));

  xor2  gate1331(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate1332(.a(gate75inter0), .b(s_112), .O(gate75inter1));
  and2  gate1333(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate1334(.a(s_112), .O(gate75inter3));
  inv1  gate1335(.a(s_113), .O(gate75inter4));
  nand2 gate1336(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate1337(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate1338(.a(G9), .O(gate75inter7));
  inv1  gate1339(.a(G317), .O(gate75inter8));
  nand2 gate1340(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate1341(.a(s_113), .b(gate75inter3), .O(gate75inter10));
  nor2  gate1342(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate1343(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate1344(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate1653(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate1654(.a(gate80inter0), .b(s_158), .O(gate80inter1));
  and2  gate1655(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate1656(.a(s_158), .O(gate80inter3));
  inv1  gate1657(.a(s_159), .O(gate80inter4));
  nand2 gate1658(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate1659(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate1660(.a(G14), .O(gate80inter7));
  inv1  gate1661(.a(G323), .O(gate80inter8));
  nand2 gate1662(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate1663(.a(s_159), .b(gate80inter3), .O(gate80inter10));
  nor2  gate1664(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate1665(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate1666(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate2409(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate2410(.a(gate82inter0), .b(s_266), .O(gate82inter1));
  and2  gate2411(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate2412(.a(s_266), .O(gate82inter3));
  inv1  gate2413(.a(s_267), .O(gate82inter4));
  nand2 gate2414(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate2415(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate2416(.a(G7), .O(gate82inter7));
  inv1  gate2417(.a(G326), .O(gate82inter8));
  nand2 gate2418(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate2419(.a(s_267), .b(gate82inter3), .O(gate82inter10));
  nor2  gate2420(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate2421(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate2422(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate1821(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate1822(.a(gate86inter0), .b(s_182), .O(gate86inter1));
  and2  gate1823(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate1824(.a(s_182), .O(gate86inter3));
  inv1  gate1825(.a(s_183), .O(gate86inter4));
  nand2 gate1826(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate1827(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate1828(.a(G8), .O(gate86inter7));
  inv1  gate1829(.a(G332), .O(gate86inter8));
  nand2 gate1830(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate1831(.a(s_183), .b(gate86inter3), .O(gate86inter10));
  nor2  gate1832(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate1833(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate1834(.a(gate86inter12), .b(gate86inter1), .O(G407));

  xor2  gate757(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate758(.a(gate87inter0), .b(s_30), .O(gate87inter1));
  and2  gate759(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate760(.a(s_30), .O(gate87inter3));
  inv1  gate761(.a(s_31), .O(gate87inter4));
  nand2 gate762(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate763(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate764(.a(G12), .O(gate87inter7));
  inv1  gate765(.a(G335), .O(gate87inter8));
  nand2 gate766(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate767(.a(s_31), .b(gate87inter3), .O(gate87inter10));
  nor2  gate768(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate769(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate770(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );

  xor2  gate2003(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate2004(.a(gate89inter0), .b(s_208), .O(gate89inter1));
  and2  gate2005(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate2006(.a(s_208), .O(gate89inter3));
  inv1  gate2007(.a(s_209), .O(gate89inter4));
  nand2 gate2008(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate2009(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate2010(.a(G17), .O(gate89inter7));
  inv1  gate2011(.a(G338), .O(gate89inter8));
  nand2 gate2012(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate2013(.a(s_209), .b(gate89inter3), .O(gate89inter10));
  nor2  gate2014(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate2015(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate2016(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate2129(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate2130(.a(gate104inter0), .b(s_226), .O(gate104inter1));
  and2  gate2131(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate2132(.a(s_226), .O(gate104inter3));
  inv1  gate2133(.a(s_227), .O(gate104inter4));
  nand2 gate2134(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate2135(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate2136(.a(G32), .O(gate104inter7));
  inv1  gate2137(.a(G359), .O(gate104inter8));
  nand2 gate2138(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate2139(.a(s_227), .b(gate104inter3), .O(gate104inter10));
  nor2  gate2140(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate2141(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate2142(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate1485(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate1486(.a(gate108inter0), .b(s_134), .O(gate108inter1));
  and2  gate1487(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate1488(.a(s_134), .O(gate108inter3));
  inv1  gate1489(.a(s_135), .O(gate108inter4));
  nand2 gate1490(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate1491(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate1492(.a(G368), .O(gate108inter7));
  inv1  gate1493(.a(G369), .O(gate108inter8));
  nand2 gate1494(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate1495(.a(s_135), .b(gate108inter3), .O(gate108inter10));
  nor2  gate1496(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate1497(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate1498(.a(gate108inter12), .b(gate108inter1), .O(G435));
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate939(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate940(.a(gate110inter0), .b(s_56), .O(gate110inter1));
  and2  gate941(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate942(.a(s_56), .O(gate110inter3));
  inv1  gate943(.a(s_57), .O(gate110inter4));
  nand2 gate944(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate945(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate946(.a(G372), .O(gate110inter7));
  inv1  gate947(.a(G373), .O(gate110inter8));
  nand2 gate948(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate949(.a(s_57), .b(gate110inter3), .O(gate110inter10));
  nor2  gate950(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate951(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate952(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate2101(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate2102(.a(gate117inter0), .b(s_222), .O(gate117inter1));
  and2  gate2103(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate2104(.a(s_222), .O(gate117inter3));
  inv1  gate2105(.a(s_223), .O(gate117inter4));
  nand2 gate2106(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate2107(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate2108(.a(G386), .O(gate117inter7));
  inv1  gate2109(.a(G387), .O(gate117inter8));
  nand2 gate2110(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate2111(.a(s_223), .b(gate117inter3), .O(gate117inter10));
  nor2  gate2112(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate2113(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate2114(.a(gate117inter12), .b(gate117inter1), .O(G462));

  xor2  gate911(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate912(.a(gate118inter0), .b(s_52), .O(gate118inter1));
  and2  gate913(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate914(.a(s_52), .O(gate118inter3));
  inv1  gate915(.a(s_53), .O(gate118inter4));
  nand2 gate916(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate917(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate918(.a(G388), .O(gate118inter7));
  inv1  gate919(.a(G389), .O(gate118inter8));
  nand2 gate920(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate921(.a(s_53), .b(gate118inter3), .O(gate118inter10));
  nor2  gate922(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate923(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate924(.a(gate118inter12), .b(gate118inter1), .O(G465));
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );

  xor2  gate2353(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate2354(.a(gate122inter0), .b(s_258), .O(gate122inter1));
  and2  gate2355(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate2356(.a(s_258), .O(gate122inter3));
  inv1  gate2357(.a(s_259), .O(gate122inter4));
  nand2 gate2358(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate2359(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate2360(.a(G396), .O(gate122inter7));
  inv1  gate2361(.a(G397), .O(gate122inter8));
  nand2 gate2362(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate2363(.a(s_259), .b(gate122inter3), .O(gate122inter10));
  nor2  gate2364(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate2365(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate2366(.a(gate122inter12), .b(gate122inter1), .O(G477));
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate1667(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate1668(.a(gate124inter0), .b(s_160), .O(gate124inter1));
  and2  gate1669(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate1670(.a(s_160), .O(gate124inter3));
  inv1  gate1671(.a(s_161), .O(gate124inter4));
  nand2 gate1672(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate1673(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate1674(.a(G400), .O(gate124inter7));
  inv1  gate1675(.a(G401), .O(gate124inter8));
  nand2 gate1676(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate1677(.a(s_161), .b(gate124inter3), .O(gate124inter10));
  nor2  gate1678(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate1679(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate1680(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate1135(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate1136(.a(gate130inter0), .b(s_84), .O(gate130inter1));
  and2  gate1137(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate1138(.a(s_84), .O(gate130inter3));
  inv1  gate1139(.a(s_85), .O(gate130inter4));
  nand2 gate1140(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate1141(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate1142(.a(G412), .O(gate130inter7));
  inv1  gate1143(.a(G413), .O(gate130inter8));
  nand2 gate1144(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate1145(.a(s_85), .b(gate130inter3), .O(gate130inter10));
  nor2  gate1146(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate1147(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate1148(.a(gate130inter12), .b(gate130inter1), .O(G501));

  xor2  gate1597(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate1598(.a(gate131inter0), .b(s_150), .O(gate131inter1));
  and2  gate1599(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate1600(.a(s_150), .O(gate131inter3));
  inv1  gate1601(.a(s_151), .O(gate131inter4));
  nand2 gate1602(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate1603(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate1604(.a(G414), .O(gate131inter7));
  inv1  gate1605(.a(G415), .O(gate131inter8));
  nand2 gate1606(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate1607(.a(s_151), .b(gate131inter3), .O(gate131inter10));
  nor2  gate1608(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate1609(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate1610(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate2241(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate2242(.a(gate138inter0), .b(s_242), .O(gate138inter1));
  and2  gate2243(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate2244(.a(s_242), .O(gate138inter3));
  inv1  gate2245(.a(s_243), .O(gate138inter4));
  nand2 gate2246(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate2247(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate2248(.a(G432), .O(gate138inter7));
  inv1  gate2249(.a(G435), .O(gate138inter8));
  nand2 gate2250(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate2251(.a(s_243), .b(gate138inter3), .O(gate138inter10));
  nor2  gate2252(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate2253(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate2254(.a(gate138inter12), .b(gate138inter1), .O(G525));

  xor2  gate1443(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate1444(.a(gate139inter0), .b(s_128), .O(gate139inter1));
  and2  gate1445(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate1446(.a(s_128), .O(gate139inter3));
  inv1  gate1447(.a(s_129), .O(gate139inter4));
  nand2 gate1448(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate1449(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate1450(.a(G438), .O(gate139inter7));
  inv1  gate1451(.a(G441), .O(gate139inter8));
  nand2 gate1452(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate1453(.a(s_129), .b(gate139inter3), .O(gate139inter10));
  nor2  gate1454(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate1455(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate1456(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );

  xor2  gate2227(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate2228(.a(gate146inter0), .b(s_240), .O(gate146inter1));
  and2  gate2229(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate2230(.a(s_240), .O(gate146inter3));
  inv1  gate2231(.a(s_241), .O(gate146inter4));
  nand2 gate2232(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate2233(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate2234(.a(G480), .O(gate146inter7));
  inv1  gate2235(.a(G483), .O(gate146inter8));
  nand2 gate2236(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate2237(.a(s_241), .b(gate146inter3), .O(gate146inter10));
  nor2  gate2238(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate2239(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate2240(.a(gate146inter12), .b(gate146inter1), .O(G549));
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate1317(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1318(.a(gate148inter0), .b(s_110), .O(gate148inter1));
  and2  gate1319(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1320(.a(s_110), .O(gate148inter3));
  inv1  gate1321(.a(s_111), .O(gate148inter4));
  nand2 gate1322(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1323(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1324(.a(G492), .O(gate148inter7));
  inv1  gate1325(.a(G495), .O(gate148inter8));
  nand2 gate1326(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1327(.a(s_111), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1328(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1329(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1330(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate2115(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate2116(.a(gate157inter0), .b(s_224), .O(gate157inter1));
  and2  gate2117(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate2118(.a(s_224), .O(gate157inter3));
  inv1  gate2119(.a(s_225), .O(gate157inter4));
  nand2 gate2120(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate2121(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate2122(.a(G438), .O(gate157inter7));
  inv1  gate2123(.a(G528), .O(gate157inter8));
  nand2 gate2124(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate2125(.a(s_225), .b(gate157inter3), .O(gate157inter10));
  nor2  gate2126(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate2127(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate2128(.a(gate157inter12), .b(gate157inter1), .O(G574));

  xor2  gate1933(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate1934(.a(gate158inter0), .b(s_198), .O(gate158inter1));
  and2  gate1935(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate1936(.a(s_198), .O(gate158inter3));
  inv1  gate1937(.a(s_199), .O(gate158inter4));
  nand2 gate1938(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate1939(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate1940(.a(G441), .O(gate158inter7));
  inv1  gate1941(.a(G528), .O(gate158inter8));
  nand2 gate1942(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate1943(.a(s_199), .b(gate158inter3), .O(gate158inter10));
  nor2  gate1944(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate1945(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate1946(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate1583(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate1584(.a(gate160inter0), .b(s_148), .O(gate160inter1));
  and2  gate1585(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate1586(.a(s_148), .O(gate160inter3));
  inv1  gate1587(.a(s_149), .O(gate160inter4));
  nand2 gate1588(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate1589(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate1590(.a(G447), .O(gate160inter7));
  inv1  gate1591(.a(G531), .O(gate160inter8));
  nand2 gate1592(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate1593(.a(s_149), .b(gate160inter3), .O(gate160inter10));
  nor2  gate1594(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate1595(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate1596(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate1891(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate1892(.a(gate162inter0), .b(s_192), .O(gate162inter1));
  and2  gate1893(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate1894(.a(s_192), .O(gate162inter3));
  inv1  gate1895(.a(s_193), .O(gate162inter4));
  nand2 gate1896(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate1897(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate1898(.a(G453), .O(gate162inter7));
  inv1  gate1899(.a(G534), .O(gate162inter8));
  nand2 gate1900(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate1901(.a(s_193), .b(gate162inter3), .O(gate162inter10));
  nor2  gate1902(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate1903(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate1904(.a(gate162inter12), .b(gate162inter1), .O(G579));

  xor2  gate2171(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate2172(.a(gate163inter0), .b(s_232), .O(gate163inter1));
  and2  gate2173(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate2174(.a(s_232), .O(gate163inter3));
  inv1  gate2175(.a(s_233), .O(gate163inter4));
  nand2 gate2176(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate2177(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate2178(.a(G456), .O(gate163inter7));
  inv1  gate2179(.a(G537), .O(gate163inter8));
  nand2 gate2180(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate2181(.a(s_233), .b(gate163inter3), .O(gate163inter10));
  nor2  gate2182(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate2183(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate2184(.a(gate163inter12), .b(gate163inter1), .O(G580));

  xor2  gate2367(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate2368(.a(gate164inter0), .b(s_260), .O(gate164inter1));
  and2  gate2369(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate2370(.a(s_260), .O(gate164inter3));
  inv1  gate2371(.a(s_261), .O(gate164inter4));
  nand2 gate2372(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate2373(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate2374(.a(G459), .O(gate164inter7));
  inv1  gate2375(.a(G537), .O(gate164inter8));
  nand2 gate2376(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate2377(.a(s_261), .b(gate164inter3), .O(gate164inter10));
  nor2  gate2378(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate2379(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate2380(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );

  xor2  gate827(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate828(.a(gate166inter0), .b(s_40), .O(gate166inter1));
  and2  gate829(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate830(.a(s_40), .O(gate166inter3));
  inv1  gate831(.a(s_41), .O(gate166inter4));
  nand2 gate832(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate833(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate834(.a(G465), .O(gate166inter7));
  inv1  gate835(.a(G540), .O(gate166inter8));
  nand2 gate836(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate837(.a(s_41), .b(gate166inter3), .O(gate166inter10));
  nor2  gate838(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate839(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate840(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate1471(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate1472(.a(gate174inter0), .b(s_132), .O(gate174inter1));
  and2  gate1473(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate1474(.a(s_132), .O(gate174inter3));
  inv1  gate1475(.a(s_133), .O(gate174inter4));
  nand2 gate1476(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate1477(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate1478(.a(G489), .O(gate174inter7));
  inv1  gate1479(.a(G552), .O(gate174inter8));
  nand2 gate1480(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate1481(.a(s_133), .b(gate174inter3), .O(gate174inter10));
  nor2  gate1482(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate1483(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate1484(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );

  xor2  gate1723(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate1724(.a(gate176inter0), .b(s_168), .O(gate176inter1));
  and2  gate1725(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate1726(.a(s_168), .O(gate176inter3));
  inv1  gate1727(.a(s_169), .O(gate176inter4));
  nand2 gate1728(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate1729(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate1730(.a(G495), .O(gate176inter7));
  inv1  gate1731(.a(G555), .O(gate176inter8));
  nand2 gate1732(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate1733(.a(s_169), .b(gate176inter3), .O(gate176inter10));
  nor2  gate1734(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate1735(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate1736(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate1919(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate1920(.a(gate180inter0), .b(s_196), .O(gate180inter1));
  and2  gate1921(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate1922(.a(s_196), .O(gate180inter3));
  inv1  gate1923(.a(s_197), .O(gate180inter4));
  nand2 gate1924(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate1925(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate1926(.a(G507), .O(gate180inter7));
  inv1  gate1927(.a(G561), .O(gate180inter8));
  nand2 gate1928(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate1929(.a(s_197), .b(gate180inter3), .O(gate180inter10));
  nor2  gate1930(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate1931(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate1932(.a(gate180inter12), .b(gate180inter1), .O(G597));
nand2 gate181( .a(G510), .b(G564), .O(G598) );

  xor2  gate575(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate576(.a(gate182inter0), .b(s_4), .O(gate182inter1));
  and2  gate577(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate578(.a(s_4), .O(gate182inter3));
  inv1  gate579(.a(s_5), .O(gate182inter4));
  nand2 gate580(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate581(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate582(.a(G513), .O(gate182inter7));
  inv1  gate583(.a(G564), .O(gate182inter8));
  nand2 gate584(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate585(.a(s_5), .b(gate182inter3), .O(gate182inter10));
  nor2  gate586(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate587(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate588(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate995(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate996(.a(gate185inter0), .b(s_64), .O(gate185inter1));
  and2  gate997(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate998(.a(s_64), .O(gate185inter3));
  inv1  gate999(.a(s_65), .O(gate185inter4));
  nand2 gate1000(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate1001(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate1002(.a(G570), .O(gate185inter7));
  inv1  gate1003(.a(G571), .O(gate185inter8));
  nand2 gate1004(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate1005(.a(s_65), .b(gate185inter3), .O(gate185inter10));
  nor2  gate1006(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate1007(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate1008(.a(gate185inter12), .b(gate185inter1), .O(G602));

  xor2  gate1765(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1766(.a(gate186inter0), .b(s_174), .O(gate186inter1));
  and2  gate1767(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1768(.a(s_174), .O(gate186inter3));
  inv1  gate1769(.a(s_175), .O(gate186inter4));
  nand2 gate1770(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1771(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1772(.a(G572), .O(gate186inter7));
  inv1  gate1773(.a(G573), .O(gate186inter8));
  nand2 gate1774(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1775(.a(s_175), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1776(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1777(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1778(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate589(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate590(.a(gate190inter0), .b(s_6), .O(gate190inter1));
  and2  gate591(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate592(.a(s_6), .O(gate190inter3));
  inv1  gate593(.a(s_7), .O(gate190inter4));
  nand2 gate594(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate595(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate596(.a(G580), .O(gate190inter7));
  inv1  gate597(.a(G581), .O(gate190inter8));
  nand2 gate598(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate599(.a(s_7), .b(gate190inter3), .O(gate190inter10));
  nor2  gate600(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate601(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate602(.a(gate190inter12), .b(gate190inter1), .O(G627));

  xor2  gate2465(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate2466(.a(gate191inter0), .b(s_274), .O(gate191inter1));
  and2  gate2467(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate2468(.a(s_274), .O(gate191inter3));
  inv1  gate2469(.a(s_275), .O(gate191inter4));
  nand2 gate2470(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate2471(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate2472(.a(G582), .O(gate191inter7));
  inv1  gate2473(.a(G583), .O(gate191inter8));
  nand2 gate2474(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate2475(.a(s_275), .b(gate191inter3), .O(gate191inter10));
  nor2  gate2476(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate2477(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate2478(.a(gate191inter12), .b(gate191inter1), .O(G632));

  xor2  gate883(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate884(.a(gate192inter0), .b(s_48), .O(gate192inter1));
  and2  gate885(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate886(.a(s_48), .O(gate192inter3));
  inv1  gate887(.a(s_49), .O(gate192inter4));
  nand2 gate888(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate889(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate890(.a(G584), .O(gate192inter7));
  inv1  gate891(.a(G585), .O(gate192inter8));
  nand2 gate892(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate893(.a(s_49), .b(gate192inter3), .O(gate192inter10));
  nor2  gate894(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate895(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate896(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate1009(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate1010(.a(gate195inter0), .b(s_66), .O(gate195inter1));
  and2  gate1011(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate1012(.a(s_66), .O(gate195inter3));
  inv1  gate1013(.a(s_67), .O(gate195inter4));
  nand2 gate1014(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate1015(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate1016(.a(G590), .O(gate195inter7));
  inv1  gate1017(.a(G591), .O(gate195inter8));
  nand2 gate1018(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate1019(.a(s_67), .b(gate195inter3), .O(gate195inter10));
  nor2  gate1020(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate1021(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate1022(.a(gate195inter12), .b(gate195inter1), .O(G648));

  xor2  gate2059(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate2060(.a(gate196inter0), .b(s_216), .O(gate196inter1));
  and2  gate2061(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate2062(.a(s_216), .O(gate196inter3));
  inv1  gate2063(.a(s_217), .O(gate196inter4));
  nand2 gate2064(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate2065(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate2066(.a(G592), .O(gate196inter7));
  inv1  gate2067(.a(G593), .O(gate196inter8));
  nand2 gate2068(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate2069(.a(s_217), .b(gate196inter3), .O(gate196inter10));
  nor2  gate2070(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate2071(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate2072(.a(gate196inter12), .b(gate196inter1), .O(G651));

  xor2  gate1205(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate1206(.a(gate197inter0), .b(s_94), .O(gate197inter1));
  and2  gate1207(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate1208(.a(s_94), .O(gate197inter3));
  inv1  gate1209(.a(s_95), .O(gate197inter4));
  nand2 gate1210(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate1211(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate1212(.a(G594), .O(gate197inter7));
  inv1  gate1213(.a(G595), .O(gate197inter8));
  nand2 gate1214(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate1215(.a(s_95), .b(gate197inter3), .O(gate197inter10));
  nor2  gate1216(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate1217(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate1218(.a(gate197inter12), .b(gate197inter1), .O(G654));

  xor2  gate715(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate716(.a(gate198inter0), .b(s_24), .O(gate198inter1));
  and2  gate717(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate718(.a(s_24), .O(gate198inter3));
  inv1  gate719(.a(s_25), .O(gate198inter4));
  nand2 gate720(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate721(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate722(.a(G596), .O(gate198inter7));
  inv1  gate723(.a(G597), .O(gate198inter8));
  nand2 gate724(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate725(.a(s_25), .b(gate198inter3), .O(gate198inter10));
  nor2  gate726(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate727(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate728(.a(gate198inter12), .b(gate198inter1), .O(G657));
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate2213(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate2214(.a(gate203inter0), .b(s_238), .O(gate203inter1));
  and2  gate2215(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate2216(.a(s_238), .O(gate203inter3));
  inv1  gate2217(.a(s_239), .O(gate203inter4));
  nand2 gate2218(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate2219(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate2220(.a(G602), .O(gate203inter7));
  inv1  gate2221(.a(G612), .O(gate203inter8));
  nand2 gate2222(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate2223(.a(s_239), .b(gate203inter3), .O(gate203inter10));
  nor2  gate2224(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate2225(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate2226(.a(gate203inter12), .b(gate203inter1), .O(G672));

  xor2  gate1219(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate1220(.a(gate204inter0), .b(s_96), .O(gate204inter1));
  and2  gate1221(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate1222(.a(s_96), .O(gate204inter3));
  inv1  gate1223(.a(s_97), .O(gate204inter4));
  nand2 gate1224(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate1225(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate1226(.a(G607), .O(gate204inter7));
  inv1  gate1227(.a(G617), .O(gate204inter8));
  nand2 gate1228(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate1229(.a(s_97), .b(gate204inter3), .O(gate204inter10));
  nor2  gate1230(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate1231(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate1232(.a(gate204inter12), .b(gate204inter1), .O(G675));

  xor2  gate1289(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate1290(.a(gate205inter0), .b(s_106), .O(gate205inter1));
  and2  gate1291(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate1292(.a(s_106), .O(gate205inter3));
  inv1  gate1293(.a(s_107), .O(gate205inter4));
  nand2 gate1294(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate1295(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate1296(.a(G622), .O(gate205inter7));
  inv1  gate1297(.a(G627), .O(gate205inter8));
  nand2 gate1298(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate1299(.a(s_107), .b(gate205inter3), .O(gate205inter10));
  nor2  gate1300(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate1301(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate1302(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );

  xor2  gate1303(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate1304(.a(gate209inter0), .b(s_108), .O(gate209inter1));
  and2  gate1305(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate1306(.a(s_108), .O(gate209inter3));
  inv1  gate1307(.a(s_109), .O(gate209inter4));
  nand2 gate1308(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate1309(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate1310(.a(G602), .O(gate209inter7));
  inv1  gate1311(.a(G666), .O(gate209inter8));
  nand2 gate1312(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate1313(.a(s_109), .b(gate209inter3), .O(gate209inter10));
  nor2  gate1314(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate1315(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate1316(.a(gate209inter12), .b(gate209inter1), .O(G690));
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );

  xor2  gate2339(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate2340(.a(gate212inter0), .b(s_256), .O(gate212inter1));
  and2  gate2341(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate2342(.a(s_256), .O(gate212inter3));
  inv1  gate2343(.a(s_257), .O(gate212inter4));
  nand2 gate2344(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate2345(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate2346(.a(G617), .O(gate212inter7));
  inv1  gate2347(.a(G669), .O(gate212inter8));
  nand2 gate2348(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate2349(.a(s_257), .b(gate212inter3), .O(gate212inter10));
  nor2  gate2350(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate2351(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate2352(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate1737(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate1738(.a(gate214inter0), .b(s_170), .O(gate214inter1));
  and2  gate1739(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate1740(.a(s_170), .O(gate214inter3));
  inv1  gate1741(.a(s_171), .O(gate214inter4));
  nand2 gate1742(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate1743(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate1744(.a(G612), .O(gate214inter7));
  inv1  gate1745(.a(G672), .O(gate214inter8));
  nand2 gate1746(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate1747(.a(s_171), .b(gate214inter3), .O(gate214inter10));
  nor2  gate1748(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate1749(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate1750(.a(gate214inter12), .b(gate214inter1), .O(G695));

  xor2  gate1905(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate1906(.a(gate215inter0), .b(s_194), .O(gate215inter1));
  and2  gate1907(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate1908(.a(s_194), .O(gate215inter3));
  inv1  gate1909(.a(s_195), .O(gate215inter4));
  nand2 gate1910(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate1911(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate1912(.a(G607), .O(gate215inter7));
  inv1  gate1913(.a(G675), .O(gate215inter8));
  nand2 gate1914(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate1915(.a(s_195), .b(gate215inter3), .O(gate215inter10));
  nor2  gate1916(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate1917(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate1918(.a(gate215inter12), .b(gate215inter1), .O(G696));

  xor2  gate1527(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate1528(.a(gate216inter0), .b(s_140), .O(gate216inter1));
  and2  gate1529(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate1530(.a(s_140), .O(gate216inter3));
  inv1  gate1531(.a(s_141), .O(gate216inter4));
  nand2 gate1532(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate1533(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate1534(.a(G617), .O(gate216inter7));
  inv1  gate1535(.a(G675), .O(gate216inter8));
  nand2 gate1536(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate1537(.a(s_141), .b(gate216inter3), .O(gate216inter10));
  nor2  gate1538(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate1539(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate1540(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate729(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate730(.a(gate218inter0), .b(s_26), .O(gate218inter1));
  and2  gate731(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate732(.a(s_26), .O(gate218inter3));
  inv1  gate733(.a(s_27), .O(gate218inter4));
  nand2 gate734(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate735(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate736(.a(G627), .O(gate218inter7));
  inv1  gate737(.a(G678), .O(gate218inter8));
  nand2 gate738(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate739(.a(s_27), .b(gate218inter3), .O(gate218inter10));
  nor2  gate740(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate741(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate742(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate1401(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate1402(.a(gate223inter0), .b(s_122), .O(gate223inter1));
  and2  gate1403(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate1404(.a(s_122), .O(gate223inter3));
  inv1  gate1405(.a(s_123), .O(gate223inter4));
  nand2 gate1406(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate1407(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate1408(.a(G627), .O(gate223inter7));
  inv1  gate1409(.a(G687), .O(gate223inter8));
  nand2 gate1410(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate1411(.a(s_123), .b(gate223inter3), .O(gate223inter10));
  nor2  gate1412(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate1413(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate1414(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );

  xor2  gate2017(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate2018(.a(gate225inter0), .b(s_210), .O(gate225inter1));
  and2  gate2019(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate2020(.a(s_210), .O(gate225inter3));
  inv1  gate2021(.a(s_211), .O(gate225inter4));
  nand2 gate2022(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate2023(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate2024(.a(G690), .O(gate225inter7));
  inv1  gate2025(.a(G691), .O(gate225inter8));
  nand2 gate2026(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate2027(.a(s_211), .b(gate225inter3), .O(gate225inter10));
  nor2  gate2028(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate2029(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate2030(.a(gate225inter12), .b(gate225inter1), .O(G706));

  xor2  gate1415(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate1416(.a(gate226inter0), .b(s_124), .O(gate226inter1));
  and2  gate1417(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate1418(.a(s_124), .O(gate226inter3));
  inv1  gate1419(.a(s_125), .O(gate226inter4));
  nand2 gate1420(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate1421(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate1422(.a(G692), .O(gate226inter7));
  inv1  gate1423(.a(G693), .O(gate226inter8));
  nand2 gate1424(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate1425(.a(s_125), .b(gate226inter3), .O(gate226inter10));
  nor2  gate1426(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate1427(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate1428(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate771(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate772(.a(gate228inter0), .b(s_32), .O(gate228inter1));
  and2  gate773(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate774(.a(s_32), .O(gate228inter3));
  inv1  gate775(.a(s_33), .O(gate228inter4));
  nand2 gate776(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate777(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate778(.a(G696), .O(gate228inter7));
  inv1  gate779(.a(G697), .O(gate228inter8));
  nand2 gate780(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate781(.a(s_33), .b(gate228inter3), .O(gate228inter10));
  nor2  gate782(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate783(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate784(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate1373(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate1374(.a(gate231inter0), .b(s_118), .O(gate231inter1));
  and2  gate1375(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate1376(.a(s_118), .O(gate231inter3));
  inv1  gate1377(.a(s_119), .O(gate231inter4));
  nand2 gate1378(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate1379(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate1380(.a(G702), .O(gate231inter7));
  inv1  gate1381(.a(G703), .O(gate231inter8));
  nand2 gate1382(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate1383(.a(s_119), .b(gate231inter3), .O(gate231inter10));
  nor2  gate1384(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate1385(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate1386(.a(gate231inter12), .b(gate231inter1), .O(G724));

  xor2  gate2283(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate2284(.a(gate232inter0), .b(s_248), .O(gate232inter1));
  and2  gate2285(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate2286(.a(s_248), .O(gate232inter3));
  inv1  gate2287(.a(s_249), .O(gate232inter4));
  nand2 gate2288(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate2289(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate2290(.a(G704), .O(gate232inter7));
  inv1  gate2291(.a(G705), .O(gate232inter8));
  nand2 gate2292(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate2293(.a(s_249), .b(gate232inter3), .O(gate232inter10));
  nor2  gate2294(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate2295(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate2296(.a(gate232inter12), .b(gate232inter1), .O(G727));
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate2031(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate2032(.a(gate234inter0), .b(s_212), .O(gate234inter1));
  and2  gate2033(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate2034(.a(s_212), .O(gate234inter3));
  inv1  gate2035(.a(s_213), .O(gate234inter4));
  nand2 gate2036(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate2037(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate2038(.a(G245), .O(gate234inter7));
  inv1  gate2039(.a(G721), .O(gate234inter8));
  nand2 gate2040(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate2041(.a(s_213), .b(gate234inter3), .O(gate234inter10));
  nor2  gate2042(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate2043(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate2044(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );

  xor2  gate1681(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate1682(.a(gate239inter0), .b(s_162), .O(gate239inter1));
  and2  gate1683(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate1684(.a(s_162), .O(gate239inter3));
  inv1  gate1685(.a(s_163), .O(gate239inter4));
  nand2 gate1686(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate1687(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate1688(.a(G260), .O(gate239inter7));
  inv1  gate1689(.a(G712), .O(gate239inter8));
  nand2 gate1690(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate1691(.a(s_163), .b(gate239inter3), .O(gate239inter10));
  nor2  gate1692(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate1693(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate1694(.a(gate239inter12), .b(gate239inter1), .O(G748));
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );

  xor2  gate1975(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate1976(.a(gate244inter0), .b(s_204), .O(gate244inter1));
  and2  gate1977(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate1978(.a(s_204), .O(gate244inter3));
  inv1  gate1979(.a(s_205), .O(gate244inter4));
  nand2 gate1980(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate1981(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate1982(.a(G721), .O(gate244inter7));
  inv1  gate1983(.a(G733), .O(gate244inter8));
  nand2 gate1984(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate1985(.a(s_205), .b(gate244inter3), .O(gate244inter10));
  nor2  gate1986(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate1987(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate1988(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate1751(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate1752(.a(gate248inter0), .b(s_172), .O(gate248inter1));
  and2  gate1753(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate1754(.a(s_172), .O(gate248inter3));
  inv1  gate1755(.a(s_173), .O(gate248inter4));
  nand2 gate1756(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate1757(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate1758(.a(G727), .O(gate248inter7));
  inv1  gate1759(.a(G739), .O(gate248inter8));
  nand2 gate1760(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate1761(.a(s_173), .b(gate248inter3), .O(gate248inter10));
  nor2  gate1762(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate1763(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate1764(.a(gate248inter12), .b(gate248inter1), .O(G761));

  xor2  gate2087(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate2088(.a(gate249inter0), .b(s_220), .O(gate249inter1));
  and2  gate2089(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate2090(.a(s_220), .O(gate249inter3));
  inv1  gate2091(.a(s_221), .O(gate249inter4));
  nand2 gate2092(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate2093(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate2094(.a(G254), .O(gate249inter7));
  inv1  gate2095(.a(G742), .O(gate249inter8));
  nand2 gate2096(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate2097(.a(s_221), .b(gate249inter3), .O(gate249inter10));
  nor2  gate2098(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate2099(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate2100(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );

  xor2  gate687(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate688(.a(gate254inter0), .b(s_20), .O(gate254inter1));
  and2  gate689(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate690(.a(s_20), .O(gate254inter3));
  inv1  gate691(.a(s_21), .O(gate254inter4));
  nand2 gate692(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate693(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate694(.a(G712), .O(gate254inter7));
  inv1  gate695(.a(G748), .O(gate254inter8));
  nand2 gate696(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate697(.a(s_21), .b(gate254inter3), .O(gate254inter10));
  nor2  gate698(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate699(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate700(.a(gate254inter12), .b(gate254inter1), .O(G767));
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate1863(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate1864(.a(gate256inter0), .b(s_188), .O(gate256inter1));
  and2  gate1865(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate1866(.a(s_188), .O(gate256inter3));
  inv1  gate1867(.a(s_189), .O(gate256inter4));
  nand2 gate1868(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate1869(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate1870(.a(G715), .O(gate256inter7));
  inv1  gate1871(.a(G751), .O(gate256inter8));
  nand2 gate1872(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate1873(.a(s_189), .b(gate256inter3), .O(gate256inter10));
  nor2  gate1874(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate1875(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate1876(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate2325(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate2326(.a(gate258inter0), .b(s_254), .O(gate258inter1));
  and2  gate2327(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate2328(.a(s_254), .O(gate258inter3));
  inv1  gate2329(.a(s_255), .O(gate258inter4));
  nand2 gate2330(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate2331(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate2332(.a(G756), .O(gate258inter7));
  inv1  gate2333(.a(G757), .O(gate258inter8));
  nand2 gate2334(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate2335(.a(s_255), .b(gate258inter3), .O(gate258inter10));
  nor2  gate2336(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate2337(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate2338(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );

  xor2  gate1947(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate1948(.a(gate264inter0), .b(s_200), .O(gate264inter1));
  and2  gate1949(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate1950(.a(s_200), .O(gate264inter3));
  inv1  gate1951(.a(s_201), .O(gate264inter4));
  nand2 gate1952(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate1953(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate1954(.a(G768), .O(gate264inter7));
  inv1  gate1955(.a(G769), .O(gate264inter8));
  nand2 gate1956(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate1957(.a(s_201), .b(gate264inter3), .O(gate264inter10));
  nor2  gate1958(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate1959(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate1960(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate1541(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate1542(.a(gate269inter0), .b(s_142), .O(gate269inter1));
  and2  gate1543(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate1544(.a(s_142), .O(gate269inter3));
  inv1  gate1545(.a(s_143), .O(gate269inter4));
  nand2 gate1546(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate1547(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate1548(.a(G654), .O(gate269inter7));
  inv1  gate1549(.a(G782), .O(gate269inter8));
  nand2 gate1550(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate1551(.a(s_143), .b(gate269inter3), .O(gate269inter10));
  nor2  gate1552(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate1553(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate1554(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );

  xor2  gate869(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate870(.a(gate275inter0), .b(s_46), .O(gate275inter1));
  and2  gate871(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate872(.a(s_46), .O(gate275inter3));
  inv1  gate873(.a(s_47), .O(gate275inter4));
  nand2 gate874(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate875(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate876(.a(G645), .O(gate275inter7));
  inv1  gate877(.a(G797), .O(gate275inter8));
  nand2 gate878(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate879(.a(s_47), .b(gate275inter3), .O(gate275inter10));
  nor2  gate880(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate881(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate882(.a(gate275inter12), .b(gate275inter1), .O(G820));

  xor2  gate1611(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate1612(.a(gate276inter0), .b(s_152), .O(gate276inter1));
  and2  gate1613(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate1614(.a(s_152), .O(gate276inter3));
  inv1  gate1615(.a(s_153), .O(gate276inter4));
  nand2 gate1616(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate1617(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate1618(.a(G773), .O(gate276inter7));
  inv1  gate1619(.a(G797), .O(gate276inter8));
  nand2 gate1620(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate1621(.a(s_153), .b(gate276inter3), .O(gate276inter10));
  nor2  gate1622(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate1623(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate1624(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate673(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate674(.a(gate279inter0), .b(s_18), .O(gate279inter1));
  and2  gate675(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate676(.a(s_18), .O(gate279inter3));
  inv1  gate677(.a(s_19), .O(gate279inter4));
  nand2 gate678(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate679(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate680(.a(G651), .O(gate279inter7));
  inv1  gate681(.a(G803), .O(gate279inter8));
  nand2 gate682(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate683(.a(s_19), .b(gate279inter3), .O(gate279inter10));
  nor2  gate684(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate685(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate686(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate1261(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate1262(.a(gate283inter0), .b(s_102), .O(gate283inter1));
  and2  gate1263(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate1264(.a(s_102), .O(gate283inter3));
  inv1  gate1265(.a(s_103), .O(gate283inter4));
  nand2 gate1266(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate1267(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate1268(.a(G657), .O(gate283inter7));
  inv1  gate1269(.a(G809), .O(gate283inter8));
  nand2 gate1270(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate1271(.a(s_103), .b(gate283inter3), .O(gate283inter10));
  nor2  gate1272(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate1273(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate1274(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate2437(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate2438(.a(gate286inter0), .b(s_270), .O(gate286inter1));
  and2  gate2439(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate2440(.a(s_270), .O(gate286inter3));
  inv1  gate2441(.a(s_271), .O(gate286inter4));
  nand2 gate2442(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate2443(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate2444(.a(G788), .O(gate286inter7));
  inv1  gate2445(.a(G812), .O(gate286inter8));
  nand2 gate2446(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate2447(.a(s_271), .b(gate286inter3), .O(gate286inter10));
  nor2  gate2448(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate2449(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate2450(.a(gate286inter12), .b(gate286inter1), .O(G831));

  xor2  gate841(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate842(.a(gate287inter0), .b(s_42), .O(gate287inter1));
  and2  gate843(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate844(.a(s_42), .O(gate287inter3));
  inv1  gate845(.a(s_43), .O(gate287inter4));
  nand2 gate846(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate847(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate848(.a(G663), .O(gate287inter7));
  inv1  gate849(.a(G815), .O(gate287inter8));
  nand2 gate850(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate851(.a(s_43), .b(gate287inter3), .O(gate287inter10));
  nor2  gate852(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate853(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate854(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate1877(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate1878(.a(gate293inter0), .b(s_190), .O(gate293inter1));
  and2  gate1879(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate1880(.a(s_190), .O(gate293inter3));
  inv1  gate1881(.a(s_191), .O(gate293inter4));
  nand2 gate1882(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate1883(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate1884(.a(G828), .O(gate293inter7));
  inv1  gate1885(.a(G829), .O(gate293inter8));
  nand2 gate1886(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate1887(.a(s_191), .b(gate293inter3), .O(gate293inter10));
  nor2  gate1888(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate1889(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate1890(.a(gate293inter12), .b(gate293inter1), .O(G886));

  xor2  gate1233(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate1234(.a(gate294inter0), .b(s_98), .O(gate294inter1));
  and2  gate1235(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate1236(.a(s_98), .O(gate294inter3));
  inv1  gate1237(.a(s_99), .O(gate294inter4));
  nand2 gate1238(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate1239(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate1240(.a(G832), .O(gate294inter7));
  inv1  gate1241(.a(G833), .O(gate294inter8));
  nand2 gate1242(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate1243(.a(s_99), .b(gate294inter3), .O(gate294inter10));
  nor2  gate1244(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate1245(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate1246(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate1275(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate1276(.a(gate387inter0), .b(s_104), .O(gate387inter1));
  and2  gate1277(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate1278(.a(s_104), .O(gate387inter3));
  inv1  gate1279(.a(s_105), .O(gate387inter4));
  nand2 gate1280(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1281(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1282(.a(G1), .O(gate387inter7));
  inv1  gate1283(.a(G1036), .O(gate387inter8));
  nand2 gate1284(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1285(.a(s_105), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1286(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1287(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate1288(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate1023(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate1024(.a(gate390inter0), .b(s_68), .O(gate390inter1));
  and2  gate1025(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate1026(.a(s_68), .O(gate390inter3));
  inv1  gate1027(.a(s_69), .O(gate390inter4));
  nand2 gate1028(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate1029(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate1030(.a(G4), .O(gate390inter7));
  inv1  gate1031(.a(G1045), .O(gate390inter8));
  nand2 gate1032(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate1033(.a(s_69), .b(gate390inter3), .O(gate390inter10));
  nor2  gate1034(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate1035(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate1036(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );

  xor2  gate2423(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate2424(.a(gate392inter0), .b(s_268), .O(gate392inter1));
  and2  gate2425(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate2426(.a(s_268), .O(gate392inter3));
  inv1  gate2427(.a(s_269), .O(gate392inter4));
  nand2 gate2428(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate2429(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate2430(.a(G6), .O(gate392inter7));
  inv1  gate2431(.a(G1051), .O(gate392inter8));
  nand2 gate2432(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate2433(.a(s_269), .b(gate392inter3), .O(gate392inter10));
  nor2  gate2434(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate2435(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate2436(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate1247(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1248(.a(gate395inter0), .b(s_100), .O(gate395inter1));
  and2  gate1249(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1250(.a(s_100), .O(gate395inter3));
  inv1  gate1251(.a(s_101), .O(gate395inter4));
  nand2 gate1252(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1253(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1254(.a(G9), .O(gate395inter7));
  inv1  gate1255(.a(G1060), .O(gate395inter8));
  nand2 gate1256(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1257(.a(s_101), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1258(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1259(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1260(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );

  xor2  gate659(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate660(.a(gate401inter0), .b(s_16), .O(gate401inter1));
  and2  gate661(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate662(.a(s_16), .O(gate401inter3));
  inv1  gate663(.a(s_17), .O(gate401inter4));
  nand2 gate664(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate665(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate666(.a(G15), .O(gate401inter7));
  inv1  gate667(.a(G1078), .O(gate401inter8));
  nand2 gate668(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate669(.a(s_17), .b(gate401inter3), .O(gate401inter10));
  nor2  gate670(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate671(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate672(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate1639(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate1640(.a(gate403inter0), .b(s_156), .O(gate403inter1));
  and2  gate1641(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate1642(.a(s_156), .O(gate403inter3));
  inv1  gate1643(.a(s_157), .O(gate403inter4));
  nand2 gate1644(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate1645(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate1646(.a(G17), .O(gate403inter7));
  inv1  gate1647(.a(G1084), .O(gate403inter8));
  nand2 gate1648(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate1649(.a(s_157), .b(gate403inter3), .O(gate403inter10));
  nor2  gate1650(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate1651(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate1652(.a(gate403inter12), .b(gate403inter1), .O(G1180));
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );

  xor2  gate1191(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate1192(.a(gate405inter0), .b(s_92), .O(gate405inter1));
  and2  gate1193(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate1194(.a(s_92), .O(gate405inter3));
  inv1  gate1195(.a(s_93), .O(gate405inter4));
  nand2 gate1196(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate1197(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate1198(.a(G19), .O(gate405inter7));
  inv1  gate1199(.a(G1090), .O(gate405inter8));
  nand2 gate1200(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate1201(.a(s_93), .b(gate405inter3), .O(gate405inter10));
  nor2  gate1202(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate1203(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate1204(.a(gate405inter12), .b(gate405inter1), .O(G1186));

  xor2  gate799(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate800(.a(gate406inter0), .b(s_36), .O(gate406inter1));
  and2  gate801(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate802(.a(s_36), .O(gate406inter3));
  inv1  gate803(.a(s_37), .O(gate406inter4));
  nand2 gate804(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate805(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate806(.a(G20), .O(gate406inter7));
  inv1  gate807(.a(G1093), .O(gate406inter8));
  nand2 gate808(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate809(.a(s_37), .b(gate406inter3), .O(gate406inter10));
  nor2  gate810(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate811(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate812(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate1569(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate1570(.a(gate410inter0), .b(s_146), .O(gate410inter1));
  and2  gate1571(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate1572(.a(s_146), .O(gate410inter3));
  inv1  gate1573(.a(s_147), .O(gate410inter4));
  nand2 gate1574(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate1575(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate1576(.a(G24), .O(gate410inter7));
  inv1  gate1577(.a(G1105), .O(gate410inter8));
  nand2 gate1578(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate1579(.a(s_147), .b(gate410inter3), .O(gate410inter10));
  nor2  gate1580(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate1581(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate1582(.a(gate410inter12), .b(gate410inter1), .O(G1201));

  xor2  gate645(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate646(.a(gate411inter0), .b(s_14), .O(gate411inter1));
  and2  gate647(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate648(.a(s_14), .O(gate411inter3));
  inv1  gate649(.a(s_15), .O(gate411inter4));
  nand2 gate650(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate651(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate652(.a(G25), .O(gate411inter7));
  inv1  gate653(.a(G1108), .O(gate411inter8));
  nand2 gate654(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate655(.a(s_15), .b(gate411inter3), .O(gate411inter10));
  nor2  gate656(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate657(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate658(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate967(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate968(.a(gate415inter0), .b(s_60), .O(gate415inter1));
  and2  gate969(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate970(.a(s_60), .O(gate415inter3));
  inv1  gate971(.a(s_61), .O(gate415inter4));
  nand2 gate972(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate973(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate974(.a(G29), .O(gate415inter7));
  inv1  gate975(.a(G1120), .O(gate415inter8));
  nand2 gate976(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate977(.a(s_61), .b(gate415inter3), .O(gate415inter10));
  nor2  gate978(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate979(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate980(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate2297(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate2298(.a(gate417inter0), .b(s_250), .O(gate417inter1));
  and2  gate2299(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate2300(.a(s_250), .O(gate417inter3));
  inv1  gate2301(.a(s_251), .O(gate417inter4));
  nand2 gate2302(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate2303(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate2304(.a(G31), .O(gate417inter7));
  inv1  gate2305(.a(G1126), .O(gate417inter8));
  nand2 gate2306(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate2307(.a(s_251), .b(gate417inter3), .O(gate417inter10));
  nor2  gate2308(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate2309(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate2310(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate1961(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate1962(.a(gate425inter0), .b(s_202), .O(gate425inter1));
  and2  gate1963(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate1964(.a(s_202), .O(gate425inter3));
  inv1  gate1965(.a(s_203), .O(gate425inter4));
  nand2 gate1966(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1967(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1968(.a(G4), .O(gate425inter7));
  inv1  gate1969(.a(G1141), .O(gate425inter8));
  nand2 gate1970(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1971(.a(s_203), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1972(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1973(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1974(.a(gate425inter12), .b(gate425inter1), .O(G1234));
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );

  xor2  gate1513(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate1514(.a(gate429inter0), .b(s_138), .O(gate429inter1));
  and2  gate1515(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate1516(.a(s_138), .O(gate429inter3));
  inv1  gate1517(.a(s_139), .O(gate429inter4));
  nand2 gate1518(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate1519(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate1520(.a(G6), .O(gate429inter7));
  inv1  gate1521(.a(G1147), .O(gate429inter8));
  nand2 gate1522(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate1523(.a(s_139), .b(gate429inter3), .O(gate429inter10));
  nor2  gate1524(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate1525(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate1526(.a(gate429inter12), .b(gate429inter1), .O(G1238));

  xor2  gate1695(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate1696(.a(gate430inter0), .b(s_164), .O(gate430inter1));
  and2  gate1697(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate1698(.a(s_164), .O(gate430inter3));
  inv1  gate1699(.a(s_165), .O(gate430inter4));
  nand2 gate1700(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate1701(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate1702(.a(G1051), .O(gate430inter7));
  inv1  gate1703(.a(G1147), .O(gate430inter8));
  nand2 gate1704(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate1705(.a(s_165), .b(gate430inter3), .O(gate430inter10));
  nor2  gate1706(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate1707(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate1708(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate953(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate954(.a(gate433inter0), .b(s_58), .O(gate433inter1));
  and2  gate955(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate956(.a(s_58), .O(gate433inter3));
  inv1  gate957(.a(s_59), .O(gate433inter4));
  nand2 gate958(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate959(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate960(.a(G8), .O(gate433inter7));
  inv1  gate961(.a(G1153), .O(gate433inter8));
  nand2 gate962(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate963(.a(s_59), .b(gate433inter3), .O(gate433inter10));
  nor2  gate964(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate965(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate966(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate1359(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate1360(.a(gate435inter0), .b(s_116), .O(gate435inter1));
  and2  gate1361(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate1362(.a(s_116), .O(gate435inter3));
  inv1  gate1363(.a(s_117), .O(gate435inter4));
  nand2 gate1364(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate1365(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate1366(.a(G9), .O(gate435inter7));
  inv1  gate1367(.a(G1156), .O(gate435inter8));
  nand2 gate1368(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate1369(.a(s_117), .b(gate435inter3), .O(gate435inter10));
  nor2  gate1370(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate1371(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate1372(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate1709(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate1710(.a(gate438inter0), .b(s_166), .O(gate438inter1));
  and2  gate1711(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate1712(.a(s_166), .O(gate438inter3));
  inv1  gate1713(.a(s_167), .O(gate438inter4));
  nand2 gate1714(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate1715(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate1716(.a(G1063), .O(gate438inter7));
  inv1  gate1717(.a(G1159), .O(gate438inter8));
  nand2 gate1718(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate1719(.a(s_167), .b(gate438inter3), .O(gate438inter10));
  nor2  gate1720(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate1721(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate1722(.a(gate438inter12), .b(gate438inter1), .O(G1247));

  xor2  gate925(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate926(.a(gate439inter0), .b(s_54), .O(gate439inter1));
  and2  gate927(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate928(.a(s_54), .O(gate439inter3));
  inv1  gate929(.a(s_55), .O(gate439inter4));
  nand2 gate930(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate931(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate932(.a(G11), .O(gate439inter7));
  inv1  gate933(.a(G1162), .O(gate439inter8));
  nand2 gate934(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate935(.a(s_55), .b(gate439inter3), .O(gate439inter10));
  nor2  gate936(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate937(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate938(.a(gate439inter12), .b(gate439inter1), .O(G1248));

  xor2  gate701(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate702(.a(gate440inter0), .b(s_22), .O(gate440inter1));
  and2  gate703(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate704(.a(s_22), .O(gate440inter3));
  inv1  gate705(.a(s_23), .O(gate440inter4));
  nand2 gate706(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate707(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate708(.a(G1066), .O(gate440inter7));
  inv1  gate709(.a(G1162), .O(gate440inter8));
  nand2 gate710(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate711(.a(s_23), .b(gate440inter3), .O(gate440inter10));
  nor2  gate712(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate713(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate714(.a(gate440inter12), .b(gate440inter1), .O(G1249));

  xor2  gate1835(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate1836(.a(gate441inter0), .b(s_184), .O(gate441inter1));
  and2  gate1837(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate1838(.a(s_184), .O(gate441inter3));
  inv1  gate1839(.a(s_185), .O(gate441inter4));
  nand2 gate1840(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate1841(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate1842(.a(G12), .O(gate441inter7));
  inv1  gate1843(.a(G1165), .O(gate441inter8));
  nand2 gate1844(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate1845(.a(s_185), .b(gate441inter3), .O(gate441inter10));
  nor2  gate1846(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate1847(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate1848(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate1457(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate1458(.a(gate443inter0), .b(s_130), .O(gate443inter1));
  and2  gate1459(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate1460(.a(s_130), .O(gate443inter3));
  inv1  gate1461(.a(s_131), .O(gate443inter4));
  nand2 gate1462(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate1463(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate1464(.a(G13), .O(gate443inter7));
  inv1  gate1465(.a(G1168), .O(gate443inter8));
  nand2 gate1466(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate1467(.a(s_131), .b(gate443inter3), .O(gate443inter10));
  nor2  gate1468(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate1469(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate1470(.a(gate443inter12), .b(gate443inter1), .O(G1252));

  xor2  gate561(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate562(.a(gate444inter0), .b(s_2), .O(gate444inter1));
  and2  gate563(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate564(.a(s_2), .O(gate444inter3));
  inv1  gate565(.a(s_3), .O(gate444inter4));
  nand2 gate566(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate567(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate568(.a(G1072), .O(gate444inter7));
  inv1  gate569(.a(G1168), .O(gate444inter8));
  nand2 gate570(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate571(.a(s_3), .b(gate444inter3), .O(gate444inter10));
  nor2  gate572(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate573(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate574(.a(gate444inter12), .b(gate444inter1), .O(G1253));

  xor2  gate1163(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate1164(.a(gate445inter0), .b(s_88), .O(gate445inter1));
  and2  gate1165(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate1166(.a(s_88), .O(gate445inter3));
  inv1  gate1167(.a(s_89), .O(gate445inter4));
  nand2 gate1168(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate1169(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate1170(.a(G14), .O(gate445inter7));
  inv1  gate1171(.a(G1171), .O(gate445inter8));
  nand2 gate1172(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate1173(.a(s_89), .b(gate445inter3), .O(gate445inter10));
  nor2  gate1174(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate1175(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate1176(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate1989(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate1990(.a(gate448inter0), .b(s_206), .O(gate448inter1));
  and2  gate1991(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate1992(.a(s_206), .O(gate448inter3));
  inv1  gate1993(.a(s_207), .O(gate448inter4));
  nand2 gate1994(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate1995(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate1996(.a(G1078), .O(gate448inter7));
  inv1  gate1997(.a(G1174), .O(gate448inter8));
  nand2 gate1998(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate1999(.a(s_207), .b(gate448inter3), .O(gate448inter10));
  nor2  gate2000(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate2001(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate2002(.a(gate448inter12), .b(gate448inter1), .O(G1257));
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );

  xor2  gate2073(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate2074(.a(gate450inter0), .b(s_218), .O(gate450inter1));
  and2  gate2075(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate2076(.a(s_218), .O(gate450inter3));
  inv1  gate2077(.a(s_219), .O(gate450inter4));
  nand2 gate2078(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate2079(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate2080(.a(G1081), .O(gate450inter7));
  inv1  gate2081(.a(G1177), .O(gate450inter8));
  nand2 gate2082(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate2083(.a(s_219), .b(gate450inter3), .O(gate450inter10));
  nor2  gate2084(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate2085(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate2086(.a(gate450inter12), .b(gate450inter1), .O(G1259));

  xor2  gate1625(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate1626(.a(gate451inter0), .b(s_154), .O(gate451inter1));
  and2  gate1627(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate1628(.a(s_154), .O(gate451inter3));
  inv1  gate1629(.a(s_155), .O(gate451inter4));
  nand2 gate1630(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate1631(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate1632(.a(G17), .O(gate451inter7));
  inv1  gate1633(.a(G1180), .O(gate451inter8));
  nand2 gate1634(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate1635(.a(s_155), .b(gate451inter3), .O(gate451inter10));
  nor2  gate1636(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate1637(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate1638(.a(gate451inter12), .b(gate451inter1), .O(G1260));

  xor2  gate1387(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate1388(.a(gate452inter0), .b(s_120), .O(gate452inter1));
  and2  gate1389(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate1390(.a(s_120), .O(gate452inter3));
  inv1  gate1391(.a(s_121), .O(gate452inter4));
  nand2 gate1392(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate1393(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate1394(.a(G1084), .O(gate452inter7));
  inv1  gate1395(.a(G1180), .O(gate452inter8));
  nand2 gate1396(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate1397(.a(s_121), .b(gate452inter3), .O(gate452inter10));
  nor2  gate1398(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate1399(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate1400(.a(gate452inter12), .b(gate452inter1), .O(G1261));

  xor2  gate631(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate632(.a(gate453inter0), .b(s_12), .O(gate453inter1));
  and2  gate633(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate634(.a(s_12), .O(gate453inter3));
  inv1  gate635(.a(s_13), .O(gate453inter4));
  nand2 gate636(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate637(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate638(.a(G18), .O(gate453inter7));
  inv1  gate639(.a(G1183), .O(gate453inter8));
  nand2 gate640(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate641(.a(s_13), .b(gate453inter3), .O(gate453inter10));
  nor2  gate642(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate643(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate644(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );

  xor2  gate1429(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate1430(.a(gate455inter0), .b(s_126), .O(gate455inter1));
  and2  gate1431(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate1432(.a(s_126), .O(gate455inter3));
  inv1  gate1433(.a(s_127), .O(gate455inter4));
  nand2 gate1434(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate1435(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate1436(.a(G19), .O(gate455inter7));
  inv1  gate1437(.a(G1186), .O(gate455inter8));
  nand2 gate1438(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate1439(.a(s_127), .b(gate455inter3), .O(gate455inter10));
  nor2  gate1440(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate1441(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate1442(.a(gate455inter12), .b(gate455inter1), .O(G1264));

  xor2  gate1177(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate1178(.a(gate456inter0), .b(s_90), .O(gate456inter1));
  and2  gate1179(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate1180(.a(s_90), .O(gate456inter3));
  inv1  gate1181(.a(s_91), .O(gate456inter4));
  nand2 gate1182(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate1183(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate1184(.a(G1090), .O(gate456inter7));
  inv1  gate1185(.a(G1186), .O(gate456inter8));
  nand2 gate1186(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate1187(.a(s_91), .b(gate456inter3), .O(gate456inter10));
  nor2  gate1188(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate1189(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate1190(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );

  xor2  gate547(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate548(.a(gate458inter0), .b(s_0), .O(gate458inter1));
  and2  gate549(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate550(.a(s_0), .O(gate458inter3));
  inv1  gate551(.a(s_1), .O(gate458inter4));
  nand2 gate552(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate553(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate554(.a(G1093), .O(gate458inter7));
  inv1  gate555(.a(G1189), .O(gate458inter8));
  nand2 gate556(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate557(.a(s_1), .b(gate458inter3), .O(gate458inter10));
  nor2  gate558(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate559(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate560(.a(gate458inter12), .b(gate458inter1), .O(G1267));
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate1149(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate1150(.a(gate461inter0), .b(s_86), .O(gate461inter1));
  and2  gate1151(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate1152(.a(s_86), .O(gate461inter3));
  inv1  gate1153(.a(s_87), .O(gate461inter4));
  nand2 gate1154(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate1155(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate1156(.a(G22), .O(gate461inter7));
  inv1  gate1157(.a(G1195), .O(gate461inter8));
  nand2 gate1158(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate1159(.a(s_87), .b(gate461inter3), .O(gate461inter10));
  nor2  gate1160(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate1161(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate1162(.a(gate461inter12), .b(gate461inter1), .O(G1270));

  xor2  gate2451(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate2452(.a(gate462inter0), .b(s_272), .O(gate462inter1));
  and2  gate2453(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate2454(.a(s_272), .O(gate462inter3));
  inv1  gate2455(.a(s_273), .O(gate462inter4));
  nand2 gate2456(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate2457(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate2458(.a(G1099), .O(gate462inter7));
  inv1  gate2459(.a(G1195), .O(gate462inter8));
  nand2 gate2460(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate2461(.a(s_273), .b(gate462inter3), .O(gate462inter10));
  nor2  gate2462(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate2463(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate2464(.a(gate462inter12), .b(gate462inter1), .O(G1271));
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate1779(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate1780(.a(gate464inter0), .b(s_176), .O(gate464inter1));
  and2  gate1781(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate1782(.a(s_176), .O(gate464inter3));
  inv1  gate1783(.a(s_177), .O(gate464inter4));
  nand2 gate1784(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate1785(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate1786(.a(G1102), .O(gate464inter7));
  inv1  gate1787(.a(G1198), .O(gate464inter8));
  nand2 gate1788(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate1789(.a(s_177), .b(gate464inter3), .O(gate464inter10));
  nor2  gate1790(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate1791(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate1792(.a(gate464inter12), .b(gate464inter1), .O(G1273));

  xor2  gate2185(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate2186(.a(gate465inter0), .b(s_234), .O(gate465inter1));
  and2  gate2187(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate2188(.a(s_234), .O(gate465inter3));
  inv1  gate2189(.a(s_235), .O(gate465inter4));
  nand2 gate2190(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate2191(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate2192(.a(G24), .O(gate465inter7));
  inv1  gate2193(.a(G1201), .O(gate465inter8));
  nand2 gate2194(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate2195(.a(s_235), .b(gate465inter3), .O(gate465inter10));
  nor2  gate2196(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate2197(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate2198(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate2479(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate2480(.a(gate467inter0), .b(s_276), .O(gate467inter1));
  and2  gate2481(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate2482(.a(s_276), .O(gate467inter3));
  inv1  gate2483(.a(s_277), .O(gate467inter4));
  nand2 gate2484(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate2485(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate2486(.a(G25), .O(gate467inter7));
  inv1  gate2487(.a(G1204), .O(gate467inter8));
  nand2 gate2488(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate2489(.a(s_277), .b(gate467inter3), .O(gate467inter10));
  nor2  gate2490(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate2491(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate2492(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );

  xor2  gate1849(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate1850(.a(gate470inter0), .b(s_186), .O(gate470inter1));
  and2  gate1851(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate1852(.a(s_186), .O(gate470inter3));
  inv1  gate1853(.a(s_187), .O(gate470inter4));
  nand2 gate1854(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate1855(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate1856(.a(G1111), .O(gate470inter7));
  inv1  gate1857(.a(G1207), .O(gate470inter8));
  nand2 gate1858(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate1859(.a(s_187), .b(gate470inter3), .O(gate470inter10));
  nor2  gate1860(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate1861(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate1862(.a(gate470inter12), .b(gate470inter1), .O(G1279));
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate2507(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate2508(.a(gate474inter0), .b(s_280), .O(gate474inter1));
  and2  gate2509(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate2510(.a(s_280), .O(gate474inter3));
  inv1  gate2511(.a(s_281), .O(gate474inter4));
  nand2 gate2512(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate2513(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate2514(.a(G1117), .O(gate474inter7));
  inv1  gate2515(.a(G1213), .O(gate474inter8));
  nand2 gate2516(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate2517(.a(s_281), .b(gate474inter3), .O(gate474inter10));
  nor2  gate2518(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate2519(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate2520(.a(gate474inter12), .b(gate474inter1), .O(G1283));
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate2255(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate2256(.a(gate480inter0), .b(s_244), .O(gate480inter1));
  and2  gate2257(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate2258(.a(s_244), .O(gate480inter3));
  inv1  gate2259(.a(s_245), .O(gate480inter4));
  nand2 gate2260(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate2261(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate2262(.a(G1126), .O(gate480inter7));
  inv1  gate2263(.a(G1222), .O(gate480inter8));
  nand2 gate2264(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate2265(.a(s_245), .b(gate480inter3), .O(gate480inter10));
  nor2  gate2266(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate2267(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate2268(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate855(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate856(.a(gate485inter0), .b(s_44), .O(gate485inter1));
  and2  gate857(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate858(.a(s_44), .O(gate485inter3));
  inv1  gate859(.a(s_45), .O(gate485inter4));
  nand2 gate860(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate861(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate862(.a(G1232), .O(gate485inter7));
  inv1  gate863(.a(G1233), .O(gate485inter8));
  nand2 gate864(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate865(.a(s_45), .b(gate485inter3), .O(gate485inter10));
  nor2  gate866(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate867(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate868(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate1065(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate1066(.a(gate488inter0), .b(s_74), .O(gate488inter1));
  and2  gate1067(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate1068(.a(s_74), .O(gate488inter3));
  inv1  gate1069(.a(s_75), .O(gate488inter4));
  nand2 gate1070(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate1071(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate1072(.a(G1238), .O(gate488inter7));
  inv1  gate1073(.a(G1239), .O(gate488inter8));
  nand2 gate1074(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate1075(.a(s_75), .b(gate488inter3), .O(gate488inter10));
  nor2  gate1076(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate1077(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate1078(.a(gate488inter12), .b(gate488inter1), .O(G1297));

  xor2  gate1079(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate1080(.a(gate489inter0), .b(s_76), .O(gate489inter1));
  and2  gate1081(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate1082(.a(s_76), .O(gate489inter3));
  inv1  gate1083(.a(s_77), .O(gate489inter4));
  nand2 gate1084(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate1085(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate1086(.a(G1240), .O(gate489inter7));
  inv1  gate1087(.a(G1241), .O(gate489inter8));
  nand2 gate1088(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate1089(.a(s_77), .b(gate489inter3), .O(gate489inter10));
  nor2  gate1090(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate1091(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate1092(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate2381(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate2382(.a(gate491inter0), .b(s_262), .O(gate491inter1));
  and2  gate2383(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate2384(.a(s_262), .O(gate491inter3));
  inv1  gate2385(.a(s_263), .O(gate491inter4));
  nand2 gate2386(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate2387(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate2388(.a(G1244), .O(gate491inter7));
  inv1  gate2389(.a(G1245), .O(gate491inter8));
  nand2 gate2390(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate2391(.a(s_263), .b(gate491inter3), .O(gate491inter10));
  nor2  gate2392(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate2393(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate2394(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );

  xor2  gate2143(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate2144(.a(gate495inter0), .b(s_228), .O(gate495inter1));
  and2  gate2145(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate2146(.a(s_228), .O(gate495inter3));
  inv1  gate2147(.a(s_229), .O(gate495inter4));
  nand2 gate2148(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate2149(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate2150(.a(G1252), .O(gate495inter7));
  inv1  gate2151(.a(G1253), .O(gate495inter8));
  nand2 gate2152(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate2153(.a(s_229), .b(gate495inter3), .O(gate495inter10));
  nor2  gate2154(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate2155(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate2156(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );

  xor2  gate2045(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate2046(.a(gate498inter0), .b(s_214), .O(gate498inter1));
  and2  gate2047(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate2048(.a(s_214), .O(gate498inter3));
  inv1  gate2049(.a(s_215), .O(gate498inter4));
  nand2 gate2050(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate2051(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate2052(.a(G1258), .O(gate498inter7));
  inv1  gate2053(.a(G1259), .O(gate498inter8));
  nand2 gate2054(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate2055(.a(s_215), .b(gate498inter3), .O(gate498inter10));
  nor2  gate2056(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate2057(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate2058(.a(gate498inter12), .b(gate498inter1), .O(G1307));
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );

  xor2  gate1093(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate1094(.a(gate507inter0), .b(s_78), .O(gate507inter1));
  and2  gate1095(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate1096(.a(s_78), .O(gate507inter3));
  inv1  gate1097(.a(s_79), .O(gate507inter4));
  nand2 gate1098(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate1099(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate1100(.a(G1276), .O(gate507inter7));
  inv1  gate1101(.a(G1277), .O(gate507inter8));
  nand2 gate1102(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate1103(.a(s_79), .b(gate507inter3), .O(gate507inter10));
  nor2  gate1104(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate1105(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate1106(.a(gate507inter12), .b(gate507inter1), .O(G1316));
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate1793(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate1794(.a(gate510inter0), .b(s_178), .O(gate510inter1));
  and2  gate1795(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate1796(.a(s_178), .O(gate510inter3));
  inv1  gate1797(.a(s_179), .O(gate510inter4));
  nand2 gate1798(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate1799(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate1800(.a(G1282), .O(gate510inter7));
  inv1  gate1801(.a(G1283), .O(gate510inter8));
  nand2 gate1802(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate1803(.a(s_179), .b(gate510inter3), .O(gate510inter10));
  nor2  gate1804(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate1805(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate1806(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule