module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate1205(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate1206(.a(gate20inter0), .b(s_94), .O(gate20inter1));
  and2  gate1207(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate1208(.a(s_94), .O(gate20inter3));
  inv1  gate1209(.a(s_95), .O(gate20inter4));
  nand2 gate1210(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate1211(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate1212(.a(G23), .O(gate20inter7));
  inv1  gate1213(.a(G24), .O(gate20inter8));
  nand2 gate1214(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate1215(.a(s_95), .b(gate20inter3), .O(gate20inter10));
  nor2  gate1216(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate1217(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate1218(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate1121(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate1122(.a(gate22inter0), .b(s_82), .O(gate22inter1));
  and2  gate1123(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate1124(.a(s_82), .O(gate22inter3));
  inv1  gate1125(.a(s_83), .O(gate22inter4));
  nand2 gate1126(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate1127(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate1128(.a(G27), .O(gate22inter7));
  inv1  gate1129(.a(G28), .O(gate22inter8));
  nand2 gate1130(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate1131(.a(s_83), .b(gate22inter3), .O(gate22inter10));
  nor2  gate1132(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate1133(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate1134(.a(gate22inter12), .b(gate22inter1), .O(G305));
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate589(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate590(.a(gate24inter0), .b(s_6), .O(gate24inter1));
  and2  gate591(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate592(.a(s_6), .O(gate24inter3));
  inv1  gate593(.a(s_7), .O(gate24inter4));
  nand2 gate594(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate595(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate596(.a(G31), .O(gate24inter7));
  inv1  gate597(.a(G32), .O(gate24inter8));
  nand2 gate598(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate599(.a(s_7), .b(gate24inter3), .O(gate24inter10));
  nor2  gate600(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate601(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate602(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate687(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate688(.a(gate29inter0), .b(s_20), .O(gate29inter1));
  and2  gate689(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate690(.a(s_20), .O(gate29inter3));
  inv1  gate691(.a(s_21), .O(gate29inter4));
  nand2 gate692(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate693(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate694(.a(G3), .O(gate29inter7));
  inv1  gate695(.a(G7), .O(gate29inter8));
  nand2 gate696(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate697(.a(s_21), .b(gate29inter3), .O(gate29inter10));
  nor2  gate698(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate699(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate700(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate575(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate576(.a(gate34inter0), .b(s_4), .O(gate34inter1));
  and2  gate577(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate578(.a(s_4), .O(gate34inter3));
  inv1  gate579(.a(s_5), .O(gate34inter4));
  nand2 gate580(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate581(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate582(.a(G25), .O(gate34inter7));
  inv1  gate583(.a(G29), .O(gate34inter8));
  nand2 gate584(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate585(.a(s_5), .b(gate34inter3), .O(gate34inter10));
  nor2  gate586(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate587(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate588(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate981(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate982(.a(gate46inter0), .b(s_62), .O(gate46inter1));
  and2  gate983(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate984(.a(s_62), .O(gate46inter3));
  inv1  gate985(.a(s_63), .O(gate46inter4));
  nand2 gate986(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate987(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate988(.a(G6), .O(gate46inter7));
  inv1  gate989(.a(G272), .O(gate46inter8));
  nand2 gate990(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate991(.a(s_63), .b(gate46inter3), .O(gate46inter10));
  nor2  gate992(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate993(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate994(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate939(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate940(.a(gate65inter0), .b(s_56), .O(gate65inter1));
  and2  gate941(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate942(.a(s_56), .O(gate65inter3));
  inv1  gate943(.a(s_57), .O(gate65inter4));
  nand2 gate944(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate945(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate946(.a(G25), .O(gate65inter7));
  inv1  gate947(.a(G302), .O(gate65inter8));
  nand2 gate948(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate949(.a(s_57), .b(gate65inter3), .O(gate65inter10));
  nor2  gate950(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate951(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate952(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );

  xor2  gate547(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate548(.a(gate83inter0), .b(s_0), .O(gate83inter1));
  and2  gate549(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate550(.a(s_0), .O(gate83inter3));
  inv1  gate551(.a(s_1), .O(gate83inter4));
  nand2 gate552(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate553(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate554(.a(G11), .O(gate83inter7));
  inv1  gate555(.a(G329), .O(gate83inter8));
  nand2 gate556(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate557(.a(s_1), .b(gate83inter3), .O(gate83inter10));
  nor2  gate558(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate559(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate560(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate925(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate926(.a(gate86inter0), .b(s_54), .O(gate86inter1));
  and2  gate927(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate928(.a(s_54), .O(gate86inter3));
  inv1  gate929(.a(s_55), .O(gate86inter4));
  nand2 gate930(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate931(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate932(.a(G8), .O(gate86inter7));
  inv1  gate933(.a(G332), .O(gate86inter8));
  nand2 gate934(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate935(.a(s_55), .b(gate86inter3), .O(gate86inter10));
  nor2  gate936(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate937(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate938(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate1275(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate1276(.a(gate100inter0), .b(s_104), .O(gate100inter1));
  and2  gate1277(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate1278(.a(s_104), .O(gate100inter3));
  inv1  gate1279(.a(s_105), .O(gate100inter4));
  nand2 gate1280(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate1281(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate1282(.a(G31), .O(gate100inter7));
  inv1  gate1283(.a(G353), .O(gate100inter8));
  nand2 gate1284(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate1285(.a(s_105), .b(gate100inter3), .O(gate100inter10));
  nor2  gate1286(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate1287(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate1288(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );

  xor2  gate1233(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate1234(.a(gate103inter0), .b(s_98), .O(gate103inter1));
  and2  gate1235(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate1236(.a(s_98), .O(gate103inter3));
  inv1  gate1237(.a(s_99), .O(gate103inter4));
  nand2 gate1238(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate1239(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate1240(.a(G28), .O(gate103inter7));
  inv1  gate1241(.a(G359), .O(gate103inter8));
  nand2 gate1242(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate1243(.a(s_99), .b(gate103inter3), .O(gate103inter10));
  nor2  gate1244(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate1245(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate1246(.a(gate103inter12), .b(gate103inter1), .O(G424));
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate1219(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate1220(.a(gate119inter0), .b(s_96), .O(gate119inter1));
  and2  gate1221(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate1222(.a(s_96), .O(gate119inter3));
  inv1  gate1223(.a(s_97), .O(gate119inter4));
  nand2 gate1224(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate1225(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate1226(.a(G390), .O(gate119inter7));
  inv1  gate1227(.a(G391), .O(gate119inter8));
  nand2 gate1228(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate1229(.a(s_97), .b(gate119inter3), .O(gate119inter10));
  nor2  gate1230(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate1231(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate1232(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );

  xor2  gate743(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate744(.a(gate133inter0), .b(s_28), .O(gate133inter1));
  and2  gate745(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate746(.a(s_28), .O(gate133inter3));
  inv1  gate747(.a(s_29), .O(gate133inter4));
  nand2 gate748(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate749(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate750(.a(G418), .O(gate133inter7));
  inv1  gate751(.a(G419), .O(gate133inter8));
  nand2 gate752(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate753(.a(s_29), .b(gate133inter3), .O(gate133inter10));
  nor2  gate754(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate755(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate756(.a(gate133inter12), .b(gate133inter1), .O(G510));
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate1107(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate1108(.a(gate144inter0), .b(s_80), .O(gate144inter1));
  and2  gate1109(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate1110(.a(s_80), .O(gate144inter3));
  inv1  gate1111(.a(s_81), .O(gate144inter4));
  nand2 gate1112(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate1113(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate1114(.a(G468), .O(gate144inter7));
  inv1  gate1115(.a(G471), .O(gate144inter8));
  nand2 gate1116(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate1117(.a(s_81), .b(gate144inter3), .O(gate144inter10));
  nor2  gate1118(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate1119(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate1120(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate1303(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate1304(.a(gate155inter0), .b(s_108), .O(gate155inter1));
  and2  gate1305(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate1306(.a(s_108), .O(gate155inter3));
  inv1  gate1307(.a(s_109), .O(gate155inter4));
  nand2 gate1308(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1309(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1310(.a(G432), .O(gate155inter7));
  inv1  gate1311(.a(G525), .O(gate155inter8));
  nand2 gate1312(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1313(.a(s_109), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1314(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1315(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1316(.a(gate155inter12), .b(gate155inter1), .O(G572));

  xor2  gate897(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate898(.a(gate156inter0), .b(s_50), .O(gate156inter1));
  and2  gate899(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate900(.a(s_50), .O(gate156inter3));
  inv1  gate901(.a(s_51), .O(gate156inter4));
  nand2 gate902(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate903(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate904(.a(G435), .O(gate156inter7));
  inv1  gate905(.a(G525), .O(gate156inter8));
  nand2 gate906(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate907(.a(s_51), .b(gate156inter3), .O(gate156inter10));
  nor2  gate908(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate909(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate910(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate701(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate702(.a(gate160inter0), .b(s_22), .O(gate160inter1));
  and2  gate703(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate704(.a(s_22), .O(gate160inter3));
  inv1  gate705(.a(s_23), .O(gate160inter4));
  nand2 gate706(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate707(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate708(.a(G447), .O(gate160inter7));
  inv1  gate709(.a(G531), .O(gate160inter8));
  nand2 gate710(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate711(.a(s_23), .b(gate160inter3), .O(gate160inter10));
  nor2  gate712(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate713(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate714(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate1079(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate1080(.a(gate174inter0), .b(s_76), .O(gate174inter1));
  and2  gate1081(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate1082(.a(s_76), .O(gate174inter3));
  inv1  gate1083(.a(s_77), .O(gate174inter4));
  nand2 gate1084(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate1085(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate1086(.a(G489), .O(gate174inter7));
  inv1  gate1087(.a(G552), .O(gate174inter8));
  nand2 gate1088(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate1089(.a(s_77), .b(gate174inter3), .O(gate174inter10));
  nor2  gate1090(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate1091(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate1092(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate673(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate674(.a(gate185inter0), .b(s_18), .O(gate185inter1));
  and2  gate675(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate676(.a(s_18), .O(gate185inter3));
  inv1  gate677(.a(s_19), .O(gate185inter4));
  nand2 gate678(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate679(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate680(.a(G570), .O(gate185inter7));
  inv1  gate681(.a(G571), .O(gate185inter8));
  nand2 gate682(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate683(.a(s_19), .b(gate185inter3), .O(gate185inter10));
  nor2  gate684(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate685(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate686(.a(gate185inter12), .b(gate185inter1), .O(G602));
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate1037(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate1038(.a(gate191inter0), .b(s_70), .O(gate191inter1));
  and2  gate1039(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate1040(.a(s_70), .O(gate191inter3));
  inv1  gate1041(.a(s_71), .O(gate191inter4));
  nand2 gate1042(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate1043(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate1044(.a(G582), .O(gate191inter7));
  inv1  gate1045(.a(G583), .O(gate191inter8));
  nand2 gate1046(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate1047(.a(s_71), .b(gate191inter3), .O(gate191inter10));
  nor2  gate1048(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate1049(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate1050(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate841(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate842(.a(gate195inter0), .b(s_42), .O(gate195inter1));
  and2  gate843(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate844(.a(s_42), .O(gate195inter3));
  inv1  gate845(.a(s_43), .O(gate195inter4));
  nand2 gate846(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate847(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate848(.a(G590), .O(gate195inter7));
  inv1  gate849(.a(G591), .O(gate195inter8));
  nand2 gate850(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate851(.a(s_43), .b(gate195inter3), .O(gate195inter10));
  nor2  gate852(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate853(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate854(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate799(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate800(.a(gate201inter0), .b(s_36), .O(gate201inter1));
  and2  gate801(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate802(.a(s_36), .O(gate201inter3));
  inv1  gate803(.a(s_37), .O(gate201inter4));
  nand2 gate804(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate805(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate806(.a(G602), .O(gate201inter7));
  inv1  gate807(.a(G607), .O(gate201inter8));
  nand2 gate808(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate809(.a(s_37), .b(gate201inter3), .O(gate201inter10));
  nor2  gate810(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate811(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate812(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate1051(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate1052(.a(gate203inter0), .b(s_72), .O(gate203inter1));
  and2  gate1053(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate1054(.a(s_72), .O(gate203inter3));
  inv1  gate1055(.a(s_73), .O(gate203inter4));
  nand2 gate1056(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate1057(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate1058(.a(G602), .O(gate203inter7));
  inv1  gate1059(.a(G612), .O(gate203inter8));
  nand2 gate1060(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate1061(.a(s_73), .b(gate203inter3), .O(gate203inter10));
  nor2  gate1062(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate1063(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate1064(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );

  xor2  gate561(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate562(.a(gate208inter0), .b(s_2), .O(gate208inter1));
  and2  gate563(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate564(.a(s_2), .O(gate208inter3));
  inv1  gate565(.a(s_3), .O(gate208inter4));
  nand2 gate566(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate567(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate568(.a(G627), .O(gate208inter7));
  inv1  gate569(.a(G637), .O(gate208inter8));
  nand2 gate570(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate571(.a(s_3), .b(gate208inter3), .O(gate208inter10));
  nor2  gate572(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate573(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate574(.a(gate208inter12), .b(gate208inter1), .O(G687));
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate1317(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate1318(.a(gate211inter0), .b(s_110), .O(gate211inter1));
  and2  gate1319(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate1320(.a(s_110), .O(gate211inter3));
  inv1  gate1321(.a(s_111), .O(gate211inter4));
  nand2 gate1322(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate1323(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate1324(.a(G612), .O(gate211inter7));
  inv1  gate1325(.a(G669), .O(gate211inter8));
  nand2 gate1326(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate1327(.a(s_111), .b(gate211inter3), .O(gate211inter10));
  nor2  gate1328(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate1329(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate1330(.a(gate211inter12), .b(gate211inter1), .O(G692));
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );

  xor2  gate827(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate828(.a(gate221inter0), .b(s_40), .O(gate221inter1));
  and2  gate829(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate830(.a(s_40), .O(gate221inter3));
  inv1  gate831(.a(s_41), .O(gate221inter4));
  nand2 gate832(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate833(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate834(.a(G622), .O(gate221inter7));
  inv1  gate835(.a(G684), .O(gate221inter8));
  nand2 gate836(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate837(.a(s_41), .b(gate221inter3), .O(gate221inter10));
  nor2  gate838(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate839(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate840(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate855(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate856(.a(gate226inter0), .b(s_44), .O(gate226inter1));
  and2  gate857(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate858(.a(s_44), .O(gate226inter3));
  inv1  gate859(.a(s_45), .O(gate226inter4));
  nand2 gate860(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate861(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate862(.a(G692), .O(gate226inter7));
  inv1  gate863(.a(G693), .O(gate226inter8));
  nand2 gate864(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate865(.a(s_45), .b(gate226inter3), .O(gate226inter10));
  nor2  gate866(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate867(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate868(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate995(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate996(.a(gate236inter0), .b(s_64), .O(gate236inter1));
  and2  gate997(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate998(.a(s_64), .O(gate236inter3));
  inv1  gate999(.a(s_65), .O(gate236inter4));
  nand2 gate1000(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate1001(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate1002(.a(G251), .O(gate236inter7));
  inv1  gate1003(.a(G727), .O(gate236inter8));
  nand2 gate1004(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate1005(.a(s_65), .b(gate236inter3), .O(gate236inter10));
  nor2  gate1006(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate1007(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate1008(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate1023(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate1024(.a(gate250inter0), .b(s_68), .O(gate250inter1));
  and2  gate1025(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate1026(.a(s_68), .O(gate250inter3));
  inv1  gate1027(.a(s_69), .O(gate250inter4));
  nand2 gate1028(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate1029(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate1030(.a(G706), .O(gate250inter7));
  inv1  gate1031(.a(G742), .O(gate250inter8));
  nand2 gate1032(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate1033(.a(s_69), .b(gate250inter3), .O(gate250inter10));
  nor2  gate1034(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate1035(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate1036(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );

  xor2  gate1247(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate1248(.a(gate264inter0), .b(s_100), .O(gate264inter1));
  and2  gate1249(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate1250(.a(s_100), .O(gate264inter3));
  inv1  gate1251(.a(s_101), .O(gate264inter4));
  nand2 gate1252(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate1253(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate1254(.a(G768), .O(gate264inter7));
  inv1  gate1255(.a(G769), .O(gate264inter8));
  nand2 gate1256(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate1257(.a(s_101), .b(gate264inter3), .O(gate264inter10));
  nor2  gate1258(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate1259(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate1260(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );

  xor2  gate785(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate786(.a(gate273inter0), .b(s_34), .O(gate273inter1));
  and2  gate787(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate788(.a(s_34), .O(gate273inter3));
  inv1  gate789(.a(s_35), .O(gate273inter4));
  nand2 gate790(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate791(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate792(.a(G642), .O(gate273inter7));
  inv1  gate793(.a(G794), .O(gate273inter8));
  nand2 gate794(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate795(.a(s_35), .b(gate273inter3), .O(gate273inter10));
  nor2  gate796(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate797(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate798(.a(gate273inter12), .b(gate273inter1), .O(G818));
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate771(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate772(.a(gate286inter0), .b(s_32), .O(gate286inter1));
  and2  gate773(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate774(.a(s_32), .O(gate286inter3));
  inv1  gate775(.a(s_33), .O(gate286inter4));
  nand2 gate776(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate777(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate778(.a(G788), .O(gate286inter7));
  inv1  gate779(.a(G812), .O(gate286inter8));
  nand2 gate780(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate781(.a(s_33), .b(gate286inter3), .O(gate286inter10));
  nor2  gate782(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate783(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate784(.a(gate286inter12), .b(gate286inter1), .O(G831));
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate603(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate604(.a(gate290inter0), .b(s_8), .O(gate290inter1));
  and2  gate605(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate606(.a(s_8), .O(gate290inter3));
  inv1  gate607(.a(s_9), .O(gate290inter4));
  nand2 gate608(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate609(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate610(.a(G820), .O(gate290inter7));
  inv1  gate611(.a(G821), .O(gate290inter8));
  nand2 gate612(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate613(.a(s_9), .b(gate290inter3), .O(gate290inter10));
  nor2  gate614(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate615(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate616(.a(gate290inter12), .b(gate290inter1), .O(G847));

  xor2  gate869(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate870(.a(gate291inter0), .b(s_46), .O(gate291inter1));
  and2  gate871(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate872(.a(s_46), .O(gate291inter3));
  inv1  gate873(.a(s_47), .O(gate291inter4));
  nand2 gate874(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate875(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate876(.a(G822), .O(gate291inter7));
  inv1  gate877(.a(G823), .O(gate291inter8));
  nand2 gate878(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate879(.a(s_47), .b(gate291inter3), .O(gate291inter10));
  nor2  gate880(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate881(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate882(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate1093(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate1094(.a(gate387inter0), .b(s_78), .O(gate387inter1));
  and2  gate1095(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate1096(.a(s_78), .O(gate387inter3));
  inv1  gate1097(.a(s_79), .O(gate387inter4));
  nand2 gate1098(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1099(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1100(.a(G1), .O(gate387inter7));
  inv1  gate1101(.a(G1036), .O(gate387inter8));
  nand2 gate1102(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1103(.a(s_79), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1104(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1105(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate1106(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );

  xor2  gate967(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate968(.a(gate392inter0), .b(s_60), .O(gate392inter1));
  and2  gate969(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate970(.a(s_60), .O(gate392inter3));
  inv1  gate971(.a(s_61), .O(gate392inter4));
  nand2 gate972(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate973(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate974(.a(G6), .O(gate392inter7));
  inv1  gate975(.a(G1051), .O(gate392inter8));
  nand2 gate976(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate977(.a(s_61), .b(gate392inter3), .O(gate392inter10));
  nor2  gate978(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate979(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate980(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate883(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate884(.a(gate397inter0), .b(s_48), .O(gate397inter1));
  and2  gate885(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate886(.a(s_48), .O(gate397inter3));
  inv1  gate887(.a(s_49), .O(gate397inter4));
  nand2 gate888(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate889(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate890(.a(G11), .O(gate397inter7));
  inv1  gate891(.a(G1066), .O(gate397inter8));
  nand2 gate892(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate893(.a(s_49), .b(gate397inter3), .O(gate397inter10));
  nor2  gate894(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate895(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate896(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate617(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate618(.a(gate402inter0), .b(s_10), .O(gate402inter1));
  and2  gate619(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate620(.a(s_10), .O(gate402inter3));
  inv1  gate621(.a(s_11), .O(gate402inter4));
  nand2 gate622(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate623(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate624(.a(G16), .O(gate402inter7));
  inv1  gate625(.a(G1081), .O(gate402inter8));
  nand2 gate626(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate627(.a(s_11), .b(gate402inter3), .O(gate402inter10));
  nor2  gate628(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate629(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate630(.a(gate402inter12), .b(gate402inter1), .O(G1177));
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate1177(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate1178(.a(gate417inter0), .b(s_90), .O(gate417inter1));
  and2  gate1179(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate1180(.a(s_90), .O(gate417inter3));
  inv1  gate1181(.a(s_91), .O(gate417inter4));
  nand2 gate1182(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate1183(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate1184(.a(G31), .O(gate417inter7));
  inv1  gate1185(.a(G1126), .O(gate417inter8));
  nand2 gate1186(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate1187(.a(s_91), .b(gate417inter3), .O(gate417inter10));
  nor2  gate1188(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate1189(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate1190(.a(gate417inter12), .b(gate417inter1), .O(G1222));

  xor2  gate1135(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate1136(.a(gate418inter0), .b(s_84), .O(gate418inter1));
  and2  gate1137(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate1138(.a(s_84), .O(gate418inter3));
  inv1  gate1139(.a(s_85), .O(gate418inter4));
  nand2 gate1140(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate1141(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate1142(.a(G32), .O(gate418inter7));
  inv1  gate1143(.a(G1129), .O(gate418inter8));
  nand2 gate1144(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate1145(.a(s_85), .b(gate418inter3), .O(gate418inter10));
  nor2  gate1146(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate1147(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate1148(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate1261(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate1262(.a(gate422inter0), .b(s_102), .O(gate422inter1));
  and2  gate1263(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate1264(.a(s_102), .O(gate422inter3));
  inv1  gate1265(.a(s_103), .O(gate422inter4));
  nand2 gate1266(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate1267(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate1268(.a(G1039), .O(gate422inter7));
  inv1  gate1269(.a(G1135), .O(gate422inter8));
  nand2 gate1270(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate1271(.a(s_103), .b(gate422inter3), .O(gate422inter10));
  nor2  gate1272(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate1273(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate1274(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate813(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate814(.a(gate437inter0), .b(s_38), .O(gate437inter1));
  and2  gate815(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate816(.a(s_38), .O(gate437inter3));
  inv1  gate817(.a(s_39), .O(gate437inter4));
  nand2 gate818(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate819(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate820(.a(G10), .O(gate437inter7));
  inv1  gate821(.a(G1159), .O(gate437inter8));
  nand2 gate822(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate823(.a(s_39), .b(gate437inter3), .O(gate437inter10));
  nor2  gate824(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate825(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate826(.a(gate437inter12), .b(gate437inter1), .O(G1246));
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate1149(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate1150(.a(gate439inter0), .b(s_86), .O(gate439inter1));
  and2  gate1151(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate1152(.a(s_86), .O(gate439inter3));
  inv1  gate1153(.a(s_87), .O(gate439inter4));
  nand2 gate1154(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate1155(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate1156(.a(G11), .O(gate439inter7));
  inv1  gate1157(.a(G1162), .O(gate439inter8));
  nand2 gate1158(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate1159(.a(s_87), .b(gate439inter3), .O(gate439inter10));
  nor2  gate1160(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate1161(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate1162(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate729(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate730(.a(gate443inter0), .b(s_26), .O(gate443inter1));
  and2  gate731(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate732(.a(s_26), .O(gate443inter3));
  inv1  gate733(.a(s_27), .O(gate443inter4));
  nand2 gate734(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate735(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate736(.a(G13), .O(gate443inter7));
  inv1  gate737(.a(G1168), .O(gate443inter8));
  nand2 gate738(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate739(.a(s_27), .b(gate443inter3), .O(gate443inter10));
  nor2  gate740(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate741(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate742(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );

  xor2  gate631(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate632(.a(gate447inter0), .b(s_12), .O(gate447inter1));
  and2  gate633(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate634(.a(s_12), .O(gate447inter3));
  inv1  gate635(.a(s_13), .O(gate447inter4));
  nand2 gate636(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate637(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate638(.a(G15), .O(gate447inter7));
  inv1  gate639(.a(G1174), .O(gate447inter8));
  nand2 gate640(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate641(.a(s_13), .b(gate447inter3), .O(gate447inter10));
  nor2  gate642(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate643(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate644(.a(gate447inter12), .b(gate447inter1), .O(G1256));
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate1191(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate1192(.a(gate456inter0), .b(s_92), .O(gate456inter1));
  and2  gate1193(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate1194(.a(s_92), .O(gate456inter3));
  inv1  gate1195(.a(s_93), .O(gate456inter4));
  nand2 gate1196(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate1197(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate1198(.a(G1090), .O(gate456inter7));
  inv1  gate1199(.a(G1186), .O(gate456inter8));
  nand2 gate1200(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate1201(.a(s_93), .b(gate456inter3), .O(gate456inter10));
  nor2  gate1202(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate1203(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate1204(.a(gate456inter12), .b(gate456inter1), .O(G1265));

  xor2  gate645(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate646(.a(gate457inter0), .b(s_14), .O(gate457inter1));
  and2  gate647(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate648(.a(s_14), .O(gate457inter3));
  inv1  gate649(.a(s_15), .O(gate457inter4));
  nand2 gate650(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate651(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate652(.a(G20), .O(gate457inter7));
  inv1  gate653(.a(G1189), .O(gate457inter8));
  nand2 gate654(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate655(.a(s_15), .b(gate457inter3), .O(gate457inter10));
  nor2  gate656(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate657(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate658(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate911(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate912(.a(gate461inter0), .b(s_52), .O(gate461inter1));
  and2  gate913(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate914(.a(s_52), .O(gate461inter3));
  inv1  gate915(.a(s_53), .O(gate461inter4));
  nand2 gate916(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate917(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate918(.a(G22), .O(gate461inter7));
  inv1  gate919(.a(G1195), .O(gate461inter8));
  nand2 gate920(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate921(.a(s_53), .b(gate461inter3), .O(gate461inter10));
  nor2  gate922(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate923(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate924(.a(gate461inter12), .b(gate461inter1), .O(G1270));
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );

  xor2  gate757(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate758(.a(gate484inter0), .b(s_30), .O(gate484inter1));
  and2  gate759(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate760(.a(s_30), .O(gate484inter3));
  inv1  gate761(.a(s_31), .O(gate484inter4));
  nand2 gate762(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate763(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate764(.a(G1230), .O(gate484inter7));
  inv1  gate765(.a(G1231), .O(gate484inter8));
  nand2 gate766(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate767(.a(s_31), .b(gate484inter3), .O(gate484inter10));
  nor2  gate768(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate769(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate770(.a(gate484inter12), .b(gate484inter1), .O(G1293));
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate1065(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate1066(.a(gate486inter0), .b(s_74), .O(gate486inter1));
  and2  gate1067(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate1068(.a(s_74), .O(gate486inter3));
  inv1  gate1069(.a(s_75), .O(gate486inter4));
  nand2 gate1070(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate1071(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate1072(.a(G1234), .O(gate486inter7));
  inv1  gate1073(.a(G1235), .O(gate486inter8));
  nand2 gate1074(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate1075(.a(s_75), .b(gate486inter3), .O(gate486inter10));
  nor2  gate1076(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate1077(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate1078(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate1163(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1164(.a(gate494inter0), .b(s_88), .O(gate494inter1));
  and2  gate1165(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1166(.a(s_88), .O(gate494inter3));
  inv1  gate1167(.a(s_89), .O(gate494inter4));
  nand2 gate1168(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1169(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1170(.a(G1250), .O(gate494inter7));
  inv1  gate1171(.a(G1251), .O(gate494inter8));
  nand2 gate1172(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1173(.a(s_89), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1174(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1175(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1176(.a(gate494inter12), .b(gate494inter1), .O(G1303));

  xor2  gate715(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate716(.a(gate495inter0), .b(s_24), .O(gate495inter1));
  and2  gate717(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate718(.a(s_24), .O(gate495inter3));
  inv1  gate719(.a(s_25), .O(gate495inter4));
  nand2 gate720(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate721(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate722(.a(G1252), .O(gate495inter7));
  inv1  gate723(.a(G1253), .O(gate495inter8));
  nand2 gate724(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate725(.a(s_25), .b(gate495inter3), .O(gate495inter10));
  nor2  gate726(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate727(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate728(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate953(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate954(.a(gate499inter0), .b(s_58), .O(gate499inter1));
  and2  gate955(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate956(.a(s_58), .O(gate499inter3));
  inv1  gate957(.a(s_59), .O(gate499inter4));
  nand2 gate958(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate959(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate960(.a(G1260), .O(gate499inter7));
  inv1  gate961(.a(G1261), .O(gate499inter8));
  nand2 gate962(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate963(.a(s_59), .b(gate499inter3), .O(gate499inter10));
  nor2  gate964(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate965(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate966(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );

  xor2  gate1289(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate1290(.a(gate505inter0), .b(s_106), .O(gate505inter1));
  and2  gate1291(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate1292(.a(s_106), .O(gate505inter3));
  inv1  gate1293(.a(s_107), .O(gate505inter4));
  nand2 gate1294(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate1295(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate1296(.a(G1272), .O(gate505inter7));
  inv1  gate1297(.a(G1273), .O(gate505inter8));
  nand2 gate1298(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate1299(.a(s_107), .b(gate505inter3), .O(gate505inter10));
  nor2  gate1300(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate1301(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate1302(.a(gate505inter12), .b(gate505inter1), .O(G1314));
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate1009(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate1010(.a(gate510inter0), .b(s_66), .O(gate510inter1));
  and2  gate1011(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate1012(.a(s_66), .O(gate510inter3));
  inv1  gate1013(.a(s_67), .O(gate510inter4));
  nand2 gate1014(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate1015(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate1016(.a(G1282), .O(gate510inter7));
  inv1  gate1017(.a(G1283), .O(gate510inter8));
  nand2 gate1018(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate1019(.a(s_67), .b(gate510inter3), .O(gate510inter10));
  nor2  gate1020(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate1021(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate1022(.a(gate510inter12), .b(gate510inter1), .O(G1319));

  xor2  gate659(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate660(.a(gate511inter0), .b(s_16), .O(gate511inter1));
  and2  gate661(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate662(.a(s_16), .O(gate511inter3));
  inv1  gate663(.a(s_17), .O(gate511inter4));
  nand2 gate664(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate665(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate666(.a(G1284), .O(gate511inter7));
  inv1  gate667(.a(G1285), .O(gate511inter8));
  nand2 gate668(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate669(.a(s_17), .b(gate511inter3), .O(gate511inter10));
  nor2  gate670(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate671(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate672(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule