module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281, s_282, s_283, s_284, s_285, s_286, s_287, s_288, s_289, s_290, s_291, s_292, s_293, s_294, s_295, s_296, s_297, s_298, s_299, s_300, s_301, s_302, s_303, s_304, s_305, s_306, s_307, s_308, s_309, s_310, s_311;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate813(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate814(.a(gate9inter0), .b(s_38), .O(gate9inter1));
  and2  gate815(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate816(.a(s_38), .O(gate9inter3));
  inv1  gate817(.a(s_39), .O(gate9inter4));
  nand2 gate818(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate819(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate820(.a(G1), .O(gate9inter7));
  inv1  gate821(.a(G2), .O(gate9inter8));
  nand2 gate822(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate823(.a(s_39), .b(gate9inter3), .O(gate9inter10));
  nor2  gate824(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate825(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate826(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate561(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate562(.a(gate11inter0), .b(s_2), .O(gate11inter1));
  and2  gate563(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate564(.a(s_2), .O(gate11inter3));
  inv1  gate565(.a(s_3), .O(gate11inter4));
  nand2 gate566(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate567(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate568(.a(G5), .O(gate11inter7));
  inv1  gate569(.a(G6), .O(gate11inter8));
  nand2 gate570(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate571(.a(s_3), .b(gate11inter3), .O(gate11inter10));
  nor2  gate572(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate573(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate574(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );

  xor2  gate1191(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate1192(.a(gate14inter0), .b(s_92), .O(gate14inter1));
  and2  gate1193(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate1194(.a(s_92), .O(gate14inter3));
  inv1  gate1195(.a(s_93), .O(gate14inter4));
  nand2 gate1196(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate1197(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate1198(.a(G11), .O(gate14inter7));
  inv1  gate1199(.a(G12), .O(gate14inter8));
  nand2 gate1200(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate1201(.a(s_93), .b(gate14inter3), .O(gate14inter10));
  nor2  gate1202(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate1203(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate1204(.a(gate14inter12), .b(gate14inter1), .O(G281));

  xor2  gate1709(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate1710(.a(gate15inter0), .b(s_166), .O(gate15inter1));
  and2  gate1711(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate1712(.a(s_166), .O(gate15inter3));
  inv1  gate1713(.a(s_167), .O(gate15inter4));
  nand2 gate1714(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate1715(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate1716(.a(G13), .O(gate15inter7));
  inv1  gate1717(.a(G14), .O(gate15inter8));
  nand2 gate1718(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate1719(.a(s_167), .b(gate15inter3), .O(gate15inter10));
  nor2  gate1720(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate1721(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate1722(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate1219(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate1220(.a(gate17inter0), .b(s_96), .O(gate17inter1));
  and2  gate1221(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate1222(.a(s_96), .O(gate17inter3));
  inv1  gate1223(.a(s_97), .O(gate17inter4));
  nand2 gate1224(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate1225(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate1226(.a(G17), .O(gate17inter7));
  inv1  gate1227(.a(G18), .O(gate17inter8));
  nand2 gate1228(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate1229(.a(s_97), .b(gate17inter3), .O(gate17inter10));
  nor2  gate1230(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate1231(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate1232(.a(gate17inter12), .b(gate17inter1), .O(G290));

  xor2  gate2269(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate2270(.a(gate18inter0), .b(s_246), .O(gate18inter1));
  and2  gate2271(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate2272(.a(s_246), .O(gate18inter3));
  inv1  gate2273(.a(s_247), .O(gate18inter4));
  nand2 gate2274(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate2275(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate2276(.a(G19), .O(gate18inter7));
  inv1  gate2277(.a(G20), .O(gate18inter8));
  nand2 gate2278(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate2279(.a(s_247), .b(gate18inter3), .O(gate18inter10));
  nor2  gate2280(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate2281(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate2282(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate1821(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate1822(.a(gate20inter0), .b(s_182), .O(gate20inter1));
  and2  gate1823(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate1824(.a(s_182), .O(gate20inter3));
  inv1  gate1825(.a(s_183), .O(gate20inter4));
  nand2 gate1826(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate1827(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate1828(.a(G23), .O(gate20inter7));
  inv1  gate1829(.a(G24), .O(gate20inter8));
  nand2 gate1830(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate1831(.a(s_183), .b(gate20inter3), .O(gate20inter10));
  nor2  gate1832(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate1833(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate1834(.a(gate20inter12), .b(gate20inter1), .O(G299));

  xor2  gate2157(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate2158(.a(gate21inter0), .b(s_230), .O(gate21inter1));
  and2  gate2159(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate2160(.a(s_230), .O(gate21inter3));
  inv1  gate2161(.a(s_231), .O(gate21inter4));
  nand2 gate2162(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate2163(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate2164(.a(G25), .O(gate21inter7));
  inv1  gate2165(.a(G26), .O(gate21inter8));
  nand2 gate2166(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate2167(.a(s_231), .b(gate21inter3), .O(gate21inter10));
  nor2  gate2168(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate2169(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate2170(.a(gate21inter12), .b(gate21inter1), .O(G302));

  xor2  gate1667(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate1668(.a(gate22inter0), .b(s_160), .O(gate22inter1));
  and2  gate1669(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate1670(.a(s_160), .O(gate22inter3));
  inv1  gate1671(.a(s_161), .O(gate22inter4));
  nand2 gate1672(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate1673(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate1674(.a(G27), .O(gate22inter7));
  inv1  gate1675(.a(G28), .O(gate22inter8));
  nand2 gate1676(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate1677(.a(s_161), .b(gate22inter3), .O(gate22inter10));
  nor2  gate1678(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate1679(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate1680(.a(gate22inter12), .b(gate22inter1), .O(G305));

  xor2  gate2395(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate2396(.a(gate23inter0), .b(s_264), .O(gate23inter1));
  and2  gate2397(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate2398(.a(s_264), .O(gate23inter3));
  inv1  gate2399(.a(s_265), .O(gate23inter4));
  nand2 gate2400(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate2401(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate2402(.a(G29), .O(gate23inter7));
  inv1  gate2403(.a(G30), .O(gate23inter8));
  nand2 gate2404(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate2405(.a(s_265), .b(gate23inter3), .O(gate23inter10));
  nor2  gate2406(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate2407(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate2408(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate2605(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate2606(.a(gate26inter0), .b(s_294), .O(gate26inter1));
  and2  gate2607(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate2608(.a(s_294), .O(gate26inter3));
  inv1  gate2609(.a(s_295), .O(gate26inter4));
  nand2 gate2610(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate2611(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate2612(.a(G9), .O(gate26inter7));
  inv1  gate2613(.a(G13), .O(gate26inter8));
  nand2 gate2614(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate2615(.a(s_295), .b(gate26inter3), .O(gate26inter10));
  nor2  gate2616(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate2617(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate2618(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate1429(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate1430(.a(gate28inter0), .b(s_126), .O(gate28inter1));
  and2  gate1431(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate1432(.a(s_126), .O(gate28inter3));
  inv1  gate1433(.a(s_127), .O(gate28inter4));
  nand2 gate1434(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate1435(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate1436(.a(G10), .O(gate28inter7));
  inv1  gate1437(.a(G14), .O(gate28inter8));
  nand2 gate1438(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate1439(.a(s_127), .b(gate28inter3), .O(gate28inter10));
  nor2  gate1440(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate1441(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate1442(.a(gate28inter12), .b(gate28inter1), .O(G323));

  xor2  gate2297(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate2298(.a(gate29inter0), .b(s_250), .O(gate29inter1));
  and2  gate2299(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate2300(.a(s_250), .O(gate29inter3));
  inv1  gate2301(.a(s_251), .O(gate29inter4));
  nand2 gate2302(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate2303(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate2304(.a(G3), .O(gate29inter7));
  inv1  gate2305(.a(G7), .O(gate29inter8));
  nand2 gate2306(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate2307(.a(s_251), .b(gate29inter3), .O(gate29inter10));
  nor2  gate2308(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate2309(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate2310(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate1793(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate1794(.a(gate31inter0), .b(s_178), .O(gate31inter1));
  and2  gate1795(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate1796(.a(s_178), .O(gate31inter3));
  inv1  gate1797(.a(s_179), .O(gate31inter4));
  nand2 gate1798(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate1799(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate1800(.a(G4), .O(gate31inter7));
  inv1  gate1801(.a(G8), .O(gate31inter8));
  nand2 gate1802(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate1803(.a(s_179), .b(gate31inter3), .O(gate31inter10));
  nor2  gate1804(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate1805(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate1806(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate2199(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate2200(.a(gate34inter0), .b(s_236), .O(gate34inter1));
  and2  gate2201(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate2202(.a(s_236), .O(gate34inter3));
  inv1  gate2203(.a(s_237), .O(gate34inter4));
  nand2 gate2204(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate2205(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate2206(.a(G25), .O(gate34inter7));
  inv1  gate2207(.a(G29), .O(gate34inter8));
  nand2 gate2208(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate2209(.a(s_237), .b(gate34inter3), .O(gate34inter10));
  nor2  gate2210(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate2211(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate2212(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate2521(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate2522(.a(gate37inter0), .b(s_282), .O(gate37inter1));
  and2  gate2523(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate2524(.a(s_282), .O(gate37inter3));
  inv1  gate2525(.a(s_283), .O(gate37inter4));
  nand2 gate2526(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate2527(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate2528(.a(G19), .O(gate37inter7));
  inv1  gate2529(.a(G23), .O(gate37inter8));
  nand2 gate2530(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate2531(.a(s_283), .b(gate37inter3), .O(gate37inter10));
  nor2  gate2532(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate2533(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate2534(.a(gate37inter12), .b(gate37inter1), .O(G350));

  xor2  gate1387(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate1388(.a(gate38inter0), .b(s_120), .O(gate38inter1));
  and2  gate1389(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate1390(.a(s_120), .O(gate38inter3));
  inv1  gate1391(.a(s_121), .O(gate38inter4));
  nand2 gate1392(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate1393(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate1394(.a(G27), .O(gate38inter7));
  inv1  gate1395(.a(G31), .O(gate38inter8));
  nand2 gate1396(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate1397(.a(s_121), .b(gate38inter3), .O(gate38inter10));
  nor2  gate1398(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate1399(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate1400(.a(gate38inter12), .b(gate38inter1), .O(G353));

  xor2  gate1359(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate1360(.a(gate39inter0), .b(s_116), .O(gate39inter1));
  and2  gate1361(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate1362(.a(s_116), .O(gate39inter3));
  inv1  gate1363(.a(s_117), .O(gate39inter4));
  nand2 gate1364(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate1365(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate1366(.a(G20), .O(gate39inter7));
  inv1  gate1367(.a(G24), .O(gate39inter8));
  nand2 gate1368(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate1369(.a(s_117), .b(gate39inter3), .O(gate39inter10));
  nor2  gate1370(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate1371(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate1372(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate2143(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate2144(.a(gate41inter0), .b(s_228), .O(gate41inter1));
  and2  gate2145(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate2146(.a(s_228), .O(gate41inter3));
  inv1  gate2147(.a(s_229), .O(gate41inter4));
  nand2 gate2148(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate2149(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate2150(.a(G1), .O(gate41inter7));
  inv1  gate2151(.a(G266), .O(gate41inter8));
  nand2 gate2152(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate2153(.a(s_229), .b(gate41inter3), .O(gate41inter10));
  nor2  gate2154(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate2155(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate2156(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );

  xor2  gate1317(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate1318(.a(gate45inter0), .b(s_110), .O(gate45inter1));
  and2  gate1319(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate1320(.a(s_110), .O(gate45inter3));
  inv1  gate1321(.a(s_111), .O(gate45inter4));
  nand2 gate1322(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate1323(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate1324(.a(G5), .O(gate45inter7));
  inv1  gate1325(.a(G272), .O(gate45inter8));
  nand2 gate1326(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate1327(.a(s_111), .b(gate45inter3), .O(gate45inter10));
  nor2  gate1328(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate1329(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate1330(.a(gate45inter12), .b(gate45inter1), .O(G366));

  xor2  gate1891(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate1892(.a(gate46inter0), .b(s_192), .O(gate46inter1));
  and2  gate1893(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate1894(.a(s_192), .O(gate46inter3));
  inv1  gate1895(.a(s_193), .O(gate46inter4));
  nand2 gate1896(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate1897(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate1898(.a(G6), .O(gate46inter7));
  inv1  gate1899(.a(G272), .O(gate46inter8));
  nand2 gate1900(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate1901(.a(s_193), .b(gate46inter3), .O(gate46inter10));
  nor2  gate1902(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate1903(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate1904(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate799(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate800(.a(gate55inter0), .b(s_36), .O(gate55inter1));
  and2  gate801(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate802(.a(s_36), .O(gate55inter3));
  inv1  gate803(.a(s_37), .O(gate55inter4));
  nand2 gate804(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate805(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate806(.a(G15), .O(gate55inter7));
  inv1  gate807(.a(G287), .O(gate55inter8));
  nand2 gate808(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate809(.a(s_37), .b(gate55inter3), .O(gate55inter10));
  nor2  gate810(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate811(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate812(.a(gate55inter12), .b(gate55inter1), .O(G376));

  xor2  gate2255(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate2256(.a(gate56inter0), .b(s_244), .O(gate56inter1));
  and2  gate2257(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate2258(.a(s_244), .O(gate56inter3));
  inv1  gate2259(.a(s_245), .O(gate56inter4));
  nand2 gate2260(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate2261(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate2262(.a(G16), .O(gate56inter7));
  inv1  gate2263(.a(G287), .O(gate56inter8));
  nand2 gate2264(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate2265(.a(s_245), .b(gate56inter3), .O(gate56inter10));
  nor2  gate2266(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate2267(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate2268(.a(gate56inter12), .b(gate56inter1), .O(G377));

  xor2  gate2227(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate2228(.a(gate57inter0), .b(s_240), .O(gate57inter1));
  and2  gate2229(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate2230(.a(s_240), .O(gate57inter3));
  inv1  gate2231(.a(s_241), .O(gate57inter4));
  nand2 gate2232(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate2233(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate2234(.a(G17), .O(gate57inter7));
  inv1  gate2235(.a(G290), .O(gate57inter8));
  nand2 gate2236(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate2237(.a(s_241), .b(gate57inter3), .O(gate57inter10));
  nor2  gate2238(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate2239(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate2240(.a(gate57inter12), .b(gate57inter1), .O(G378));
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );

  xor2  gate2171(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate2172(.a(gate61inter0), .b(s_232), .O(gate61inter1));
  and2  gate2173(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate2174(.a(s_232), .O(gate61inter3));
  inv1  gate2175(.a(s_233), .O(gate61inter4));
  nand2 gate2176(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate2177(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate2178(.a(G21), .O(gate61inter7));
  inv1  gate2179(.a(G296), .O(gate61inter8));
  nand2 gate2180(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate2181(.a(s_233), .b(gate61inter3), .O(gate61inter10));
  nor2  gate2182(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate2183(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate2184(.a(gate61inter12), .b(gate61inter1), .O(G382));
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate1415(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate1416(.a(gate63inter0), .b(s_124), .O(gate63inter1));
  and2  gate1417(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate1418(.a(s_124), .O(gate63inter3));
  inv1  gate1419(.a(s_125), .O(gate63inter4));
  nand2 gate1420(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate1421(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate1422(.a(G23), .O(gate63inter7));
  inv1  gate1423(.a(G299), .O(gate63inter8));
  nand2 gate1424(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate1425(.a(s_125), .b(gate63inter3), .O(gate63inter10));
  nor2  gate1426(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate1427(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate1428(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate1625(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate1626(.a(gate65inter0), .b(s_154), .O(gate65inter1));
  and2  gate1627(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate1628(.a(s_154), .O(gate65inter3));
  inv1  gate1629(.a(s_155), .O(gate65inter4));
  nand2 gate1630(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate1631(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate1632(.a(G25), .O(gate65inter7));
  inv1  gate1633(.a(G302), .O(gate65inter8));
  nand2 gate1634(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate1635(.a(s_155), .b(gate65inter3), .O(gate65inter10));
  nor2  gate1636(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate1637(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate1638(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate2535(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate2536(.a(gate67inter0), .b(s_284), .O(gate67inter1));
  and2  gate2537(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate2538(.a(s_284), .O(gate67inter3));
  inv1  gate2539(.a(s_285), .O(gate67inter4));
  nand2 gate2540(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate2541(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate2542(.a(G27), .O(gate67inter7));
  inv1  gate2543(.a(G305), .O(gate67inter8));
  nand2 gate2544(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate2545(.a(s_285), .b(gate67inter3), .O(gate67inter10));
  nor2  gate2546(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate2547(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate2548(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate2339(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate2340(.a(gate70inter0), .b(s_256), .O(gate70inter1));
  and2  gate2341(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate2342(.a(s_256), .O(gate70inter3));
  inv1  gate2343(.a(s_257), .O(gate70inter4));
  nand2 gate2344(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate2345(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate2346(.a(G30), .O(gate70inter7));
  inv1  gate2347(.a(G308), .O(gate70inter8));
  nand2 gate2348(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate2349(.a(s_257), .b(gate70inter3), .O(gate70inter10));
  nor2  gate2350(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate2351(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate2352(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate1135(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate1136(.a(gate80inter0), .b(s_84), .O(gate80inter1));
  and2  gate1137(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate1138(.a(s_84), .O(gate80inter3));
  inv1  gate1139(.a(s_85), .O(gate80inter4));
  nand2 gate1140(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate1141(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate1142(.a(G14), .O(gate80inter7));
  inv1  gate1143(.a(G323), .O(gate80inter8));
  nand2 gate1144(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate1145(.a(s_85), .b(gate80inter3), .O(gate80inter10));
  nor2  gate1146(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate1147(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate1148(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );

  xor2  gate883(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate884(.a(gate83inter0), .b(s_48), .O(gate83inter1));
  and2  gate885(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate886(.a(s_48), .O(gate83inter3));
  inv1  gate887(.a(s_49), .O(gate83inter4));
  nand2 gate888(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate889(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate890(.a(G11), .O(gate83inter7));
  inv1  gate891(.a(G329), .O(gate83inter8));
  nand2 gate892(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate893(.a(s_49), .b(gate83inter3), .O(gate83inter10));
  nor2  gate894(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate895(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate896(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate1163(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate1164(.a(gate85inter0), .b(s_88), .O(gate85inter1));
  and2  gate1165(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate1166(.a(s_88), .O(gate85inter3));
  inv1  gate1167(.a(s_89), .O(gate85inter4));
  nand2 gate1168(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate1169(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate1170(.a(G4), .O(gate85inter7));
  inv1  gate1171(.a(G332), .O(gate85inter8));
  nand2 gate1172(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate1173(.a(s_89), .b(gate85inter3), .O(gate85inter10));
  nor2  gate1174(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate1175(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate1176(.a(gate85inter12), .b(gate85inter1), .O(G406));

  xor2  gate2003(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate2004(.a(gate86inter0), .b(s_208), .O(gate86inter1));
  and2  gate2005(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate2006(.a(s_208), .O(gate86inter3));
  inv1  gate2007(.a(s_209), .O(gate86inter4));
  nand2 gate2008(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate2009(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate2010(.a(G8), .O(gate86inter7));
  inv1  gate2011(.a(G332), .O(gate86inter8));
  nand2 gate2012(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate2013(.a(s_209), .b(gate86inter3), .O(gate86inter10));
  nor2  gate2014(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate2015(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate2016(.a(gate86inter12), .b(gate86inter1), .O(G407));

  xor2  gate1009(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate1010(.a(gate87inter0), .b(s_66), .O(gate87inter1));
  and2  gate1011(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate1012(.a(s_66), .O(gate87inter3));
  inv1  gate1013(.a(s_67), .O(gate87inter4));
  nand2 gate1014(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate1015(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate1016(.a(G12), .O(gate87inter7));
  inv1  gate1017(.a(G335), .O(gate87inter8));
  nand2 gate1018(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate1019(.a(s_67), .b(gate87inter3), .O(gate87inter10));
  nor2  gate1020(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate1021(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate1022(.a(gate87inter12), .b(gate87inter1), .O(G408));

  xor2  gate1331(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate1332(.a(gate88inter0), .b(s_112), .O(gate88inter1));
  and2  gate1333(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate1334(.a(s_112), .O(gate88inter3));
  inv1  gate1335(.a(s_113), .O(gate88inter4));
  nand2 gate1336(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate1337(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate1338(.a(G16), .O(gate88inter7));
  inv1  gate1339(.a(G335), .O(gate88inter8));
  nand2 gate1340(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate1341(.a(s_113), .b(gate88inter3), .O(gate88inter10));
  nor2  gate1342(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate1343(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate1344(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );

  xor2  gate2073(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate2074(.a(gate93inter0), .b(s_218), .O(gate93inter1));
  and2  gate2075(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate2076(.a(s_218), .O(gate93inter3));
  inv1  gate2077(.a(s_219), .O(gate93inter4));
  nand2 gate2078(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate2079(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate2080(.a(G18), .O(gate93inter7));
  inv1  gate2081(.a(G344), .O(gate93inter8));
  nand2 gate2082(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate2083(.a(s_219), .b(gate93inter3), .O(gate93inter10));
  nor2  gate2084(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate2085(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate2086(.a(gate93inter12), .b(gate93inter1), .O(G414));

  xor2  gate673(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate674(.a(gate94inter0), .b(s_18), .O(gate94inter1));
  and2  gate675(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate676(.a(s_18), .O(gate94inter3));
  inv1  gate677(.a(s_19), .O(gate94inter4));
  nand2 gate678(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate679(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate680(.a(G22), .O(gate94inter7));
  inv1  gate681(.a(G344), .O(gate94inter8));
  nand2 gate682(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate683(.a(s_19), .b(gate94inter3), .O(gate94inter10));
  nor2  gate684(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate685(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate686(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate995(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate996(.a(gate96inter0), .b(s_64), .O(gate96inter1));
  and2  gate997(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate998(.a(s_64), .O(gate96inter3));
  inv1  gate999(.a(s_65), .O(gate96inter4));
  nand2 gate1000(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate1001(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate1002(.a(G30), .O(gate96inter7));
  inv1  gate1003(.a(G347), .O(gate96inter8));
  nand2 gate1004(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate1005(.a(s_65), .b(gate96inter3), .O(gate96inter10));
  nor2  gate1006(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate1007(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate1008(.a(gate96inter12), .b(gate96inter1), .O(G417));
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate1527(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate1528(.a(gate99inter0), .b(s_140), .O(gate99inter1));
  and2  gate1529(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate1530(.a(s_140), .O(gate99inter3));
  inv1  gate1531(.a(s_141), .O(gate99inter4));
  nand2 gate1532(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate1533(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate1534(.a(G27), .O(gate99inter7));
  inv1  gate1535(.a(G353), .O(gate99inter8));
  nand2 gate1536(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate1537(.a(s_141), .b(gate99inter3), .O(gate99inter10));
  nor2  gate1538(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate1539(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate1540(.a(gate99inter12), .b(gate99inter1), .O(G420));

  xor2  gate2577(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate2578(.a(gate100inter0), .b(s_290), .O(gate100inter1));
  and2  gate2579(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate2580(.a(s_290), .O(gate100inter3));
  inv1  gate2581(.a(s_291), .O(gate100inter4));
  nand2 gate2582(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate2583(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate2584(.a(G31), .O(gate100inter7));
  inv1  gate2585(.a(G353), .O(gate100inter8));
  nand2 gate2586(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate2587(.a(s_291), .b(gate100inter3), .O(gate100inter10));
  nor2  gate2588(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate2589(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate2590(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate2619(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate2620(.a(gate102inter0), .b(s_296), .O(gate102inter1));
  and2  gate2621(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate2622(.a(s_296), .O(gate102inter3));
  inv1  gate2623(.a(s_297), .O(gate102inter4));
  nand2 gate2624(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate2625(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate2626(.a(G24), .O(gate102inter7));
  inv1  gate2627(.a(G356), .O(gate102inter8));
  nand2 gate2628(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate2629(.a(s_297), .b(gate102inter3), .O(gate102inter10));
  nor2  gate2630(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate2631(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate2632(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate1849(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate1850(.a(gate107inter0), .b(s_186), .O(gate107inter1));
  and2  gate1851(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate1852(.a(s_186), .O(gate107inter3));
  inv1  gate1853(.a(s_187), .O(gate107inter4));
  nand2 gate1854(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate1855(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate1856(.a(G366), .O(gate107inter7));
  inv1  gate1857(.a(G367), .O(gate107inter8));
  nand2 gate1858(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate1859(.a(s_187), .b(gate107inter3), .O(gate107inter10));
  nor2  gate1860(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate1861(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate1862(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );

  xor2  gate1261(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate1262(.a(gate113inter0), .b(s_102), .O(gate113inter1));
  and2  gate1263(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate1264(.a(s_102), .O(gate113inter3));
  inv1  gate1265(.a(s_103), .O(gate113inter4));
  nand2 gate1266(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate1267(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate1268(.a(G378), .O(gate113inter7));
  inv1  gate1269(.a(G379), .O(gate113inter8));
  nand2 gate1270(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate1271(.a(s_103), .b(gate113inter3), .O(gate113inter10));
  nor2  gate1272(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate1273(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate1274(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate2367(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate2368(.a(gate115inter0), .b(s_260), .O(gate115inter1));
  and2  gate2369(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate2370(.a(s_260), .O(gate115inter3));
  inv1  gate2371(.a(s_261), .O(gate115inter4));
  nand2 gate2372(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate2373(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate2374(.a(G382), .O(gate115inter7));
  inv1  gate2375(.a(G383), .O(gate115inter8));
  nand2 gate2376(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate2377(.a(s_261), .b(gate115inter3), .O(gate115inter10));
  nor2  gate2378(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate2379(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate2380(.a(gate115inter12), .b(gate115inter1), .O(G456));

  xor2  gate1919(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate1920(.a(gate116inter0), .b(s_196), .O(gate116inter1));
  and2  gate1921(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate1922(.a(s_196), .O(gate116inter3));
  inv1  gate1923(.a(s_197), .O(gate116inter4));
  nand2 gate1924(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate1925(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate1926(.a(G384), .O(gate116inter7));
  inv1  gate1927(.a(G385), .O(gate116inter8));
  nand2 gate1928(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate1929(.a(s_197), .b(gate116inter3), .O(gate116inter10));
  nor2  gate1930(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate1931(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate1932(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate2325(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate2326(.a(gate119inter0), .b(s_254), .O(gate119inter1));
  and2  gate2327(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate2328(.a(s_254), .O(gate119inter3));
  inv1  gate2329(.a(s_255), .O(gate119inter4));
  nand2 gate2330(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate2331(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate2332(.a(G390), .O(gate119inter7));
  inv1  gate2333(.a(G391), .O(gate119inter8));
  nand2 gate2334(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate2335(.a(s_255), .b(gate119inter3), .O(gate119inter10));
  nor2  gate2336(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate2337(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate2338(.a(gate119inter12), .b(gate119inter1), .O(G468));

  xor2  gate1093(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate1094(.a(gate120inter0), .b(s_78), .O(gate120inter1));
  and2  gate1095(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate1096(.a(s_78), .O(gate120inter3));
  inv1  gate1097(.a(s_79), .O(gate120inter4));
  nand2 gate1098(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate1099(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate1100(.a(G392), .O(gate120inter7));
  inv1  gate1101(.a(G393), .O(gate120inter8));
  nand2 gate1102(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate1103(.a(s_79), .b(gate120inter3), .O(gate120inter10));
  nor2  gate1104(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate1105(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate1106(.a(gate120inter12), .b(gate120inter1), .O(G471));
nand2 gate121( .a(G394), .b(G395), .O(G474) );

  xor2  gate925(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate926(.a(gate122inter0), .b(s_54), .O(gate122inter1));
  and2  gate927(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate928(.a(s_54), .O(gate122inter3));
  inv1  gate929(.a(s_55), .O(gate122inter4));
  nand2 gate930(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate931(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate932(.a(G396), .O(gate122inter7));
  inv1  gate933(.a(G397), .O(gate122inter8));
  nand2 gate934(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate935(.a(s_55), .b(gate122inter3), .O(gate122inter10));
  nor2  gate936(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate937(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate938(.a(gate122inter12), .b(gate122inter1), .O(G477));

  xor2  gate967(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate968(.a(gate123inter0), .b(s_60), .O(gate123inter1));
  and2  gate969(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate970(.a(s_60), .O(gate123inter3));
  inv1  gate971(.a(s_61), .O(gate123inter4));
  nand2 gate972(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate973(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate974(.a(G398), .O(gate123inter7));
  inv1  gate975(.a(G399), .O(gate123inter8));
  nand2 gate976(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate977(.a(s_61), .b(gate123inter3), .O(gate123inter10));
  nor2  gate978(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate979(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate980(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );

  xor2  gate981(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate982(.a(gate127inter0), .b(s_62), .O(gate127inter1));
  and2  gate983(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate984(.a(s_62), .O(gate127inter3));
  inv1  gate985(.a(s_63), .O(gate127inter4));
  nand2 gate986(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate987(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate988(.a(G406), .O(gate127inter7));
  inv1  gate989(.a(G407), .O(gate127inter8));
  nand2 gate990(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate991(.a(s_63), .b(gate127inter3), .O(gate127inter10));
  nor2  gate992(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate993(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate994(.a(gate127inter12), .b(gate127inter1), .O(G492));

  xor2  gate2087(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate2088(.a(gate128inter0), .b(s_220), .O(gate128inter1));
  and2  gate2089(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate2090(.a(s_220), .O(gate128inter3));
  inv1  gate2091(.a(s_221), .O(gate128inter4));
  nand2 gate2092(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate2093(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate2094(.a(G408), .O(gate128inter7));
  inv1  gate2095(.a(G409), .O(gate128inter8));
  nand2 gate2096(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate2097(.a(s_221), .b(gate128inter3), .O(gate128inter10));
  nor2  gate2098(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate2099(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate2100(.a(gate128inter12), .b(gate128inter1), .O(G495));
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate2129(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate2130(.a(gate132inter0), .b(s_226), .O(gate132inter1));
  and2  gate2131(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate2132(.a(s_226), .O(gate132inter3));
  inv1  gate2133(.a(s_227), .O(gate132inter4));
  nand2 gate2134(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate2135(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate2136(.a(G416), .O(gate132inter7));
  inv1  gate2137(.a(G417), .O(gate132inter8));
  nand2 gate2138(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate2139(.a(s_227), .b(gate132inter3), .O(gate132inter10));
  nor2  gate2140(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate2141(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate2142(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate939(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate940(.a(gate135inter0), .b(s_56), .O(gate135inter1));
  and2  gate941(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate942(.a(s_56), .O(gate135inter3));
  inv1  gate943(.a(s_57), .O(gate135inter4));
  nand2 gate944(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate945(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate946(.a(G422), .O(gate135inter7));
  inv1  gate947(.a(G423), .O(gate135inter8));
  nand2 gate948(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate949(.a(s_57), .b(gate135inter3), .O(gate135inter10));
  nor2  gate950(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate951(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate952(.a(gate135inter12), .b(gate135inter1), .O(G516));
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate2353(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate2354(.a(gate143inter0), .b(s_258), .O(gate143inter1));
  and2  gate2355(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate2356(.a(s_258), .O(gate143inter3));
  inv1  gate2357(.a(s_259), .O(gate143inter4));
  nand2 gate2358(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate2359(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate2360(.a(G462), .O(gate143inter7));
  inv1  gate2361(.a(G465), .O(gate143inter8));
  nand2 gate2362(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate2363(.a(s_259), .b(gate143inter3), .O(gate143inter10));
  nor2  gate2364(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate2365(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate2366(.a(gate143inter12), .b(gate143inter1), .O(G540));

  xor2  gate1513(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate1514(.a(gate144inter0), .b(s_138), .O(gate144inter1));
  and2  gate1515(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate1516(.a(s_138), .O(gate144inter3));
  inv1  gate1517(.a(s_139), .O(gate144inter4));
  nand2 gate1518(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate1519(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate1520(.a(G468), .O(gate144inter7));
  inv1  gate1521(.a(G471), .O(gate144inter8));
  nand2 gate1522(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate1523(.a(s_139), .b(gate144inter3), .O(gate144inter10));
  nor2  gate1524(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate1525(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate1526(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate1373(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1374(.a(gate148inter0), .b(s_118), .O(gate148inter1));
  and2  gate1375(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1376(.a(s_118), .O(gate148inter3));
  inv1  gate1377(.a(s_119), .O(gate148inter4));
  nand2 gate1378(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1379(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1380(.a(G492), .O(gate148inter7));
  inv1  gate1381(.a(G495), .O(gate148inter8));
  nand2 gate1382(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1383(.a(s_119), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1384(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1385(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1386(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate869(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate870(.a(gate150inter0), .b(s_46), .O(gate150inter1));
  and2  gate871(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate872(.a(s_46), .O(gate150inter3));
  inv1  gate873(.a(s_47), .O(gate150inter4));
  nand2 gate874(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate875(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate876(.a(G504), .O(gate150inter7));
  inv1  gate877(.a(G507), .O(gate150inter8));
  nand2 gate878(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate879(.a(s_47), .b(gate150inter3), .O(gate150inter10));
  nor2  gate880(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate881(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate882(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );

  xor2  gate1653(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate1654(.a(gate152inter0), .b(s_158), .O(gate152inter1));
  and2  gate1655(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate1656(.a(s_158), .O(gate152inter3));
  inv1  gate1657(.a(s_159), .O(gate152inter4));
  nand2 gate1658(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate1659(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate1660(.a(G516), .O(gate152inter7));
  inv1  gate1661(.a(G519), .O(gate152inter8));
  nand2 gate1662(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate1663(.a(s_159), .b(gate152inter3), .O(gate152inter10));
  nor2  gate1664(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate1665(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate1666(.a(gate152inter12), .b(gate152inter1), .O(G567));
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate645(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate646(.a(gate155inter0), .b(s_14), .O(gate155inter1));
  and2  gate647(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate648(.a(s_14), .O(gate155inter3));
  inv1  gate649(.a(s_15), .O(gate155inter4));
  nand2 gate650(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate651(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate652(.a(G432), .O(gate155inter7));
  inv1  gate653(.a(G525), .O(gate155inter8));
  nand2 gate654(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate655(.a(s_15), .b(gate155inter3), .O(gate155inter10));
  nor2  gate656(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate657(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate658(.a(gate155inter12), .b(gate155inter1), .O(G572));

  xor2  gate1807(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate1808(.a(gate156inter0), .b(s_180), .O(gate156inter1));
  and2  gate1809(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate1810(.a(s_180), .O(gate156inter3));
  inv1  gate1811(.a(s_181), .O(gate156inter4));
  nand2 gate1812(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate1813(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate1814(.a(G435), .O(gate156inter7));
  inv1  gate1815(.a(G525), .O(gate156inter8));
  nand2 gate1816(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate1817(.a(s_181), .b(gate156inter3), .O(gate156inter10));
  nor2  gate1818(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate1819(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate1820(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate1611(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate1612(.a(gate159inter0), .b(s_152), .O(gate159inter1));
  and2  gate1613(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate1614(.a(s_152), .O(gate159inter3));
  inv1  gate1615(.a(s_153), .O(gate159inter4));
  nand2 gate1616(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate1617(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate1618(.a(G444), .O(gate159inter7));
  inv1  gate1619(.a(G531), .O(gate159inter8));
  nand2 gate1620(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate1621(.a(s_153), .b(gate159inter3), .O(gate159inter10));
  nor2  gate1622(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate1623(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate1624(.a(gate159inter12), .b(gate159inter1), .O(G576));

  xor2  gate2101(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate2102(.a(gate160inter0), .b(s_222), .O(gate160inter1));
  and2  gate2103(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate2104(.a(s_222), .O(gate160inter3));
  inv1  gate2105(.a(s_223), .O(gate160inter4));
  nand2 gate2106(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate2107(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate2108(.a(G447), .O(gate160inter7));
  inv1  gate2109(.a(G531), .O(gate160inter8));
  nand2 gate2110(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate2111(.a(s_223), .b(gate160inter3), .O(gate160inter10));
  nor2  gate2112(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate2113(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate2114(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate2059(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate2060(.a(gate164inter0), .b(s_216), .O(gate164inter1));
  and2  gate2061(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate2062(.a(s_216), .O(gate164inter3));
  inv1  gate2063(.a(s_217), .O(gate164inter4));
  nand2 gate2064(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate2065(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate2066(.a(G459), .O(gate164inter7));
  inv1  gate2067(.a(G537), .O(gate164inter8));
  nand2 gate2068(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate2069(.a(s_217), .b(gate164inter3), .O(gate164inter10));
  nor2  gate2070(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate2071(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate2072(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );

  xor2  gate771(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate772(.a(gate166inter0), .b(s_32), .O(gate166inter1));
  and2  gate773(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate774(.a(s_32), .O(gate166inter3));
  inv1  gate775(.a(s_33), .O(gate166inter4));
  nand2 gate776(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate777(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate778(.a(G465), .O(gate166inter7));
  inv1  gate779(.a(G540), .O(gate166inter8));
  nand2 gate780(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate781(.a(s_33), .b(gate166inter3), .O(gate166inter10));
  nor2  gate782(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate783(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate784(.a(gate166inter12), .b(gate166inter1), .O(G583));

  xor2  gate1079(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate1080(.a(gate167inter0), .b(s_76), .O(gate167inter1));
  and2  gate1081(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate1082(.a(s_76), .O(gate167inter3));
  inv1  gate1083(.a(s_77), .O(gate167inter4));
  nand2 gate1084(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate1085(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate1086(.a(G468), .O(gate167inter7));
  inv1  gate1087(.a(G543), .O(gate167inter8));
  nand2 gate1088(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate1089(.a(s_77), .b(gate167inter3), .O(gate167inter10));
  nor2  gate1090(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate1091(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate1092(.a(gate167inter12), .b(gate167inter1), .O(G584));

  xor2  gate1905(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate1906(.a(gate168inter0), .b(s_194), .O(gate168inter1));
  and2  gate1907(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate1908(.a(s_194), .O(gate168inter3));
  inv1  gate1909(.a(s_195), .O(gate168inter4));
  nand2 gate1910(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate1911(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate1912(.a(G471), .O(gate168inter7));
  inv1  gate1913(.a(G543), .O(gate168inter8));
  nand2 gate1914(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate1915(.a(s_195), .b(gate168inter3), .O(gate168inter10));
  nor2  gate1916(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate1917(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate1918(.a(gate168inter12), .b(gate168inter1), .O(G585));

  xor2  gate2549(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate2550(.a(gate169inter0), .b(s_286), .O(gate169inter1));
  and2  gate2551(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate2552(.a(s_286), .O(gate169inter3));
  inv1  gate2553(.a(s_287), .O(gate169inter4));
  nand2 gate2554(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate2555(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate2556(.a(G474), .O(gate169inter7));
  inv1  gate2557(.a(G546), .O(gate169inter8));
  nand2 gate2558(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate2559(.a(s_287), .b(gate169inter3), .O(gate169inter10));
  nor2  gate2560(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate2561(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate2562(.a(gate169inter12), .b(gate169inter1), .O(G586));
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate1023(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate1024(.a(gate172inter0), .b(s_68), .O(gate172inter1));
  and2  gate1025(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate1026(.a(s_68), .O(gate172inter3));
  inv1  gate1027(.a(s_69), .O(gate172inter4));
  nand2 gate1028(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate1029(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate1030(.a(G483), .O(gate172inter7));
  inv1  gate1031(.a(G549), .O(gate172inter8));
  nand2 gate1032(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate1033(.a(s_69), .b(gate172inter3), .O(gate172inter10));
  nor2  gate1034(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate1035(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate1036(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate2661(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate2662(.a(gate174inter0), .b(s_302), .O(gate174inter1));
  and2  gate2663(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate2664(.a(s_302), .O(gate174inter3));
  inv1  gate2665(.a(s_303), .O(gate174inter4));
  nand2 gate2666(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate2667(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate2668(.a(G489), .O(gate174inter7));
  inv1  gate2669(.a(G552), .O(gate174inter8));
  nand2 gate2670(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate2671(.a(s_303), .b(gate174inter3), .O(gate174inter10));
  nor2  gate2672(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate2673(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate2674(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );

  xor2  gate603(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate604(.a(gate177inter0), .b(s_8), .O(gate177inter1));
  and2  gate605(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate606(.a(s_8), .O(gate177inter3));
  inv1  gate607(.a(s_9), .O(gate177inter4));
  nand2 gate608(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate609(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate610(.a(G498), .O(gate177inter7));
  inv1  gate611(.a(G558), .O(gate177inter8));
  nand2 gate612(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate613(.a(s_9), .b(gate177inter3), .O(gate177inter10));
  nor2  gate614(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate615(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate616(.a(gate177inter12), .b(gate177inter1), .O(G594));
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate1583(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate1584(.a(gate181inter0), .b(s_148), .O(gate181inter1));
  and2  gate1585(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate1586(.a(s_148), .O(gate181inter3));
  inv1  gate1587(.a(s_149), .O(gate181inter4));
  nand2 gate1588(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate1589(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate1590(.a(G510), .O(gate181inter7));
  inv1  gate1591(.a(G564), .O(gate181inter8));
  nand2 gate1592(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate1593(.a(s_149), .b(gate181inter3), .O(gate181inter10));
  nor2  gate1594(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate1595(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate1596(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate2311(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate2312(.a(gate188inter0), .b(s_252), .O(gate188inter1));
  and2  gate2313(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate2314(.a(s_252), .O(gate188inter3));
  inv1  gate2315(.a(s_253), .O(gate188inter4));
  nand2 gate2316(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate2317(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate2318(.a(G576), .O(gate188inter7));
  inv1  gate2319(.a(G577), .O(gate188inter8));
  nand2 gate2320(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate2321(.a(s_253), .b(gate188inter3), .O(gate188inter10));
  nor2  gate2322(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate2323(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate2324(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate547(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate548(.a(gate191inter0), .b(s_0), .O(gate191inter1));
  and2  gate549(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate550(.a(s_0), .O(gate191inter3));
  inv1  gate551(.a(s_1), .O(gate191inter4));
  nand2 gate552(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate553(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate554(.a(G582), .O(gate191inter7));
  inv1  gate555(.a(G583), .O(gate191inter8));
  nand2 gate556(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate557(.a(s_1), .b(gate191inter3), .O(gate191inter10));
  nor2  gate558(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate559(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate560(.a(gate191inter12), .b(gate191inter1), .O(G632));

  xor2  gate2717(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate2718(.a(gate192inter0), .b(s_310), .O(gate192inter1));
  and2  gate2719(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate2720(.a(s_310), .O(gate192inter3));
  inv1  gate2721(.a(s_311), .O(gate192inter4));
  nand2 gate2722(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate2723(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate2724(.a(G584), .O(gate192inter7));
  inv1  gate2725(.a(G585), .O(gate192inter8));
  nand2 gate2726(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate2727(.a(s_311), .b(gate192inter3), .O(gate192inter10));
  nor2  gate2728(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate2729(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate2730(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate575(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate576(.a(gate197inter0), .b(s_4), .O(gate197inter1));
  and2  gate577(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate578(.a(s_4), .O(gate197inter3));
  inv1  gate579(.a(s_5), .O(gate197inter4));
  nand2 gate580(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate581(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate582(.a(G594), .O(gate197inter7));
  inv1  gate583(.a(G595), .O(gate197inter8));
  nand2 gate584(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate585(.a(s_5), .b(gate197inter3), .O(gate197inter10));
  nor2  gate586(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate587(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate588(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );

  xor2  gate743(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate744(.a(gate202inter0), .b(s_28), .O(gate202inter1));
  and2  gate745(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate746(.a(s_28), .O(gate202inter3));
  inv1  gate747(.a(s_29), .O(gate202inter4));
  nand2 gate748(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate749(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate750(.a(G612), .O(gate202inter7));
  inv1  gate751(.a(G617), .O(gate202inter8));
  nand2 gate752(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate753(.a(s_29), .b(gate202inter3), .O(gate202inter10));
  nor2  gate754(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate755(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate756(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );

  xor2  gate1149(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate1150(.a(gate204inter0), .b(s_86), .O(gate204inter1));
  and2  gate1151(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate1152(.a(s_86), .O(gate204inter3));
  inv1  gate1153(.a(s_87), .O(gate204inter4));
  nand2 gate1154(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate1155(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate1156(.a(G607), .O(gate204inter7));
  inv1  gate1157(.a(G617), .O(gate204inter8));
  nand2 gate1158(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate1159(.a(s_87), .b(gate204inter3), .O(gate204inter10));
  nor2  gate1160(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate1161(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate1162(.a(gate204inter12), .b(gate204inter1), .O(G675));
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );

  xor2  gate2675(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate2676(.a(gate208inter0), .b(s_304), .O(gate208inter1));
  and2  gate2677(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate2678(.a(s_304), .O(gate208inter3));
  inv1  gate2679(.a(s_305), .O(gate208inter4));
  nand2 gate2680(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate2681(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate2682(.a(G627), .O(gate208inter7));
  inv1  gate2683(.a(G637), .O(gate208inter8));
  nand2 gate2684(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate2685(.a(s_305), .b(gate208inter3), .O(gate208inter10));
  nor2  gate2686(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate2687(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate2688(.a(gate208inter12), .b(gate208inter1), .O(G687));

  xor2  gate1835(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate1836(.a(gate209inter0), .b(s_184), .O(gate209inter1));
  and2  gate1837(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate1838(.a(s_184), .O(gate209inter3));
  inv1  gate1839(.a(s_185), .O(gate209inter4));
  nand2 gate1840(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate1841(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate1842(.a(G602), .O(gate209inter7));
  inv1  gate1843(.a(G666), .O(gate209inter8));
  nand2 gate1844(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate1845(.a(s_185), .b(gate209inter3), .O(gate209inter10));
  nor2  gate1846(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate1847(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate1848(.a(gate209inter12), .b(gate209inter1), .O(G690));

  xor2  gate911(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate912(.a(gate210inter0), .b(s_52), .O(gate210inter1));
  and2  gate913(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate914(.a(s_52), .O(gate210inter3));
  inv1  gate915(.a(s_53), .O(gate210inter4));
  nand2 gate916(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate917(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate918(.a(G607), .O(gate210inter7));
  inv1  gate919(.a(G666), .O(gate210inter8));
  nand2 gate920(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate921(.a(s_53), .b(gate210inter3), .O(gate210inter10));
  nor2  gate922(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate923(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate924(.a(gate210inter12), .b(gate210inter1), .O(G691));
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate2647(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate2648(.a(gate214inter0), .b(s_300), .O(gate214inter1));
  and2  gate2649(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate2650(.a(s_300), .O(gate214inter3));
  inv1  gate2651(.a(s_301), .O(gate214inter4));
  nand2 gate2652(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate2653(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate2654(.a(G612), .O(gate214inter7));
  inv1  gate2655(.a(G672), .O(gate214inter8));
  nand2 gate2656(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate2657(.a(s_301), .b(gate214inter3), .O(gate214inter10));
  nor2  gate2658(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate2659(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate2660(.a(gate214inter12), .b(gate214inter1), .O(G695));

  xor2  gate1751(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate1752(.a(gate215inter0), .b(s_172), .O(gate215inter1));
  and2  gate1753(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate1754(.a(s_172), .O(gate215inter3));
  inv1  gate1755(.a(s_173), .O(gate215inter4));
  nand2 gate1756(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate1757(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate1758(.a(G607), .O(gate215inter7));
  inv1  gate1759(.a(G675), .O(gate215inter8));
  nand2 gate1760(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate1761(.a(s_173), .b(gate215inter3), .O(gate215inter10));
  nor2  gate1762(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate1763(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate1764(.a(gate215inter12), .b(gate215inter1), .O(G696));

  xor2  gate1485(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate1486(.a(gate216inter0), .b(s_134), .O(gate216inter1));
  and2  gate1487(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate1488(.a(s_134), .O(gate216inter3));
  inv1  gate1489(.a(s_135), .O(gate216inter4));
  nand2 gate1490(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate1491(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate1492(.a(G617), .O(gate216inter7));
  inv1  gate1493(.a(G675), .O(gate216inter8));
  nand2 gate1494(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate1495(.a(s_135), .b(gate216inter3), .O(gate216inter10));
  nor2  gate1496(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate1497(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate1498(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate589(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate590(.a(gate218inter0), .b(s_6), .O(gate218inter1));
  and2  gate591(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate592(.a(s_6), .O(gate218inter3));
  inv1  gate593(.a(s_7), .O(gate218inter4));
  nand2 gate594(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate595(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate596(.a(G627), .O(gate218inter7));
  inv1  gate597(.a(G678), .O(gate218inter8));
  nand2 gate598(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate599(.a(s_7), .b(gate218inter3), .O(gate218inter10));
  nor2  gate600(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate601(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate602(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate1989(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate1990(.a(gate220inter0), .b(s_206), .O(gate220inter1));
  and2  gate1991(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate1992(.a(s_206), .O(gate220inter3));
  inv1  gate1993(.a(s_207), .O(gate220inter4));
  nand2 gate1994(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate1995(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate1996(.a(G637), .O(gate220inter7));
  inv1  gate1997(.a(G681), .O(gate220inter8));
  nand2 gate1998(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate1999(.a(s_207), .b(gate220inter3), .O(gate220inter10));
  nor2  gate2000(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate2001(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate2002(.a(gate220inter12), .b(gate220inter1), .O(G701));
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate785(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate786(.a(gate224inter0), .b(s_34), .O(gate224inter1));
  and2  gate787(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate788(.a(s_34), .O(gate224inter3));
  inv1  gate789(.a(s_35), .O(gate224inter4));
  nand2 gate790(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate791(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate792(.a(G637), .O(gate224inter7));
  inv1  gate793(.a(G687), .O(gate224inter8));
  nand2 gate794(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate795(.a(s_35), .b(gate224inter3), .O(gate224inter10));
  nor2  gate796(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate797(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate798(.a(gate224inter12), .b(gate224inter1), .O(G705));

  xor2  gate897(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate898(.a(gate225inter0), .b(s_50), .O(gate225inter1));
  and2  gate899(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate900(.a(s_50), .O(gate225inter3));
  inv1  gate901(.a(s_51), .O(gate225inter4));
  nand2 gate902(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate903(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate904(.a(G690), .O(gate225inter7));
  inv1  gate905(.a(G691), .O(gate225inter8));
  nand2 gate906(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate907(.a(s_51), .b(gate225inter3), .O(gate225inter10));
  nor2  gate908(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate909(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate910(.a(gate225inter12), .b(gate225inter1), .O(G706));
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate2381(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate2382(.a(gate228inter0), .b(s_262), .O(gate228inter1));
  and2  gate2383(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate2384(.a(s_262), .O(gate228inter3));
  inv1  gate2385(.a(s_263), .O(gate228inter4));
  nand2 gate2386(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate2387(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate2388(.a(G696), .O(gate228inter7));
  inv1  gate2389(.a(G697), .O(gate228inter8));
  nand2 gate2390(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate2391(.a(s_263), .b(gate228inter3), .O(gate228inter10));
  nor2  gate2392(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate2393(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate2394(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate1065(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate1066(.a(gate231inter0), .b(s_74), .O(gate231inter1));
  and2  gate1067(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate1068(.a(s_74), .O(gate231inter3));
  inv1  gate1069(.a(s_75), .O(gate231inter4));
  nand2 gate1070(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate1071(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate1072(.a(G702), .O(gate231inter7));
  inv1  gate1073(.a(G703), .O(gate231inter8));
  nand2 gate1074(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate1075(.a(s_75), .b(gate231inter3), .O(gate231inter10));
  nor2  gate1076(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate1077(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate1078(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate1177(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate1178(.a(gate233inter0), .b(s_90), .O(gate233inter1));
  and2  gate1179(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate1180(.a(s_90), .O(gate233inter3));
  inv1  gate1181(.a(s_91), .O(gate233inter4));
  nand2 gate1182(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1183(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1184(.a(G242), .O(gate233inter7));
  inv1  gate1185(.a(G718), .O(gate233inter8));
  nand2 gate1186(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1187(.a(s_91), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1188(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1189(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1190(.a(gate233inter12), .b(gate233inter1), .O(G730));

  xor2  gate2563(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate2564(.a(gate234inter0), .b(s_288), .O(gate234inter1));
  and2  gate2565(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate2566(.a(s_288), .O(gate234inter3));
  inv1  gate2567(.a(s_289), .O(gate234inter4));
  nand2 gate2568(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate2569(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate2570(.a(G245), .O(gate234inter7));
  inv1  gate2571(.a(G721), .O(gate234inter8));
  nand2 gate2572(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate2573(.a(s_289), .b(gate234inter3), .O(gate234inter10));
  nor2  gate2574(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate2575(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate2576(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate1121(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate1122(.a(gate237inter0), .b(s_82), .O(gate237inter1));
  and2  gate1123(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate1124(.a(s_82), .O(gate237inter3));
  inv1  gate1125(.a(s_83), .O(gate237inter4));
  nand2 gate1126(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1127(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1128(.a(G254), .O(gate237inter7));
  inv1  gate1129(.a(G706), .O(gate237inter8));
  nand2 gate1130(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1131(.a(s_83), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1132(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1133(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1134(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate827(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate828(.a(gate249inter0), .b(s_40), .O(gate249inter1));
  and2  gate829(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate830(.a(s_40), .O(gate249inter3));
  inv1  gate831(.a(s_41), .O(gate249inter4));
  nand2 gate832(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate833(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate834(.a(G254), .O(gate249inter7));
  inv1  gate835(.a(G742), .O(gate249inter8));
  nand2 gate836(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate837(.a(s_41), .b(gate249inter3), .O(gate249inter10));
  nor2  gate838(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate839(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate840(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate2031(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate2032(.a(gate255inter0), .b(s_212), .O(gate255inter1));
  and2  gate2033(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate2034(.a(s_212), .O(gate255inter3));
  inv1  gate2035(.a(s_213), .O(gate255inter4));
  nand2 gate2036(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate2037(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate2038(.a(G263), .O(gate255inter7));
  inv1  gate2039(.a(G751), .O(gate255inter8));
  nand2 gate2040(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate2041(.a(s_213), .b(gate255inter3), .O(gate255inter10));
  nor2  gate2042(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate2043(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate2044(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );

  xor2  gate1569(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate1570(.a(gate259inter0), .b(s_146), .O(gate259inter1));
  and2  gate1571(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate1572(.a(s_146), .O(gate259inter3));
  inv1  gate1573(.a(s_147), .O(gate259inter4));
  nand2 gate1574(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate1575(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate1576(.a(G758), .O(gate259inter7));
  inv1  gate1577(.a(G759), .O(gate259inter8));
  nand2 gate1578(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate1579(.a(s_147), .b(gate259inter3), .O(gate259inter10));
  nor2  gate1580(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate1581(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate1582(.a(gate259inter12), .b(gate259inter1), .O(G776));
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate715(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate716(.a(gate262inter0), .b(s_24), .O(gate262inter1));
  and2  gate717(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate718(.a(s_24), .O(gate262inter3));
  inv1  gate719(.a(s_25), .O(gate262inter4));
  nand2 gate720(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate721(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate722(.a(G764), .O(gate262inter7));
  inv1  gate723(.a(G765), .O(gate262inter8));
  nand2 gate724(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate725(.a(s_25), .b(gate262inter3), .O(gate262inter10));
  nor2  gate726(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate727(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate728(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate953(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate954(.a(gate265inter0), .b(s_58), .O(gate265inter1));
  and2  gate955(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate956(.a(s_58), .O(gate265inter3));
  inv1  gate957(.a(s_59), .O(gate265inter4));
  nand2 gate958(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate959(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate960(.a(G642), .O(gate265inter7));
  inv1  gate961(.a(G770), .O(gate265inter8));
  nand2 gate962(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate963(.a(s_59), .b(gate265inter3), .O(gate265inter10));
  nor2  gate964(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate965(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate966(.a(gate265inter12), .b(gate265inter1), .O(G794));

  xor2  gate2185(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate2186(.a(gate266inter0), .b(s_234), .O(gate266inter1));
  and2  gate2187(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate2188(.a(s_234), .O(gate266inter3));
  inv1  gate2189(.a(s_235), .O(gate266inter4));
  nand2 gate2190(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate2191(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate2192(.a(G645), .O(gate266inter7));
  inv1  gate2193(.a(G773), .O(gate266inter8));
  nand2 gate2194(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate2195(.a(s_235), .b(gate266inter3), .O(gate266inter10));
  nor2  gate2196(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate2197(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate2198(.a(gate266inter12), .b(gate266inter1), .O(G797));

  xor2  gate1345(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate1346(.a(gate267inter0), .b(s_114), .O(gate267inter1));
  and2  gate1347(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate1348(.a(s_114), .O(gate267inter3));
  inv1  gate1349(.a(s_115), .O(gate267inter4));
  nand2 gate1350(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate1351(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate1352(.a(G648), .O(gate267inter7));
  inv1  gate1353(.a(G776), .O(gate267inter8));
  nand2 gate1354(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate1355(.a(s_115), .b(gate267inter3), .O(gate267inter10));
  nor2  gate1356(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate1357(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate1358(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );

  xor2  gate1205(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate1206(.a(gate275inter0), .b(s_94), .O(gate275inter1));
  and2  gate1207(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate1208(.a(s_94), .O(gate275inter3));
  inv1  gate1209(.a(s_95), .O(gate275inter4));
  nand2 gate1210(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate1211(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate1212(.a(G645), .O(gate275inter7));
  inv1  gate1213(.a(G797), .O(gate275inter8));
  nand2 gate1214(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate1215(.a(s_95), .b(gate275inter3), .O(gate275inter10));
  nor2  gate1216(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate1217(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate1218(.a(gate275inter12), .b(gate275inter1), .O(G820));
nand2 gate276( .a(G773), .b(G797), .O(G821) );

  xor2  gate687(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate688(.a(gate277inter0), .b(s_20), .O(gate277inter1));
  and2  gate689(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate690(.a(s_20), .O(gate277inter3));
  inv1  gate691(.a(s_21), .O(gate277inter4));
  nand2 gate692(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate693(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate694(.a(G648), .O(gate277inter7));
  inv1  gate695(.a(G800), .O(gate277inter8));
  nand2 gate696(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate697(.a(s_21), .b(gate277inter3), .O(gate277inter10));
  nor2  gate698(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate699(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate700(.a(gate277inter12), .b(gate277inter1), .O(G822));

  xor2  gate1107(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate1108(.a(gate278inter0), .b(s_80), .O(gate278inter1));
  and2  gate1109(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate1110(.a(s_80), .O(gate278inter3));
  inv1  gate1111(.a(s_81), .O(gate278inter4));
  nand2 gate1112(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate1113(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate1114(.a(G776), .O(gate278inter7));
  inv1  gate1115(.a(G800), .O(gate278inter8));
  nand2 gate1116(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate1117(.a(s_81), .b(gate278inter3), .O(gate278inter10));
  nor2  gate1118(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate1119(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate1120(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );

  xor2  gate1765(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate1766(.a(gate284inter0), .b(s_174), .O(gate284inter1));
  and2  gate1767(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate1768(.a(s_174), .O(gate284inter3));
  inv1  gate1769(.a(s_175), .O(gate284inter4));
  nand2 gate1770(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate1771(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate1772(.a(G785), .O(gate284inter7));
  inv1  gate1773(.a(G809), .O(gate284inter8));
  nand2 gate1774(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate1775(.a(s_175), .b(gate284inter3), .O(gate284inter10));
  nor2  gate1776(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate1777(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate1778(.a(gate284inter12), .b(gate284inter1), .O(G829));

  xor2  gate2437(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate2438(.a(gate285inter0), .b(s_270), .O(gate285inter1));
  and2  gate2439(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate2440(.a(s_270), .O(gate285inter3));
  inv1  gate2441(.a(s_271), .O(gate285inter4));
  nand2 gate2442(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate2443(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate2444(.a(G660), .O(gate285inter7));
  inv1  gate2445(.a(G812), .O(gate285inter8));
  nand2 gate2446(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate2447(.a(s_271), .b(gate285inter3), .O(gate285inter10));
  nor2  gate2448(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate2449(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate2450(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate1723(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate1724(.a(gate287inter0), .b(s_168), .O(gate287inter1));
  and2  gate1725(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate1726(.a(s_168), .O(gate287inter3));
  inv1  gate1727(.a(s_169), .O(gate287inter4));
  nand2 gate1728(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate1729(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate1730(.a(G663), .O(gate287inter7));
  inv1  gate1731(.a(G815), .O(gate287inter8));
  nand2 gate1732(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate1733(.a(s_169), .b(gate287inter3), .O(gate287inter10));
  nor2  gate1734(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate1735(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate1736(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate2409(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate2410(.a(gate289inter0), .b(s_266), .O(gate289inter1));
  and2  gate2411(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate2412(.a(s_266), .O(gate289inter3));
  inv1  gate2413(.a(s_267), .O(gate289inter4));
  nand2 gate2414(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate2415(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate2416(.a(G818), .O(gate289inter7));
  inv1  gate2417(.a(G819), .O(gate289inter8));
  nand2 gate2418(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate2419(.a(s_267), .b(gate289inter3), .O(gate289inter10));
  nor2  gate2420(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate2421(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate2422(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate1877(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate1878(.a(gate292inter0), .b(s_190), .O(gate292inter1));
  and2  gate1879(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate1880(.a(s_190), .O(gate292inter3));
  inv1  gate1881(.a(s_191), .O(gate292inter4));
  nand2 gate1882(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate1883(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate1884(.a(G824), .O(gate292inter7));
  inv1  gate1885(.a(G825), .O(gate292inter8));
  nand2 gate1886(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate1887(.a(s_191), .b(gate292inter3), .O(gate292inter10));
  nor2  gate1888(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate1889(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate1890(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate1275(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate1276(.a(gate295inter0), .b(s_104), .O(gate295inter1));
  and2  gate1277(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate1278(.a(s_104), .O(gate295inter3));
  inv1  gate1279(.a(s_105), .O(gate295inter4));
  nand2 gate1280(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate1281(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate1282(.a(G830), .O(gate295inter7));
  inv1  gate1283(.a(G831), .O(gate295inter8));
  nand2 gate1284(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate1285(.a(s_105), .b(gate295inter3), .O(gate295inter10));
  nor2  gate1286(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate1287(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate1288(.a(gate295inter12), .b(gate295inter1), .O(G912));
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate1681(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate1682(.a(gate393inter0), .b(s_162), .O(gate393inter1));
  and2  gate1683(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate1684(.a(s_162), .O(gate393inter3));
  inv1  gate1685(.a(s_163), .O(gate393inter4));
  nand2 gate1686(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate1687(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate1688(.a(G7), .O(gate393inter7));
  inv1  gate1689(.a(G1054), .O(gate393inter8));
  nand2 gate1690(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate1691(.a(s_163), .b(gate393inter3), .O(gate393inter10));
  nor2  gate1692(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate1693(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate1694(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate2479(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate2480(.a(gate395inter0), .b(s_276), .O(gate395inter1));
  and2  gate2481(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate2482(.a(s_276), .O(gate395inter3));
  inv1  gate2483(.a(s_277), .O(gate395inter4));
  nand2 gate2484(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate2485(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate2486(.a(G9), .O(gate395inter7));
  inv1  gate2487(.a(G1060), .O(gate395inter8));
  nand2 gate2488(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate2489(.a(s_277), .b(gate395inter3), .O(gate395inter10));
  nor2  gate2490(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate2491(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate2492(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate631(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate632(.a(gate397inter0), .b(s_12), .O(gate397inter1));
  and2  gate633(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate634(.a(s_12), .O(gate397inter3));
  inv1  gate635(.a(s_13), .O(gate397inter4));
  nand2 gate636(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate637(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate638(.a(G11), .O(gate397inter7));
  inv1  gate639(.a(G1066), .O(gate397inter8));
  nand2 gate640(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate641(.a(s_13), .b(gate397inter3), .O(gate397inter10));
  nor2  gate642(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate643(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate644(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate1947(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate1948(.a(gate399inter0), .b(s_200), .O(gate399inter1));
  and2  gate1949(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate1950(.a(s_200), .O(gate399inter3));
  inv1  gate1951(.a(s_201), .O(gate399inter4));
  nand2 gate1952(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate1953(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate1954(.a(G13), .O(gate399inter7));
  inv1  gate1955(.a(G1072), .O(gate399inter8));
  nand2 gate1956(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate1957(.a(s_201), .b(gate399inter3), .O(gate399inter10));
  nor2  gate1958(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate1959(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate1960(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );

  xor2  gate2115(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate2116(.a(gate401inter0), .b(s_224), .O(gate401inter1));
  and2  gate2117(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate2118(.a(s_224), .O(gate401inter3));
  inv1  gate2119(.a(s_225), .O(gate401inter4));
  nand2 gate2120(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate2121(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate2122(.a(G15), .O(gate401inter7));
  inv1  gate2123(.a(G1078), .O(gate401inter8));
  nand2 gate2124(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate2125(.a(s_225), .b(gate401inter3), .O(gate401inter10));
  nor2  gate2126(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate2127(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate2128(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );

  xor2  gate2451(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate2452(.a(gate405inter0), .b(s_272), .O(gate405inter1));
  and2  gate2453(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate2454(.a(s_272), .O(gate405inter3));
  inv1  gate2455(.a(s_273), .O(gate405inter4));
  nand2 gate2456(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate2457(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate2458(.a(G19), .O(gate405inter7));
  inv1  gate2459(.a(G1090), .O(gate405inter8));
  nand2 gate2460(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate2461(.a(s_273), .b(gate405inter3), .O(gate405inter10));
  nor2  gate2462(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate2463(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate2464(.a(gate405inter12), .b(gate405inter1), .O(G1186));

  xor2  gate2633(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate2634(.a(gate406inter0), .b(s_298), .O(gate406inter1));
  and2  gate2635(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate2636(.a(s_298), .O(gate406inter3));
  inv1  gate2637(.a(s_299), .O(gate406inter4));
  nand2 gate2638(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate2639(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate2640(.a(G20), .O(gate406inter7));
  inv1  gate2641(.a(G1093), .O(gate406inter8));
  nand2 gate2642(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate2643(.a(s_299), .b(gate406inter3), .O(gate406inter10));
  nor2  gate2644(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate2645(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate2646(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate729(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate730(.a(gate410inter0), .b(s_26), .O(gate410inter1));
  and2  gate731(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate732(.a(s_26), .O(gate410inter3));
  inv1  gate733(.a(s_27), .O(gate410inter4));
  nand2 gate734(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate735(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate736(.a(G24), .O(gate410inter7));
  inv1  gate737(.a(G1105), .O(gate410inter8));
  nand2 gate738(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate739(.a(s_27), .b(gate410inter3), .O(gate410inter10));
  nor2  gate740(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate741(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate742(.a(gate410inter12), .b(gate410inter1), .O(G1201));

  xor2  gate1933(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate1934(.a(gate411inter0), .b(s_198), .O(gate411inter1));
  and2  gate1935(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate1936(.a(s_198), .O(gate411inter3));
  inv1  gate1937(.a(s_199), .O(gate411inter4));
  nand2 gate1938(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate1939(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate1940(.a(G25), .O(gate411inter7));
  inv1  gate1941(.a(G1108), .O(gate411inter8));
  nand2 gate1942(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate1943(.a(s_199), .b(gate411inter3), .O(gate411inter10));
  nor2  gate1944(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate1945(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate1946(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate1737(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate1738(.a(gate413inter0), .b(s_170), .O(gate413inter1));
  and2  gate1739(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate1740(.a(s_170), .O(gate413inter3));
  inv1  gate1741(.a(s_171), .O(gate413inter4));
  nand2 gate1742(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1743(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1744(.a(G27), .O(gate413inter7));
  inv1  gate1745(.a(G1114), .O(gate413inter8));
  nand2 gate1746(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1747(.a(s_171), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1748(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1749(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1750(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate1443(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate1444(.a(gate417inter0), .b(s_128), .O(gate417inter1));
  and2  gate1445(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate1446(.a(s_128), .O(gate417inter3));
  inv1  gate1447(.a(s_129), .O(gate417inter4));
  nand2 gate1448(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate1449(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate1450(.a(G31), .O(gate417inter7));
  inv1  gate1451(.a(G1126), .O(gate417inter8));
  nand2 gate1452(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate1453(.a(s_129), .b(gate417inter3), .O(gate417inter10));
  nor2  gate1454(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate1455(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate1456(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate757(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate758(.a(gate419inter0), .b(s_30), .O(gate419inter1));
  and2  gate759(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate760(.a(s_30), .O(gate419inter3));
  inv1  gate761(.a(s_31), .O(gate419inter4));
  nand2 gate762(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate763(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate764(.a(G1), .O(gate419inter7));
  inv1  gate765(.a(G1132), .O(gate419inter8));
  nand2 gate766(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate767(.a(s_31), .b(gate419inter3), .O(gate419inter10));
  nor2  gate768(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate769(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate770(.a(gate419inter12), .b(gate419inter1), .O(G1228));
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate2591(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate2592(.a(gate425inter0), .b(s_292), .O(gate425inter1));
  and2  gate2593(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate2594(.a(s_292), .O(gate425inter3));
  inv1  gate2595(.a(s_293), .O(gate425inter4));
  nand2 gate2596(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate2597(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate2598(.a(G4), .O(gate425inter7));
  inv1  gate2599(.a(G1141), .O(gate425inter8));
  nand2 gate2600(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate2601(.a(s_293), .b(gate425inter3), .O(gate425inter10));
  nor2  gate2602(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate2603(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate2604(.a(gate425inter12), .b(gate425inter1), .O(G1234));

  xor2  gate2423(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate2424(.a(gate426inter0), .b(s_268), .O(gate426inter1));
  and2  gate2425(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate2426(.a(s_268), .O(gate426inter3));
  inv1  gate2427(.a(s_269), .O(gate426inter4));
  nand2 gate2428(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate2429(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate2430(.a(G1045), .O(gate426inter7));
  inv1  gate2431(.a(G1141), .O(gate426inter8));
  nand2 gate2432(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate2433(.a(s_269), .b(gate426inter3), .O(gate426inter10));
  nor2  gate2434(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate2435(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate2436(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate2045(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate2046(.a(gate428inter0), .b(s_214), .O(gate428inter1));
  and2  gate2047(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate2048(.a(s_214), .O(gate428inter3));
  inv1  gate2049(.a(s_215), .O(gate428inter4));
  nand2 gate2050(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate2051(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate2052(.a(G1048), .O(gate428inter7));
  inv1  gate2053(.a(G1144), .O(gate428inter8));
  nand2 gate2054(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate2055(.a(s_215), .b(gate428inter3), .O(gate428inter10));
  nor2  gate2056(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate2057(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate2058(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate1695(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate1696(.a(gate430inter0), .b(s_164), .O(gate430inter1));
  and2  gate1697(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate1698(.a(s_164), .O(gate430inter3));
  inv1  gate1699(.a(s_165), .O(gate430inter4));
  nand2 gate1700(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate1701(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate1702(.a(G1051), .O(gate430inter7));
  inv1  gate1703(.a(G1147), .O(gate430inter8));
  nand2 gate1704(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate1705(.a(s_165), .b(gate430inter3), .O(gate430inter10));
  nor2  gate1706(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate1707(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate1708(.a(gate430inter12), .b(gate430inter1), .O(G1239));

  xor2  gate1863(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate1864(.a(gate431inter0), .b(s_188), .O(gate431inter1));
  and2  gate1865(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate1866(.a(s_188), .O(gate431inter3));
  inv1  gate1867(.a(s_189), .O(gate431inter4));
  nand2 gate1868(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate1869(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate1870(.a(G7), .O(gate431inter7));
  inv1  gate1871(.a(G1150), .O(gate431inter8));
  nand2 gate1872(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate1873(.a(s_189), .b(gate431inter3), .O(gate431inter10));
  nor2  gate1874(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate1875(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate1876(.a(gate431inter12), .b(gate431inter1), .O(G1240));

  xor2  gate1779(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate1780(.a(gate432inter0), .b(s_176), .O(gate432inter1));
  and2  gate1781(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate1782(.a(s_176), .O(gate432inter3));
  inv1  gate1783(.a(s_177), .O(gate432inter4));
  nand2 gate1784(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate1785(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate1786(.a(G1054), .O(gate432inter7));
  inv1  gate1787(.a(G1150), .O(gate432inter8));
  nand2 gate1788(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate1789(.a(s_177), .b(gate432inter3), .O(gate432inter10));
  nor2  gate1790(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate1791(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate1792(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate1233(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate1234(.a(gate434inter0), .b(s_98), .O(gate434inter1));
  and2  gate1235(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate1236(.a(s_98), .O(gate434inter3));
  inv1  gate1237(.a(s_99), .O(gate434inter4));
  nand2 gate1238(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate1239(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate1240(.a(G1057), .O(gate434inter7));
  inv1  gate1241(.a(G1153), .O(gate434inter8));
  nand2 gate1242(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate1243(.a(s_99), .b(gate434inter3), .O(gate434inter10));
  nor2  gate1244(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate1245(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate1246(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate2493(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate2494(.a(gate438inter0), .b(s_278), .O(gate438inter1));
  and2  gate2495(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate2496(.a(s_278), .O(gate438inter3));
  inv1  gate2497(.a(s_279), .O(gate438inter4));
  nand2 gate2498(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate2499(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate2500(.a(G1063), .O(gate438inter7));
  inv1  gate2501(.a(G1159), .O(gate438inter8));
  nand2 gate2502(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate2503(.a(s_279), .b(gate438inter3), .O(gate438inter10));
  nor2  gate2504(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate2505(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate2506(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate1247(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate1248(.a(gate443inter0), .b(s_100), .O(gate443inter1));
  and2  gate1249(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate1250(.a(s_100), .O(gate443inter3));
  inv1  gate1251(.a(s_101), .O(gate443inter4));
  nand2 gate1252(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate1253(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate1254(.a(G13), .O(gate443inter7));
  inv1  gate1255(.a(G1168), .O(gate443inter8));
  nand2 gate1256(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate1257(.a(s_101), .b(gate443inter3), .O(gate443inter10));
  nor2  gate1258(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate1259(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate1260(.a(gate443inter12), .b(gate443inter1), .O(G1252));

  xor2  gate2507(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate2508(.a(gate444inter0), .b(s_280), .O(gate444inter1));
  and2  gate2509(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate2510(.a(s_280), .O(gate444inter3));
  inv1  gate2511(.a(s_281), .O(gate444inter4));
  nand2 gate2512(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate2513(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate2514(.a(G1072), .O(gate444inter7));
  inv1  gate2515(.a(G1168), .O(gate444inter8));
  nand2 gate2516(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate2517(.a(s_281), .b(gate444inter3), .O(gate444inter10));
  nor2  gate2518(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate2519(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate2520(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );

  xor2  gate2241(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate2242(.a(gate447inter0), .b(s_242), .O(gate447inter1));
  and2  gate2243(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate2244(.a(s_242), .O(gate447inter3));
  inv1  gate2245(.a(s_243), .O(gate447inter4));
  nand2 gate2246(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate2247(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate2248(.a(G15), .O(gate447inter7));
  inv1  gate2249(.a(G1174), .O(gate447inter8));
  nand2 gate2250(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate2251(.a(s_243), .b(gate447inter3), .O(gate447inter10));
  nor2  gate2252(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate2253(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate2254(.a(gate447inter12), .b(gate447inter1), .O(G1256));
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );

  xor2  gate1555(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate1556(.a(gate451inter0), .b(s_144), .O(gate451inter1));
  and2  gate1557(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate1558(.a(s_144), .O(gate451inter3));
  inv1  gate1559(.a(s_145), .O(gate451inter4));
  nand2 gate1560(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate1561(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate1562(.a(G17), .O(gate451inter7));
  inv1  gate1563(.a(G1180), .O(gate451inter8));
  nand2 gate1564(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate1565(.a(s_145), .b(gate451inter3), .O(gate451inter10));
  nor2  gate1566(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate1567(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate1568(.a(gate451inter12), .b(gate451inter1), .O(G1260));
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );

  xor2  gate2213(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate2214(.a(gate455inter0), .b(s_238), .O(gate455inter1));
  and2  gate2215(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate2216(.a(s_238), .O(gate455inter3));
  inv1  gate2217(.a(s_239), .O(gate455inter4));
  nand2 gate2218(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate2219(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate2220(.a(G19), .O(gate455inter7));
  inv1  gate2221(.a(G1186), .O(gate455inter8));
  nand2 gate2222(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate2223(.a(s_239), .b(gate455inter3), .O(gate455inter10));
  nor2  gate2224(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate2225(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate2226(.a(gate455inter12), .b(gate455inter1), .O(G1264));

  xor2  gate1639(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate1640(.a(gate456inter0), .b(s_156), .O(gate456inter1));
  and2  gate1641(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate1642(.a(s_156), .O(gate456inter3));
  inv1  gate1643(.a(s_157), .O(gate456inter4));
  nand2 gate1644(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate1645(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate1646(.a(G1090), .O(gate456inter7));
  inv1  gate1647(.a(G1186), .O(gate456inter8));
  nand2 gate1648(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate1649(.a(s_157), .b(gate456inter3), .O(gate456inter10));
  nor2  gate1650(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate1651(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate1652(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate841(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate842(.a(gate459inter0), .b(s_42), .O(gate459inter1));
  and2  gate843(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate844(.a(s_42), .O(gate459inter3));
  inv1  gate845(.a(s_43), .O(gate459inter4));
  nand2 gate846(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate847(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate848(.a(G21), .O(gate459inter7));
  inv1  gate849(.a(G1192), .O(gate459inter8));
  nand2 gate850(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate851(.a(s_43), .b(gate459inter3), .O(gate459inter10));
  nor2  gate852(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate853(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate854(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate1975(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate1976(.a(gate463inter0), .b(s_204), .O(gate463inter1));
  and2  gate1977(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate1978(.a(s_204), .O(gate463inter3));
  inv1  gate1979(.a(s_205), .O(gate463inter4));
  nand2 gate1980(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate1981(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate1982(.a(G23), .O(gate463inter7));
  inv1  gate1983(.a(G1198), .O(gate463inter8));
  nand2 gate1984(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate1985(.a(s_205), .b(gate463inter3), .O(gate463inter10));
  nor2  gate1986(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate1987(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate1988(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate1457(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate1458(.a(gate467inter0), .b(s_130), .O(gate467inter1));
  and2  gate1459(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate1460(.a(s_130), .O(gate467inter3));
  inv1  gate1461(.a(s_131), .O(gate467inter4));
  nand2 gate1462(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate1463(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate1464(.a(G25), .O(gate467inter7));
  inv1  gate1465(.a(G1204), .O(gate467inter8));
  nand2 gate1466(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate1467(.a(s_131), .b(gate467inter3), .O(gate467inter10));
  nor2  gate1468(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate1469(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate1470(.a(gate467inter12), .b(gate467inter1), .O(G1276));

  xor2  gate1037(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate1038(.a(gate468inter0), .b(s_70), .O(gate468inter1));
  and2  gate1039(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate1040(.a(s_70), .O(gate468inter3));
  inv1  gate1041(.a(s_71), .O(gate468inter4));
  nand2 gate1042(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate1043(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate1044(.a(G1108), .O(gate468inter7));
  inv1  gate1045(.a(G1204), .O(gate468inter8));
  nand2 gate1046(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate1047(.a(s_71), .b(gate468inter3), .O(gate468inter10));
  nor2  gate1048(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate1049(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate1050(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );

  xor2  gate1051(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate1052(.a(gate470inter0), .b(s_72), .O(gate470inter1));
  and2  gate1053(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate1054(.a(s_72), .O(gate470inter3));
  inv1  gate1055(.a(s_73), .O(gate470inter4));
  nand2 gate1056(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate1057(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate1058(.a(G1111), .O(gate470inter7));
  inv1  gate1059(.a(G1207), .O(gate470inter8));
  nand2 gate1060(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate1061(.a(s_73), .b(gate470inter3), .O(gate470inter10));
  nor2  gate1062(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate1063(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate1064(.a(gate470inter12), .b(gate470inter1), .O(G1279));

  xor2  gate1289(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate1290(.a(gate471inter0), .b(s_106), .O(gate471inter1));
  and2  gate1291(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate1292(.a(s_106), .O(gate471inter3));
  inv1  gate1293(.a(s_107), .O(gate471inter4));
  nand2 gate1294(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate1295(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate1296(.a(G27), .O(gate471inter7));
  inv1  gate1297(.a(G1210), .O(gate471inter8));
  nand2 gate1298(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate1299(.a(s_107), .b(gate471inter3), .O(gate471inter10));
  nor2  gate1300(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate1301(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate1302(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate1303(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate1304(.a(gate474inter0), .b(s_108), .O(gate474inter1));
  and2  gate1305(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate1306(.a(s_108), .O(gate474inter3));
  inv1  gate1307(.a(s_109), .O(gate474inter4));
  nand2 gate1308(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate1309(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate1310(.a(G1117), .O(gate474inter7));
  inv1  gate1311(.a(G1213), .O(gate474inter8));
  nand2 gate1312(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate1313(.a(s_109), .b(gate474inter3), .O(gate474inter10));
  nor2  gate1314(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate1315(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate1316(.a(gate474inter12), .b(gate474inter1), .O(G1283));

  xor2  gate2703(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate2704(.a(gate475inter0), .b(s_308), .O(gate475inter1));
  and2  gate2705(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate2706(.a(s_308), .O(gate475inter3));
  inv1  gate2707(.a(s_309), .O(gate475inter4));
  nand2 gate2708(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate2709(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate2710(.a(G29), .O(gate475inter7));
  inv1  gate2711(.a(G1216), .O(gate475inter8));
  nand2 gate2712(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate2713(.a(s_309), .b(gate475inter3), .O(gate475inter10));
  nor2  gate2714(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate2715(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate2716(.a(gate475inter12), .b(gate475inter1), .O(G1284));

  xor2  gate1499(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate1500(.a(gate476inter0), .b(s_136), .O(gate476inter1));
  and2  gate1501(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate1502(.a(s_136), .O(gate476inter3));
  inv1  gate1503(.a(s_137), .O(gate476inter4));
  nand2 gate1504(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate1505(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate1506(.a(G1120), .O(gate476inter7));
  inv1  gate1507(.a(G1216), .O(gate476inter8));
  nand2 gate1508(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate1509(.a(s_137), .b(gate476inter3), .O(gate476inter10));
  nor2  gate1510(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate1511(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate1512(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );

  xor2  gate701(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate702(.a(gate478inter0), .b(s_22), .O(gate478inter1));
  and2  gate703(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate704(.a(s_22), .O(gate478inter3));
  inv1  gate705(.a(s_23), .O(gate478inter4));
  nand2 gate706(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate707(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate708(.a(G1123), .O(gate478inter7));
  inv1  gate709(.a(G1219), .O(gate478inter8));
  nand2 gate710(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate711(.a(s_23), .b(gate478inter3), .O(gate478inter10));
  nor2  gate712(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate713(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate714(.a(gate478inter12), .b(gate478inter1), .O(G1287));
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate1961(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate1962(.a(gate480inter0), .b(s_202), .O(gate480inter1));
  and2  gate1963(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate1964(.a(s_202), .O(gate480inter3));
  inv1  gate1965(.a(s_203), .O(gate480inter4));
  nand2 gate1966(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate1967(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate1968(.a(G1126), .O(gate480inter7));
  inv1  gate1969(.a(G1222), .O(gate480inter8));
  nand2 gate1970(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate1971(.a(s_203), .b(gate480inter3), .O(gate480inter10));
  nor2  gate1972(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate1973(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate1974(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate2283(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate2284(.a(gate482inter0), .b(s_248), .O(gate482inter1));
  and2  gate2285(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate2286(.a(s_248), .O(gate482inter3));
  inv1  gate2287(.a(s_249), .O(gate482inter4));
  nand2 gate2288(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate2289(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate2290(.a(G1129), .O(gate482inter7));
  inv1  gate2291(.a(G1225), .O(gate482inter8));
  nand2 gate2292(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate2293(.a(s_249), .b(gate482inter3), .O(gate482inter10));
  nor2  gate2294(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate2295(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate2296(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );

  xor2  gate659(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate660(.a(gate484inter0), .b(s_16), .O(gate484inter1));
  and2  gate661(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate662(.a(s_16), .O(gate484inter3));
  inv1  gate663(.a(s_17), .O(gate484inter4));
  nand2 gate664(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate665(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate666(.a(G1230), .O(gate484inter7));
  inv1  gate667(.a(G1231), .O(gate484inter8));
  nand2 gate668(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate669(.a(s_17), .b(gate484inter3), .O(gate484inter10));
  nor2  gate670(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate671(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate672(.a(gate484inter12), .b(gate484inter1), .O(G1293));
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate2689(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate2690(.a(gate488inter0), .b(s_306), .O(gate488inter1));
  and2  gate2691(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate2692(.a(s_306), .O(gate488inter3));
  inv1  gate2693(.a(s_307), .O(gate488inter4));
  nand2 gate2694(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate2695(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate2696(.a(G1238), .O(gate488inter7));
  inv1  gate2697(.a(G1239), .O(gate488inter8));
  nand2 gate2698(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate2699(.a(s_307), .b(gate488inter3), .O(gate488inter10));
  nor2  gate2700(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate2701(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate2702(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate1471(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate1472(.a(gate491inter0), .b(s_132), .O(gate491inter1));
  and2  gate1473(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate1474(.a(s_132), .O(gate491inter3));
  inv1  gate1475(.a(s_133), .O(gate491inter4));
  nand2 gate1476(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate1477(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate1478(.a(G1244), .O(gate491inter7));
  inv1  gate1479(.a(G1245), .O(gate491inter8));
  nand2 gate1480(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate1481(.a(s_133), .b(gate491inter3), .O(gate491inter10));
  nor2  gate1482(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate1483(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate1484(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate2465(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate2466(.a(gate494inter0), .b(s_274), .O(gate494inter1));
  and2  gate2467(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate2468(.a(s_274), .O(gate494inter3));
  inv1  gate2469(.a(s_275), .O(gate494inter4));
  nand2 gate2470(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate2471(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate2472(.a(G1250), .O(gate494inter7));
  inv1  gate2473(.a(G1251), .O(gate494inter8));
  nand2 gate2474(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate2475(.a(s_275), .b(gate494inter3), .O(gate494inter10));
  nor2  gate2476(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate2477(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate2478(.a(gate494inter12), .b(gate494inter1), .O(G1303));

  xor2  gate1401(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate1402(.a(gate495inter0), .b(s_122), .O(gate495inter1));
  and2  gate1403(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate1404(.a(s_122), .O(gate495inter3));
  inv1  gate1405(.a(s_123), .O(gate495inter4));
  nand2 gate1406(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate1407(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate1408(.a(G1252), .O(gate495inter7));
  inv1  gate1409(.a(G1253), .O(gate495inter8));
  nand2 gate1410(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate1411(.a(s_123), .b(gate495inter3), .O(gate495inter10));
  nor2  gate1412(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate1413(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate1414(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate1597(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate1598(.a(gate497inter0), .b(s_150), .O(gate497inter1));
  and2  gate1599(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate1600(.a(s_150), .O(gate497inter3));
  inv1  gate1601(.a(s_151), .O(gate497inter4));
  nand2 gate1602(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate1603(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate1604(.a(G1256), .O(gate497inter7));
  inv1  gate1605(.a(G1257), .O(gate497inter8));
  nand2 gate1606(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate1607(.a(s_151), .b(gate497inter3), .O(gate497inter10));
  nor2  gate1608(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate1609(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate1610(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate2017(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate2018(.a(gate501inter0), .b(s_210), .O(gate501inter1));
  and2  gate2019(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate2020(.a(s_210), .O(gate501inter3));
  inv1  gate2021(.a(s_211), .O(gate501inter4));
  nand2 gate2022(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate2023(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate2024(.a(G1264), .O(gate501inter7));
  inv1  gate2025(.a(G1265), .O(gate501inter8));
  nand2 gate2026(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate2027(.a(s_211), .b(gate501inter3), .O(gate501inter10));
  nor2  gate2028(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate2029(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate2030(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate1541(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate1542(.a(gate504inter0), .b(s_142), .O(gate504inter1));
  and2  gate1543(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate1544(.a(s_142), .O(gate504inter3));
  inv1  gate1545(.a(s_143), .O(gate504inter4));
  nand2 gate1546(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate1547(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate1548(.a(G1270), .O(gate504inter7));
  inv1  gate1549(.a(G1271), .O(gate504inter8));
  nand2 gate1550(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate1551(.a(s_143), .b(gate504inter3), .O(gate504inter10));
  nor2  gate1552(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate1553(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate1554(.a(gate504inter12), .b(gate504inter1), .O(G1313));

  xor2  gate617(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate618(.a(gate505inter0), .b(s_10), .O(gate505inter1));
  and2  gate619(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate620(.a(s_10), .O(gate505inter3));
  inv1  gate621(.a(s_11), .O(gate505inter4));
  nand2 gate622(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate623(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate624(.a(G1272), .O(gate505inter7));
  inv1  gate625(.a(G1273), .O(gate505inter8));
  nand2 gate626(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate627(.a(s_11), .b(gate505inter3), .O(gate505inter10));
  nor2  gate628(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate629(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate630(.a(gate505inter12), .b(gate505inter1), .O(G1314));
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate855(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate856(.a(gate508inter0), .b(s_44), .O(gate508inter1));
  and2  gate857(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate858(.a(s_44), .O(gate508inter3));
  inv1  gate859(.a(s_45), .O(gate508inter4));
  nand2 gate860(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate861(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate862(.a(G1278), .O(gate508inter7));
  inv1  gate863(.a(G1279), .O(gate508inter8));
  nand2 gate864(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate865(.a(s_45), .b(gate508inter3), .O(gate508inter10));
  nor2  gate866(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate867(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate868(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule