module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );

  xor2  gate561(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate562(.a(gate14inter0), .b(s_2), .O(gate14inter1));
  and2  gate563(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate564(.a(s_2), .O(gate14inter3));
  inv1  gate565(.a(s_3), .O(gate14inter4));
  nand2 gate566(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate567(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate568(.a(G11), .O(gate14inter7));
  inv1  gate569(.a(G12), .O(gate14inter8));
  nand2 gate570(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate571(.a(s_3), .b(gate14inter3), .O(gate14inter10));
  nor2  gate572(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate573(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate574(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate1443(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate1444(.a(gate22inter0), .b(s_128), .O(gate22inter1));
  and2  gate1445(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate1446(.a(s_128), .O(gate22inter3));
  inv1  gate1447(.a(s_129), .O(gate22inter4));
  nand2 gate1448(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate1449(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate1450(.a(G27), .O(gate22inter7));
  inv1  gate1451(.a(G28), .O(gate22inter8));
  nand2 gate1452(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate1453(.a(s_129), .b(gate22inter3), .O(gate22inter10));
  nor2  gate1454(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate1455(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate1456(.a(gate22inter12), .b(gate22inter1), .O(G305));
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate687(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate688(.a(gate24inter0), .b(s_20), .O(gate24inter1));
  and2  gate689(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate690(.a(s_20), .O(gate24inter3));
  inv1  gate691(.a(s_21), .O(gate24inter4));
  nand2 gate692(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate693(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate694(.a(G31), .O(gate24inter7));
  inv1  gate695(.a(G32), .O(gate24inter8));
  nand2 gate696(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate697(.a(s_21), .b(gate24inter3), .O(gate24inter10));
  nor2  gate698(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate699(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate700(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate1065(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate1066(.a(gate28inter0), .b(s_74), .O(gate28inter1));
  and2  gate1067(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate1068(.a(s_74), .O(gate28inter3));
  inv1  gate1069(.a(s_75), .O(gate28inter4));
  nand2 gate1070(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate1071(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate1072(.a(G10), .O(gate28inter7));
  inv1  gate1073(.a(G14), .O(gate28inter8));
  nand2 gate1074(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate1075(.a(s_75), .b(gate28inter3), .O(gate28inter10));
  nor2  gate1076(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate1077(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate1078(.a(gate28inter12), .b(gate28inter1), .O(G323));

  xor2  gate1387(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate1388(.a(gate29inter0), .b(s_120), .O(gate29inter1));
  and2  gate1389(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate1390(.a(s_120), .O(gate29inter3));
  inv1  gate1391(.a(s_121), .O(gate29inter4));
  nand2 gate1392(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate1393(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate1394(.a(G3), .O(gate29inter7));
  inv1  gate1395(.a(G7), .O(gate29inter8));
  nand2 gate1396(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate1397(.a(s_121), .b(gate29inter3), .O(gate29inter10));
  nor2  gate1398(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate1399(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate1400(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );

  xor2  gate1051(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate1052(.a(gate32inter0), .b(s_72), .O(gate32inter1));
  and2  gate1053(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate1054(.a(s_72), .O(gate32inter3));
  inv1  gate1055(.a(s_73), .O(gate32inter4));
  nand2 gate1056(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate1057(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate1058(.a(G12), .O(gate32inter7));
  inv1  gate1059(.a(G16), .O(gate32inter8));
  nand2 gate1060(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate1061(.a(s_73), .b(gate32inter3), .O(gate32inter10));
  nor2  gate1062(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate1063(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate1064(.a(gate32inter12), .b(gate32inter1), .O(G335));
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate1247(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate1248(.a(gate34inter0), .b(s_100), .O(gate34inter1));
  and2  gate1249(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate1250(.a(s_100), .O(gate34inter3));
  inv1  gate1251(.a(s_101), .O(gate34inter4));
  nand2 gate1252(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate1253(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate1254(.a(G25), .O(gate34inter7));
  inv1  gate1255(.a(G29), .O(gate34inter8));
  nand2 gate1256(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate1257(.a(s_101), .b(gate34inter3), .O(gate34inter10));
  nor2  gate1258(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate1259(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate1260(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );

  xor2  gate771(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate772(.a(gate40inter0), .b(s_32), .O(gate40inter1));
  and2  gate773(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate774(.a(s_32), .O(gate40inter3));
  inv1  gate775(.a(s_33), .O(gate40inter4));
  nand2 gate776(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate777(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate778(.a(G28), .O(gate40inter7));
  inv1  gate779(.a(G32), .O(gate40inter8));
  nand2 gate780(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate781(.a(s_33), .b(gate40inter3), .O(gate40inter10));
  nor2  gate782(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate783(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate784(.a(gate40inter12), .b(gate40inter1), .O(G359));
nand2 gate41( .a(G1), .b(G266), .O(G362) );

  xor2  gate673(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate674(.a(gate42inter0), .b(s_18), .O(gate42inter1));
  and2  gate675(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate676(.a(s_18), .O(gate42inter3));
  inv1  gate677(.a(s_19), .O(gate42inter4));
  nand2 gate678(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate679(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate680(.a(G2), .O(gate42inter7));
  inv1  gate681(.a(G266), .O(gate42inter8));
  nand2 gate682(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate683(.a(s_19), .b(gate42inter3), .O(gate42inter10));
  nor2  gate684(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate685(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate686(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );

  xor2  gate617(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate618(.a(gate48inter0), .b(s_10), .O(gate48inter1));
  and2  gate619(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate620(.a(s_10), .O(gate48inter3));
  inv1  gate621(.a(s_11), .O(gate48inter4));
  nand2 gate622(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate623(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate624(.a(G8), .O(gate48inter7));
  inv1  gate625(.a(G275), .O(gate48inter8));
  nand2 gate626(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate627(.a(s_11), .b(gate48inter3), .O(gate48inter10));
  nor2  gate628(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate629(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate630(.a(gate48inter12), .b(gate48inter1), .O(G369));
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate995(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate996(.a(gate52inter0), .b(s_64), .O(gate52inter1));
  and2  gate997(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate998(.a(s_64), .O(gate52inter3));
  inv1  gate999(.a(s_65), .O(gate52inter4));
  nand2 gate1000(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate1001(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate1002(.a(G12), .O(gate52inter7));
  inv1  gate1003(.a(G281), .O(gate52inter8));
  nand2 gate1004(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate1005(.a(s_65), .b(gate52inter3), .O(gate52inter10));
  nor2  gate1006(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate1007(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate1008(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );

  xor2  gate967(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate968(.a(gate68inter0), .b(s_60), .O(gate68inter1));
  and2  gate969(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate970(.a(s_60), .O(gate68inter3));
  inv1  gate971(.a(s_61), .O(gate68inter4));
  nand2 gate972(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate973(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate974(.a(G28), .O(gate68inter7));
  inv1  gate975(.a(G305), .O(gate68inter8));
  nand2 gate976(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate977(.a(s_61), .b(gate68inter3), .O(gate68inter10));
  nor2  gate978(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate979(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate980(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate1359(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate1360(.a(gate77inter0), .b(s_116), .O(gate77inter1));
  and2  gate1361(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate1362(.a(s_116), .O(gate77inter3));
  inv1  gate1363(.a(s_117), .O(gate77inter4));
  nand2 gate1364(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate1365(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate1366(.a(G2), .O(gate77inter7));
  inv1  gate1367(.a(G320), .O(gate77inter8));
  nand2 gate1368(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate1369(.a(s_117), .b(gate77inter3), .O(gate77inter10));
  nor2  gate1370(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate1371(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate1372(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );

  xor2  gate1331(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate1332(.a(gate83inter0), .b(s_112), .O(gate83inter1));
  and2  gate1333(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate1334(.a(s_112), .O(gate83inter3));
  inv1  gate1335(.a(s_113), .O(gate83inter4));
  nand2 gate1336(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate1337(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate1338(.a(G11), .O(gate83inter7));
  inv1  gate1339(.a(G329), .O(gate83inter8));
  nand2 gate1340(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate1341(.a(s_113), .b(gate83inter3), .O(gate83inter10));
  nor2  gate1342(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate1343(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate1344(.a(gate83inter12), .b(gate83inter1), .O(G404));

  xor2  gate547(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate548(.a(gate84inter0), .b(s_0), .O(gate84inter1));
  and2  gate549(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate550(.a(s_0), .O(gate84inter3));
  inv1  gate551(.a(s_1), .O(gate84inter4));
  nand2 gate552(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate553(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate554(.a(G15), .O(gate84inter7));
  inv1  gate555(.a(G329), .O(gate84inter8));
  nand2 gate556(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate557(.a(s_1), .b(gate84inter3), .O(gate84inter10));
  nor2  gate558(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate559(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate560(.a(gate84inter12), .b(gate84inter1), .O(G405));
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );

  xor2  gate785(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate786(.a(gate87inter0), .b(s_34), .O(gate87inter1));
  and2  gate787(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate788(.a(s_34), .O(gate87inter3));
  inv1  gate789(.a(s_35), .O(gate87inter4));
  nand2 gate790(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate791(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate792(.a(G12), .O(gate87inter7));
  inv1  gate793(.a(G335), .O(gate87inter8));
  nand2 gate794(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate795(.a(s_35), .b(gate87inter3), .O(gate87inter10));
  nor2  gate796(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate797(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate798(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate1275(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate1276(.a(gate102inter0), .b(s_104), .O(gate102inter1));
  and2  gate1277(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate1278(.a(s_104), .O(gate102inter3));
  inv1  gate1279(.a(s_105), .O(gate102inter4));
  nand2 gate1280(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate1281(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate1282(.a(G24), .O(gate102inter7));
  inv1  gate1283(.a(G356), .O(gate102inter8));
  nand2 gate1284(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate1285(.a(s_105), .b(gate102inter3), .O(gate102inter10));
  nor2  gate1286(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate1287(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate1288(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate981(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate982(.a(gate108inter0), .b(s_62), .O(gate108inter1));
  and2  gate983(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate984(.a(s_62), .O(gate108inter3));
  inv1  gate985(.a(s_63), .O(gate108inter4));
  nand2 gate986(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate987(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate988(.a(G368), .O(gate108inter7));
  inv1  gate989(.a(G369), .O(gate108inter8));
  nand2 gate990(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate991(.a(s_63), .b(gate108inter3), .O(gate108inter10));
  nor2  gate992(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate993(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate994(.a(gate108inter12), .b(gate108inter1), .O(G435));

  xor2  gate1415(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate1416(.a(gate109inter0), .b(s_124), .O(gate109inter1));
  and2  gate1417(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate1418(.a(s_124), .O(gate109inter3));
  inv1  gate1419(.a(s_125), .O(gate109inter4));
  nand2 gate1420(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate1421(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate1422(.a(G370), .O(gate109inter7));
  inv1  gate1423(.a(G371), .O(gate109inter8));
  nand2 gate1424(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate1425(.a(s_125), .b(gate109inter3), .O(gate109inter10));
  nor2  gate1426(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate1427(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate1428(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );

  xor2  gate1177(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate1178(.a(gate122inter0), .b(s_90), .O(gate122inter1));
  and2  gate1179(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate1180(.a(s_90), .O(gate122inter3));
  inv1  gate1181(.a(s_91), .O(gate122inter4));
  nand2 gate1182(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate1183(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate1184(.a(G396), .O(gate122inter7));
  inv1  gate1185(.a(G397), .O(gate122inter8));
  nand2 gate1186(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate1187(.a(s_91), .b(gate122inter3), .O(gate122inter10));
  nor2  gate1188(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate1189(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate1190(.a(gate122inter12), .b(gate122inter1), .O(G477));
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate1527(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate1528(.a(gate124inter0), .b(s_140), .O(gate124inter1));
  and2  gate1529(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate1530(.a(s_140), .O(gate124inter3));
  inv1  gate1531(.a(s_141), .O(gate124inter4));
  nand2 gate1532(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate1533(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate1534(.a(G400), .O(gate124inter7));
  inv1  gate1535(.a(G401), .O(gate124inter8));
  nand2 gate1536(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate1537(.a(s_141), .b(gate124inter3), .O(gate124inter10));
  nor2  gate1538(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate1539(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate1540(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate603(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate604(.a(gate130inter0), .b(s_8), .O(gate130inter1));
  and2  gate605(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate606(.a(s_8), .O(gate130inter3));
  inv1  gate607(.a(s_9), .O(gate130inter4));
  nand2 gate608(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate609(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate610(.a(G412), .O(gate130inter7));
  inv1  gate611(.a(G413), .O(gate130inter8));
  nand2 gate612(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate613(.a(s_9), .b(gate130inter3), .O(gate130inter10));
  nor2  gate614(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate615(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate616(.a(gate130inter12), .b(gate130inter1), .O(G501));

  xor2  gate813(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate814(.a(gate131inter0), .b(s_38), .O(gate131inter1));
  and2  gate815(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate816(.a(s_38), .O(gate131inter3));
  inv1  gate817(.a(s_39), .O(gate131inter4));
  nand2 gate818(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate819(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate820(.a(G414), .O(gate131inter7));
  inv1  gate821(.a(G415), .O(gate131inter8));
  nand2 gate822(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate823(.a(s_39), .b(gate131inter3), .O(gate131inter10));
  nor2  gate824(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate825(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate826(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );

  xor2  gate1429(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate1430(.a(gate133inter0), .b(s_126), .O(gate133inter1));
  and2  gate1431(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate1432(.a(s_126), .O(gate133inter3));
  inv1  gate1433(.a(s_127), .O(gate133inter4));
  nand2 gate1434(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate1435(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate1436(.a(G418), .O(gate133inter7));
  inv1  gate1437(.a(G419), .O(gate133inter8));
  nand2 gate1438(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate1439(.a(s_127), .b(gate133inter3), .O(gate133inter10));
  nor2  gate1440(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate1441(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate1442(.a(gate133inter12), .b(gate133inter1), .O(G510));
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate1205(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate1206(.a(gate154inter0), .b(s_94), .O(gate154inter1));
  and2  gate1207(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate1208(.a(s_94), .O(gate154inter3));
  inv1  gate1209(.a(s_95), .O(gate154inter4));
  nand2 gate1210(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate1211(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate1212(.a(G429), .O(gate154inter7));
  inv1  gate1213(.a(G522), .O(gate154inter8));
  nand2 gate1214(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate1215(.a(s_95), .b(gate154inter3), .O(gate154inter10));
  nor2  gate1216(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate1217(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate1218(.a(gate154inter12), .b(gate154inter1), .O(G571));

  xor2  gate1611(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate1612(.a(gate155inter0), .b(s_152), .O(gate155inter1));
  and2  gate1613(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate1614(.a(s_152), .O(gate155inter3));
  inv1  gate1615(.a(s_153), .O(gate155inter4));
  nand2 gate1616(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1617(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1618(.a(G432), .O(gate155inter7));
  inv1  gate1619(.a(G525), .O(gate155inter8));
  nand2 gate1620(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1621(.a(s_153), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1622(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1623(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1624(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate743(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate744(.a(gate157inter0), .b(s_28), .O(gate157inter1));
  and2  gate745(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate746(.a(s_28), .O(gate157inter3));
  inv1  gate747(.a(s_29), .O(gate157inter4));
  nand2 gate748(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate749(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate750(.a(G438), .O(gate157inter7));
  inv1  gate751(.a(G528), .O(gate157inter8));
  nand2 gate752(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate753(.a(s_29), .b(gate157inter3), .O(gate157inter10));
  nor2  gate754(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate755(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate756(.a(gate157inter12), .b(gate157inter1), .O(G574));

  xor2  gate1107(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate1108(.a(gate158inter0), .b(s_80), .O(gate158inter1));
  and2  gate1109(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate1110(.a(s_80), .O(gate158inter3));
  inv1  gate1111(.a(s_81), .O(gate158inter4));
  nand2 gate1112(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate1113(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate1114(.a(G441), .O(gate158inter7));
  inv1  gate1115(.a(G528), .O(gate158inter8));
  nand2 gate1116(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate1117(.a(s_81), .b(gate158inter3), .O(gate158inter10));
  nor2  gate1118(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate1119(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate1120(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate1597(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate1598(.a(gate160inter0), .b(s_150), .O(gate160inter1));
  and2  gate1599(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate1600(.a(s_150), .O(gate160inter3));
  inv1  gate1601(.a(s_151), .O(gate160inter4));
  nand2 gate1602(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate1603(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate1604(.a(G447), .O(gate160inter7));
  inv1  gate1605(.a(G531), .O(gate160inter8));
  nand2 gate1606(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate1607(.a(s_151), .b(gate160inter3), .O(gate160inter10));
  nor2  gate1608(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate1609(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate1610(.a(gate160inter12), .b(gate160inter1), .O(G577));

  xor2  gate1639(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate1640(.a(gate161inter0), .b(s_156), .O(gate161inter1));
  and2  gate1641(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate1642(.a(s_156), .O(gate161inter3));
  inv1  gate1643(.a(s_157), .O(gate161inter4));
  nand2 gate1644(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate1645(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate1646(.a(G450), .O(gate161inter7));
  inv1  gate1647(.a(G534), .O(gate161inter8));
  nand2 gate1648(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate1649(.a(s_157), .b(gate161inter3), .O(gate161inter10));
  nor2  gate1650(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate1651(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate1652(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );

  xor2  gate1541(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate1542(.a(gate168inter0), .b(s_142), .O(gate168inter1));
  and2  gate1543(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate1544(.a(s_142), .O(gate168inter3));
  inv1  gate1545(.a(s_143), .O(gate168inter4));
  nand2 gate1546(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate1547(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate1548(.a(G471), .O(gate168inter7));
  inv1  gate1549(.a(G543), .O(gate168inter8));
  nand2 gate1550(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate1551(.a(s_143), .b(gate168inter3), .O(gate168inter10));
  nor2  gate1552(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate1553(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate1554(.a(gate168inter12), .b(gate168inter1), .O(G585));
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );

  xor2  gate1457(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate1458(.a(gate202inter0), .b(s_130), .O(gate202inter1));
  and2  gate1459(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate1460(.a(s_130), .O(gate202inter3));
  inv1  gate1461(.a(s_131), .O(gate202inter4));
  nand2 gate1462(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate1463(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate1464(.a(G612), .O(gate202inter7));
  inv1  gate1465(.a(G617), .O(gate202inter8));
  nand2 gate1466(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate1467(.a(s_131), .b(gate202inter3), .O(gate202inter10));
  nor2  gate1468(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate1469(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate1470(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate1345(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate1346(.a(gate205inter0), .b(s_114), .O(gate205inter1));
  and2  gate1347(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate1348(.a(s_114), .O(gate205inter3));
  inv1  gate1349(.a(s_115), .O(gate205inter4));
  nand2 gate1350(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate1351(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate1352(.a(G622), .O(gate205inter7));
  inv1  gate1353(.a(G627), .O(gate205inter8));
  nand2 gate1354(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate1355(.a(s_115), .b(gate205inter3), .O(gate205inter10));
  nor2  gate1356(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate1357(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate1358(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );

  xor2  gate939(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate940(.a(gate210inter0), .b(s_56), .O(gate210inter1));
  and2  gate941(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate942(.a(s_56), .O(gate210inter3));
  inv1  gate943(.a(s_57), .O(gate210inter4));
  nand2 gate944(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate945(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate946(.a(G607), .O(gate210inter7));
  inv1  gate947(.a(G666), .O(gate210inter8));
  nand2 gate948(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate949(.a(s_57), .b(gate210inter3), .O(gate210inter10));
  nor2  gate950(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate951(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate952(.a(gate210inter12), .b(gate210inter1), .O(G691));
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate1009(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate1010(.a(gate215inter0), .b(s_66), .O(gate215inter1));
  and2  gate1011(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate1012(.a(s_66), .O(gate215inter3));
  inv1  gate1013(.a(s_67), .O(gate215inter4));
  nand2 gate1014(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate1015(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate1016(.a(G607), .O(gate215inter7));
  inv1  gate1017(.a(G675), .O(gate215inter8));
  nand2 gate1018(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate1019(.a(s_67), .b(gate215inter3), .O(gate215inter10));
  nor2  gate1020(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate1021(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate1022(.a(gate215inter12), .b(gate215inter1), .O(G696));

  xor2  gate631(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate632(.a(gate216inter0), .b(s_12), .O(gate216inter1));
  and2  gate633(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate634(.a(s_12), .O(gate216inter3));
  inv1  gate635(.a(s_13), .O(gate216inter4));
  nand2 gate636(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate637(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate638(.a(G617), .O(gate216inter7));
  inv1  gate639(.a(G675), .O(gate216inter8));
  nand2 gate640(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate641(.a(s_13), .b(gate216inter3), .O(gate216inter10));
  nor2  gate642(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate643(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate644(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate645(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate646(.a(gate224inter0), .b(s_14), .O(gate224inter1));
  and2  gate647(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate648(.a(s_14), .O(gate224inter3));
  inv1  gate649(.a(s_15), .O(gate224inter4));
  nand2 gate650(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate651(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate652(.a(G637), .O(gate224inter7));
  inv1  gate653(.a(G687), .O(gate224inter8));
  nand2 gate654(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate655(.a(s_15), .b(gate224inter3), .O(gate224inter10));
  nor2  gate656(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate657(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate658(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate1513(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate1514(.a(gate227inter0), .b(s_138), .O(gate227inter1));
  and2  gate1515(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate1516(.a(s_138), .O(gate227inter3));
  inv1  gate1517(.a(s_139), .O(gate227inter4));
  nand2 gate1518(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate1519(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate1520(.a(G694), .O(gate227inter7));
  inv1  gate1521(.a(G695), .O(gate227inter8));
  nand2 gate1522(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate1523(.a(s_139), .b(gate227inter3), .O(gate227inter10));
  nor2  gate1524(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate1525(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate1526(.a(gate227inter12), .b(gate227inter1), .O(G712));
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );

  xor2  gate1499(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate1500(.a(gate230inter0), .b(s_136), .O(gate230inter1));
  and2  gate1501(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate1502(.a(s_136), .O(gate230inter3));
  inv1  gate1503(.a(s_137), .O(gate230inter4));
  nand2 gate1504(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate1505(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate1506(.a(G700), .O(gate230inter7));
  inv1  gate1507(.a(G701), .O(gate230inter8));
  nand2 gate1508(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate1509(.a(s_137), .b(gate230inter3), .O(gate230inter10));
  nor2  gate1510(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate1511(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate1512(.a(gate230inter12), .b(gate230inter1), .O(G721));
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );

  xor2  gate1149(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate1150(.a(gate235inter0), .b(s_86), .O(gate235inter1));
  and2  gate1151(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate1152(.a(s_86), .O(gate235inter3));
  inv1  gate1153(.a(s_87), .O(gate235inter4));
  nand2 gate1154(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate1155(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate1156(.a(G248), .O(gate235inter7));
  inv1  gate1157(.a(G724), .O(gate235inter8));
  nand2 gate1158(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate1159(.a(s_87), .b(gate235inter3), .O(gate235inter10));
  nor2  gate1160(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate1161(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate1162(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );

  xor2  gate701(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate702(.a(gate239inter0), .b(s_22), .O(gate239inter1));
  and2  gate703(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate704(.a(s_22), .O(gate239inter3));
  inv1  gate705(.a(s_23), .O(gate239inter4));
  nand2 gate706(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate707(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate708(.a(G260), .O(gate239inter7));
  inv1  gate709(.a(G712), .O(gate239inter8));
  nand2 gate710(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate711(.a(s_23), .b(gate239inter3), .O(gate239inter10));
  nor2  gate712(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate713(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate714(.a(gate239inter12), .b(gate239inter1), .O(G748));
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );

  xor2  gate953(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate954(.a(gate242inter0), .b(s_58), .O(gate242inter1));
  and2  gate955(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate956(.a(s_58), .O(gate242inter3));
  inv1  gate957(.a(s_59), .O(gate242inter4));
  nand2 gate958(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate959(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate960(.a(G718), .O(gate242inter7));
  inv1  gate961(.a(G730), .O(gate242inter8));
  nand2 gate962(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate963(.a(s_59), .b(gate242inter3), .O(gate242inter10));
  nor2  gate964(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate965(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate966(.a(gate242inter12), .b(gate242inter1), .O(G755));
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate575(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate576(.a(gate248inter0), .b(s_4), .O(gate248inter1));
  and2  gate577(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate578(.a(s_4), .O(gate248inter3));
  inv1  gate579(.a(s_5), .O(gate248inter4));
  nand2 gate580(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate581(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate582(.a(G727), .O(gate248inter7));
  inv1  gate583(.a(G739), .O(gate248inter8));
  nand2 gate584(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate585(.a(s_5), .b(gate248inter3), .O(gate248inter10));
  nor2  gate586(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate587(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate588(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate1485(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate1486(.a(gate252inter0), .b(s_134), .O(gate252inter1));
  and2  gate1487(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate1488(.a(s_134), .O(gate252inter3));
  inv1  gate1489(.a(s_135), .O(gate252inter4));
  nand2 gate1490(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate1491(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate1492(.a(G709), .O(gate252inter7));
  inv1  gate1493(.a(G745), .O(gate252inter8));
  nand2 gate1494(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate1495(.a(s_135), .b(gate252inter3), .O(gate252inter10));
  nor2  gate1496(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate1497(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate1498(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );

  xor2  gate1079(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate1080(.a(gate259inter0), .b(s_76), .O(gate259inter1));
  and2  gate1081(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate1082(.a(s_76), .O(gate259inter3));
  inv1  gate1083(.a(s_77), .O(gate259inter4));
  nand2 gate1084(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate1085(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate1086(.a(G758), .O(gate259inter7));
  inv1  gate1087(.a(G759), .O(gate259inter8));
  nand2 gate1088(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate1089(.a(s_77), .b(gate259inter3), .O(gate259inter10));
  nor2  gate1090(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate1091(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate1092(.a(gate259inter12), .b(gate259inter1), .O(G776));
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate827(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate828(.a(gate261inter0), .b(s_40), .O(gate261inter1));
  and2  gate829(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate830(.a(s_40), .O(gate261inter3));
  inv1  gate831(.a(s_41), .O(gate261inter4));
  nand2 gate832(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate833(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate834(.a(G762), .O(gate261inter7));
  inv1  gate835(.a(G763), .O(gate261inter8));
  nand2 gate836(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate837(.a(s_41), .b(gate261inter3), .O(gate261inter10));
  nor2  gate838(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate839(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate840(.a(gate261inter12), .b(gate261inter1), .O(G782));

  xor2  gate1135(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate1136(.a(gate262inter0), .b(s_84), .O(gate262inter1));
  and2  gate1137(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate1138(.a(s_84), .O(gate262inter3));
  inv1  gate1139(.a(s_85), .O(gate262inter4));
  nand2 gate1140(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate1141(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate1142(.a(G764), .O(gate262inter7));
  inv1  gate1143(.a(G765), .O(gate262inter8));
  nand2 gate1144(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate1145(.a(s_85), .b(gate262inter3), .O(gate262inter10));
  nor2  gate1146(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate1147(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate1148(.a(gate262inter12), .b(gate262inter1), .O(G785));

  xor2  gate1219(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate1220(.a(gate263inter0), .b(s_96), .O(gate263inter1));
  and2  gate1221(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate1222(.a(s_96), .O(gate263inter3));
  inv1  gate1223(.a(s_97), .O(gate263inter4));
  nand2 gate1224(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate1225(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate1226(.a(G766), .O(gate263inter7));
  inv1  gate1227(.a(G767), .O(gate263inter8));
  nand2 gate1228(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate1229(.a(s_97), .b(gate263inter3), .O(gate263inter10));
  nor2  gate1230(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate1231(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate1232(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate897(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate898(.a(gate265inter0), .b(s_50), .O(gate265inter1));
  and2  gate899(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate900(.a(s_50), .O(gate265inter3));
  inv1  gate901(.a(s_51), .O(gate265inter4));
  nand2 gate902(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate903(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate904(.a(G642), .O(gate265inter7));
  inv1  gate905(.a(G770), .O(gate265inter8));
  nand2 gate906(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate907(.a(s_51), .b(gate265inter3), .O(gate265inter10));
  nor2  gate908(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate909(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate910(.a(gate265inter12), .b(gate265inter1), .O(G794));

  xor2  gate729(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate730(.a(gate266inter0), .b(s_26), .O(gate266inter1));
  and2  gate731(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate732(.a(s_26), .O(gate266inter3));
  inv1  gate733(.a(s_27), .O(gate266inter4));
  nand2 gate734(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate735(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate736(.a(G645), .O(gate266inter7));
  inv1  gate737(.a(G773), .O(gate266inter8));
  nand2 gate738(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate739(.a(s_27), .b(gate266inter3), .O(gate266inter10));
  nor2  gate740(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate741(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate742(.a(gate266inter12), .b(gate266inter1), .O(G797));

  xor2  gate1261(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate1262(.a(gate267inter0), .b(s_102), .O(gate267inter1));
  and2  gate1263(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate1264(.a(s_102), .O(gate267inter3));
  inv1  gate1265(.a(s_103), .O(gate267inter4));
  nand2 gate1266(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate1267(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate1268(.a(G648), .O(gate267inter7));
  inv1  gate1269(.a(G776), .O(gate267inter8));
  nand2 gate1270(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate1271(.a(s_103), .b(gate267inter3), .O(gate267inter10));
  nor2  gate1272(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate1273(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate1274(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate1555(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate1556(.a(gate282inter0), .b(s_144), .O(gate282inter1));
  and2  gate1557(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate1558(.a(s_144), .O(gate282inter3));
  inv1  gate1559(.a(s_145), .O(gate282inter4));
  nand2 gate1560(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate1561(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate1562(.a(G782), .O(gate282inter7));
  inv1  gate1563(.a(G806), .O(gate282inter8));
  nand2 gate1564(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate1565(.a(s_145), .b(gate282inter3), .O(gate282inter10));
  nor2  gate1566(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate1567(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate1568(.a(gate282inter12), .b(gate282inter1), .O(G827));

  xor2  gate1625(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate1626(.a(gate283inter0), .b(s_154), .O(gate283inter1));
  and2  gate1627(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate1628(.a(s_154), .O(gate283inter3));
  inv1  gate1629(.a(s_155), .O(gate283inter4));
  nand2 gate1630(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate1631(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate1632(.a(G657), .O(gate283inter7));
  inv1  gate1633(.a(G809), .O(gate283inter8));
  nand2 gate1634(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate1635(.a(s_155), .b(gate283inter3), .O(gate283inter10));
  nor2  gate1636(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate1637(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate1638(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate589(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate590(.a(gate285inter0), .b(s_6), .O(gate285inter1));
  and2  gate591(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate592(.a(s_6), .O(gate285inter3));
  inv1  gate593(.a(s_7), .O(gate285inter4));
  nand2 gate594(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate595(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate596(.a(G660), .O(gate285inter7));
  inv1  gate597(.a(G812), .O(gate285inter8));
  nand2 gate598(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate599(.a(s_7), .b(gate285inter3), .O(gate285inter10));
  nor2  gate600(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate601(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate602(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate1037(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate1038(.a(gate289inter0), .b(s_70), .O(gate289inter1));
  and2  gate1039(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate1040(.a(s_70), .O(gate289inter3));
  inv1  gate1041(.a(s_71), .O(gate289inter4));
  nand2 gate1042(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate1043(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate1044(.a(G818), .O(gate289inter7));
  inv1  gate1045(.a(G819), .O(gate289inter8));
  nand2 gate1046(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate1047(.a(s_71), .b(gate289inter3), .O(gate289inter10));
  nor2  gate1048(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate1049(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate1050(.a(gate289inter12), .b(gate289inter1), .O(G834));

  xor2  gate1583(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate1584(.a(gate290inter0), .b(s_148), .O(gate290inter1));
  and2  gate1585(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate1586(.a(s_148), .O(gate290inter3));
  inv1  gate1587(.a(s_149), .O(gate290inter4));
  nand2 gate1588(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate1589(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate1590(.a(G820), .O(gate290inter7));
  inv1  gate1591(.a(G821), .O(gate290inter8));
  nand2 gate1592(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate1593(.a(s_149), .b(gate290inter3), .O(gate290inter10));
  nor2  gate1594(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate1595(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate1596(.a(gate290inter12), .b(gate290inter1), .O(G847));

  xor2  gate659(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate660(.a(gate291inter0), .b(s_16), .O(gate291inter1));
  and2  gate661(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate662(.a(s_16), .O(gate291inter3));
  inv1  gate663(.a(s_17), .O(gate291inter4));
  nand2 gate664(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate665(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate666(.a(G822), .O(gate291inter7));
  inv1  gate667(.a(G823), .O(gate291inter8));
  nand2 gate668(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate669(.a(s_17), .b(gate291inter3), .O(gate291inter10));
  nor2  gate670(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate671(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate672(.a(gate291inter12), .b(gate291inter1), .O(G860));

  xor2  gate1163(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate1164(.a(gate292inter0), .b(s_88), .O(gate292inter1));
  and2  gate1165(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate1166(.a(s_88), .O(gate292inter3));
  inv1  gate1167(.a(s_89), .O(gate292inter4));
  nand2 gate1168(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate1169(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate1170(.a(G824), .O(gate292inter7));
  inv1  gate1171(.a(G825), .O(gate292inter8));
  nand2 gate1172(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate1173(.a(s_89), .b(gate292inter3), .O(gate292inter10));
  nor2  gate1174(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate1175(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate1176(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate1121(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate1122(.a(gate295inter0), .b(s_82), .O(gate295inter1));
  and2  gate1123(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate1124(.a(s_82), .O(gate295inter3));
  inv1  gate1125(.a(s_83), .O(gate295inter4));
  nand2 gate1126(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate1127(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate1128(.a(G830), .O(gate295inter7));
  inv1  gate1129(.a(G831), .O(gate295inter8));
  nand2 gate1130(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate1131(.a(s_83), .b(gate295inter3), .O(gate295inter10));
  nor2  gate1132(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate1133(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate1134(.a(gate295inter12), .b(gate295inter1), .O(G912));
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate1093(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate1094(.a(gate390inter0), .b(s_78), .O(gate390inter1));
  and2  gate1095(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate1096(.a(s_78), .O(gate390inter3));
  inv1  gate1097(.a(s_79), .O(gate390inter4));
  nand2 gate1098(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate1099(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate1100(.a(G4), .O(gate390inter7));
  inv1  gate1101(.a(G1045), .O(gate390inter8));
  nand2 gate1102(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate1103(.a(s_79), .b(gate390inter3), .O(gate390inter10));
  nor2  gate1104(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate1105(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate1106(.a(gate390inter12), .b(gate390inter1), .O(G1141));

  xor2  gate1191(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate1192(.a(gate391inter0), .b(s_92), .O(gate391inter1));
  and2  gate1193(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate1194(.a(s_92), .O(gate391inter3));
  inv1  gate1195(.a(s_93), .O(gate391inter4));
  nand2 gate1196(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate1197(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate1198(.a(G5), .O(gate391inter7));
  inv1  gate1199(.a(G1048), .O(gate391inter8));
  nand2 gate1200(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate1201(.a(s_93), .b(gate391inter3), .O(gate391inter10));
  nor2  gate1202(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate1203(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate1204(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate869(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate870(.a(gate398inter0), .b(s_46), .O(gate398inter1));
  and2  gate871(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate872(.a(s_46), .O(gate398inter3));
  inv1  gate873(.a(s_47), .O(gate398inter4));
  nand2 gate874(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate875(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate876(.a(G12), .O(gate398inter7));
  inv1  gate877(.a(G1069), .O(gate398inter8));
  nand2 gate878(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate879(.a(s_47), .b(gate398inter3), .O(gate398inter10));
  nor2  gate880(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate881(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate882(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate715(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate716(.a(gate411inter0), .b(s_24), .O(gate411inter1));
  and2  gate717(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate718(.a(s_24), .O(gate411inter3));
  inv1  gate719(.a(s_25), .O(gate411inter4));
  nand2 gate720(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate721(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate722(.a(G25), .O(gate411inter7));
  inv1  gate723(.a(G1108), .O(gate411inter8));
  nand2 gate724(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate725(.a(s_25), .b(gate411inter3), .O(gate411inter10));
  nor2  gate726(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate727(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate728(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate1233(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate1234(.a(gate421inter0), .b(s_98), .O(gate421inter1));
  and2  gate1235(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate1236(.a(s_98), .O(gate421inter3));
  inv1  gate1237(.a(s_99), .O(gate421inter4));
  nand2 gate1238(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate1239(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate1240(.a(G2), .O(gate421inter7));
  inv1  gate1241(.a(G1135), .O(gate421inter8));
  nand2 gate1242(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate1243(.a(s_99), .b(gate421inter3), .O(gate421inter10));
  nor2  gate1244(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate1245(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate1246(.a(gate421inter12), .b(gate421inter1), .O(G1230));
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );

  xor2  gate1569(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate1570(.a(gate426inter0), .b(s_146), .O(gate426inter1));
  and2  gate1571(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate1572(.a(s_146), .O(gate426inter3));
  inv1  gate1573(.a(s_147), .O(gate426inter4));
  nand2 gate1574(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate1575(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate1576(.a(G1045), .O(gate426inter7));
  inv1  gate1577(.a(G1141), .O(gate426inter8));
  nand2 gate1578(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate1579(.a(s_147), .b(gate426inter3), .O(gate426inter10));
  nor2  gate1580(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate1581(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate1582(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate1471(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate1472(.a(gate428inter0), .b(s_132), .O(gate428inter1));
  and2  gate1473(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate1474(.a(s_132), .O(gate428inter3));
  inv1  gate1475(.a(s_133), .O(gate428inter4));
  nand2 gate1476(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate1477(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate1478(.a(G1048), .O(gate428inter7));
  inv1  gate1479(.a(G1144), .O(gate428inter8));
  nand2 gate1480(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate1481(.a(s_133), .b(gate428inter3), .O(gate428inter10));
  nor2  gate1482(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate1483(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate1484(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );

  xor2  gate757(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate758(.a(gate449inter0), .b(s_30), .O(gate449inter1));
  and2  gate759(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate760(.a(s_30), .O(gate449inter3));
  inv1  gate761(.a(s_31), .O(gate449inter4));
  nand2 gate762(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate763(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate764(.a(G16), .O(gate449inter7));
  inv1  gate765(.a(G1177), .O(gate449inter8));
  nand2 gate766(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate767(.a(s_31), .b(gate449inter3), .O(gate449inter10));
  nor2  gate768(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate769(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate770(.a(gate449inter12), .b(gate449inter1), .O(G1258));

  xor2  gate1667(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate1668(.a(gate450inter0), .b(s_160), .O(gate450inter1));
  and2  gate1669(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate1670(.a(s_160), .O(gate450inter3));
  inv1  gate1671(.a(s_161), .O(gate450inter4));
  nand2 gate1672(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate1673(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate1674(.a(G1081), .O(gate450inter7));
  inv1  gate1675(.a(G1177), .O(gate450inter8));
  nand2 gate1676(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate1677(.a(s_161), .b(gate450inter3), .O(gate450inter10));
  nor2  gate1678(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate1679(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate1680(.a(gate450inter12), .b(gate450inter1), .O(G1259));

  xor2  gate841(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate842(.a(gate451inter0), .b(s_42), .O(gate451inter1));
  and2  gate843(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate844(.a(s_42), .O(gate451inter3));
  inv1  gate845(.a(s_43), .O(gate451inter4));
  nand2 gate846(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate847(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate848(.a(G17), .O(gate451inter7));
  inv1  gate849(.a(G1180), .O(gate451inter8));
  nand2 gate850(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate851(.a(s_43), .b(gate451inter3), .O(gate451inter10));
  nor2  gate852(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate853(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate854(.a(gate451inter12), .b(gate451inter1), .O(G1260));
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );

  xor2  gate925(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate926(.a(gate455inter0), .b(s_54), .O(gate455inter1));
  and2  gate927(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate928(.a(s_54), .O(gate455inter3));
  inv1  gate929(.a(s_55), .O(gate455inter4));
  nand2 gate930(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate931(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate932(.a(G19), .O(gate455inter7));
  inv1  gate933(.a(G1186), .O(gate455inter8));
  nand2 gate934(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate935(.a(s_55), .b(gate455inter3), .O(gate455inter10));
  nor2  gate936(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate937(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate938(.a(gate455inter12), .b(gate455inter1), .O(G1264));
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate1653(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate1654(.a(gate463inter0), .b(s_158), .O(gate463inter1));
  and2  gate1655(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate1656(.a(s_158), .O(gate463inter3));
  inv1  gate1657(.a(s_159), .O(gate463inter4));
  nand2 gate1658(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate1659(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate1660(.a(G23), .O(gate463inter7));
  inv1  gate1661(.a(G1198), .O(gate463inter8));
  nand2 gate1662(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate1663(.a(s_159), .b(gate463inter3), .O(gate463inter10));
  nor2  gate1664(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate1665(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate1666(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );

  xor2  gate1317(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate1318(.a(gate470inter0), .b(s_110), .O(gate470inter1));
  and2  gate1319(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate1320(.a(s_110), .O(gate470inter3));
  inv1  gate1321(.a(s_111), .O(gate470inter4));
  nand2 gate1322(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate1323(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate1324(.a(G1111), .O(gate470inter7));
  inv1  gate1325(.a(G1207), .O(gate470inter8));
  nand2 gate1326(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate1327(.a(s_111), .b(gate470inter3), .O(gate470inter10));
  nor2  gate1328(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate1329(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate1330(.a(gate470inter12), .b(gate470inter1), .O(G1279));
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate1373(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate1374(.a(gate472inter0), .b(s_118), .O(gate472inter1));
  and2  gate1375(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate1376(.a(s_118), .O(gate472inter3));
  inv1  gate1377(.a(s_119), .O(gate472inter4));
  nand2 gate1378(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate1379(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate1380(.a(G1114), .O(gate472inter7));
  inv1  gate1381(.a(G1210), .O(gate472inter8));
  nand2 gate1382(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate1383(.a(s_119), .b(gate472inter3), .O(gate472inter10));
  nor2  gate1384(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate1385(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate1386(.a(gate472inter12), .b(gate472inter1), .O(G1281));

  xor2  gate911(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate912(.a(gate473inter0), .b(s_52), .O(gate473inter1));
  and2  gate913(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate914(.a(s_52), .O(gate473inter3));
  inv1  gate915(.a(s_53), .O(gate473inter4));
  nand2 gate916(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate917(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate918(.a(G28), .O(gate473inter7));
  inv1  gate919(.a(G1213), .O(gate473inter8));
  nand2 gate920(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate921(.a(s_53), .b(gate473inter3), .O(gate473inter10));
  nor2  gate922(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate923(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate924(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate1023(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate1024(.a(gate477inter0), .b(s_68), .O(gate477inter1));
  and2  gate1025(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate1026(.a(s_68), .O(gate477inter3));
  inv1  gate1027(.a(s_69), .O(gate477inter4));
  nand2 gate1028(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate1029(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate1030(.a(G30), .O(gate477inter7));
  inv1  gate1031(.a(G1219), .O(gate477inter8));
  nand2 gate1032(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate1033(.a(s_69), .b(gate477inter3), .O(gate477inter10));
  nor2  gate1034(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate1035(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate1036(.a(gate477inter12), .b(gate477inter1), .O(G1286));

  xor2  gate1303(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate1304(.a(gate478inter0), .b(s_108), .O(gate478inter1));
  and2  gate1305(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate1306(.a(s_108), .O(gate478inter3));
  inv1  gate1307(.a(s_109), .O(gate478inter4));
  nand2 gate1308(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate1309(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate1310(.a(G1123), .O(gate478inter7));
  inv1  gate1311(.a(G1219), .O(gate478inter8));
  nand2 gate1312(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate1313(.a(s_109), .b(gate478inter3), .O(gate478inter10));
  nor2  gate1314(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate1315(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate1316(.a(gate478inter12), .b(gate478inter1), .O(G1287));

  xor2  gate1289(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate1290(.a(gate479inter0), .b(s_106), .O(gate479inter1));
  and2  gate1291(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate1292(.a(s_106), .O(gate479inter3));
  inv1  gate1293(.a(s_107), .O(gate479inter4));
  nand2 gate1294(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate1295(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate1296(.a(G31), .O(gate479inter7));
  inv1  gate1297(.a(G1222), .O(gate479inter8));
  nand2 gate1298(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate1299(.a(s_107), .b(gate479inter3), .O(gate479inter10));
  nor2  gate1300(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate1301(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate1302(.a(gate479inter12), .b(gate479inter1), .O(G1288));

  xor2  gate1401(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate1402(.a(gate480inter0), .b(s_122), .O(gate480inter1));
  and2  gate1403(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate1404(.a(s_122), .O(gate480inter3));
  inv1  gate1405(.a(s_123), .O(gate480inter4));
  nand2 gate1406(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate1407(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate1408(.a(G1126), .O(gate480inter7));
  inv1  gate1409(.a(G1222), .O(gate480inter8));
  nand2 gate1410(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate1411(.a(s_123), .b(gate480inter3), .O(gate480inter10));
  nor2  gate1412(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate1413(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate1414(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate883(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate884(.a(gate488inter0), .b(s_48), .O(gate488inter1));
  and2  gate885(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate886(.a(s_48), .O(gate488inter3));
  inv1  gate887(.a(s_49), .O(gate488inter4));
  nand2 gate888(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate889(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate890(.a(G1238), .O(gate488inter7));
  inv1  gate891(.a(G1239), .O(gate488inter8));
  nand2 gate892(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate893(.a(s_49), .b(gate488inter3), .O(gate488inter10));
  nor2  gate894(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate895(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate896(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate855(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate856(.a(gate499inter0), .b(s_44), .O(gate499inter1));
  and2  gate857(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate858(.a(s_44), .O(gate499inter3));
  inv1  gate859(.a(s_45), .O(gate499inter4));
  nand2 gate860(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate861(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate862(.a(G1260), .O(gate499inter7));
  inv1  gate863(.a(G1261), .O(gate499inter8));
  nand2 gate864(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate865(.a(s_45), .b(gate499inter3), .O(gate499inter10));
  nor2  gate866(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate867(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate868(.a(gate499inter12), .b(gate499inter1), .O(G1308));

  xor2  gate799(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate800(.a(gate500inter0), .b(s_36), .O(gate500inter1));
  and2  gate801(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate802(.a(s_36), .O(gate500inter3));
  inv1  gate803(.a(s_37), .O(gate500inter4));
  nand2 gate804(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate805(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate806(.a(G1262), .O(gate500inter7));
  inv1  gate807(.a(G1263), .O(gate500inter8));
  nand2 gate808(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate809(.a(s_37), .b(gate500inter3), .O(gate500inter10));
  nor2  gate810(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate811(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate812(.a(gate500inter12), .b(gate500inter1), .O(G1309));
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule