module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281, s_282, s_283, s_284, s_285, s_286, s_287, s_288, s_289, s_290, s_291;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );

  xor2  gate1611(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate1612(.a(gate10inter0), .b(s_152), .O(gate10inter1));
  and2  gate1613(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate1614(.a(s_152), .O(gate10inter3));
  inv1  gate1615(.a(s_153), .O(gate10inter4));
  nand2 gate1616(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate1617(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate1618(.a(G3), .O(gate10inter7));
  inv1  gate1619(.a(G4), .O(gate10inter8));
  nand2 gate1620(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate1621(.a(s_153), .b(gate10inter3), .O(gate10inter10));
  nor2  gate1622(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate1623(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate1624(.a(gate10inter12), .b(gate10inter1), .O(G269));

  xor2  gate729(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate730(.a(gate11inter0), .b(s_26), .O(gate11inter1));
  and2  gate731(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate732(.a(s_26), .O(gate11inter3));
  inv1  gate733(.a(s_27), .O(gate11inter4));
  nand2 gate734(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate735(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate736(.a(G5), .O(gate11inter7));
  inv1  gate737(.a(G6), .O(gate11inter8));
  nand2 gate738(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate739(.a(s_27), .b(gate11inter3), .O(gate11inter10));
  nor2  gate740(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate741(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate742(.a(gate11inter12), .b(gate11inter1), .O(G272));

  xor2  gate1933(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate1934(.a(gate12inter0), .b(s_198), .O(gate12inter1));
  and2  gate1935(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate1936(.a(s_198), .O(gate12inter3));
  inv1  gate1937(.a(s_199), .O(gate12inter4));
  nand2 gate1938(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate1939(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate1940(.a(G7), .O(gate12inter7));
  inv1  gate1941(.a(G8), .O(gate12inter8));
  nand2 gate1942(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate1943(.a(s_199), .b(gate12inter3), .O(gate12inter10));
  nor2  gate1944(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate1945(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate1946(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );

  xor2  gate2185(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate2186(.a(gate14inter0), .b(s_234), .O(gate14inter1));
  and2  gate2187(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate2188(.a(s_234), .O(gate14inter3));
  inv1  gate2189(.a(s_235), .O(gate14inter4));
  nand2 gate2190(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate2191(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate2192(.a(G11), .O(gate14inter7));
  inv1  gate2193(.a(G12), .O(gate14inter8));
  nand2 gate2194(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate2195(.a(s_235), .b(gate14inter3), .O(gate14inter10));
  nor2  gate2196(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate2197(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate2198(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate1499(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate1500(.a(gate16inter0), .b(s_136), .O(gate16inter1));
  and2  gate1501(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate1502(.a(s_136), .O(gate16inter3));
  inv1  gate1503(.a(s_137), .O(gate16inter4));
  nand2 gate1504(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate1505(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate1506(.a(G15), .O(gate16inter7));
  inv1  gate1507(.a(G16), .O(gate16inter8));
  nand2 gate1508(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate1509(.a(s_137), .b(gate16inter3), .O(gate16inter10));
  nor2  gate1510(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate1511(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate1512(.a(gate16inter12), .b(gate16inter1), .O(G287));

  xor2  gate757(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate758(.a(gate17inter0), .b(s_30), .O(gate17inter1));
  and2  gate759(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate760(.a(s_30), .O(gate17inter3));
  inv1  gate761(.a(s_31), .O(gate17inter4));
  nand2 gate762(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate763(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate764(.a(G17), .O(gate17inter7));
  inv1  gate765(.a(G18), .O(gate17inter8));
  nand2 gate766(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate767(.a(s_31), .b(gate17inter3), .O(gate17inter10));
  nor2  gate768(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate769(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate770(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate1107(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate1108(.a(gate19inter0), .b(s_80), .O(gate19inter1));
  and2  gate1109(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate1110(.a(s_80), .O(gate19inter3));
  inv1  gate1111(.a(s_81), .O(gate19inter4));
  nand2 gate1112(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate1113(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate1114(.a(G21), .O(gate19inter7));
  inv1  gate1115(.a(G22), .O(gate19inter8));
  nand2 gate1116(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate1117(.a(s_81), .b(gate19inter3), .O(gate19inter10));
  nor2  gate1118(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate1119(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate1120(.a(gate19inter12), .b(gate19inter1), .O(G296));

  xor2  gate743(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate744(.a(gate20inter0), .b(s_28), .O(gate20inter1));
  and2  gate745(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate746(.a(s_28), .O(gate20inter3));
  inv1  gate747(.a(s_29), .O(gate20inter4));
  nand2 gate748(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate749(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate750(.a(G23), .O(gate20inter7));
  inv1  gate751(.a(G24), .O(gate20inter8));
  nand2 gate752(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate753(.a(s_29), .b(gate20inter3), .O(gate20inter10));
  nor2  gate754(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate755(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate756(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate2395(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate2396(.a(gate22inter0), .b(s_264), .O(gate22inter1));
  and2  gate2397(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate2398(.a(s_264), .O(gate22inter3));
  inv1  gate2399(.a(s_265), .O(gate22inter4));
  nand2 gate2400(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate2401(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate2402(.a(G27), .O(gate22inter7));
  inv1  gate2403(.a(G28), .O(gate22inter8));
  nand2 gate2404(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate2405(.a(s_265), .b(gate22inter3), .O(gate22inter10));
  nor2  gate2406(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate2407(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate2408(.a(gate22inter12), .b(gate22inter1), .O(G305));
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate2493(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate2494(.a(gate25inter0), .b(s_278), .O(gate25inter1));
  and2  gate2495(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate2496(.a(s_278), .O(gate25inter3));
  inv1  gate2497(.a(s_279), .O(gate25inter4));
  nand2 gate2498(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate2499(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate2500(.a(G1), .O(gate25inter7));
  inv1  gate2501(.a(G5), .O(gate25inter8));
  nand2 gate2502(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate2503(.a(s_279), .b(gate25inter3), .O(gate25inter10));
  nor2  gate2504(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate2505(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate2506(.a(gate25inter12), .b(gate25inter1), .O(G314));

  xor2  gate967(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate968(.a(gate26inter0), .b(s_60), .O(gate26inter1));
  and2  gate969(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate970(.a(s_60), .O(gate26inter3));
  inv1  gate971(.a(s_61), .O(gate26inter4));
  nand2 gate972(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate973(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate974(.a(G9), .O(gate26inter7));
  inv1  gate975(.a(G13), .O(gate26inter8));
  nand2 gate976(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate977(.a(s_61), .b(gate26inter3), .O(gate26inter10));
  nor2  gate978(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate979(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate980(.a(gate26inter12), .b(gate26inter1), .O(G317));

  xor2  gate1079(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate1080(.a(gate27inter0), .b(s_76), .O(gate27inter1));
  and2  gate1081(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate1082(.a(s_76), .O(gate27inter3));
  inv1  gate1083(.a(s_77), .O(gate27inter4));
  nand2 gate1084(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate1085(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate1086(.a(G2), .O(gate27inter7));
  inv1  gate1087(.a(G6), .O(gate27inter8));
  nand2 gate1088(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate1089(.a(s_77), .b(gate27inter3), .O(gate27inter10));
  nor2  gate1090(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate1091(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate1092(.a(gate27inter12), .b(gate27inter1), .O(G320));

  xor2  gate1751(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate1752(.a(gate28inter0), .b(s_172), .O(gate28inter1));
  and2  gate1753(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate1754(.a(s_172), .O(gate28inter3));
  inv1  gate1755(.a(s_173), .O(gate28inter4));
  nand2 gate1756(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate1757(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate1758(.a(G10), .O(gate28inter7));
  inv1  gate1759(.a(G14), .O(gate28inter8));
  nand2 gate1760(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate1761(.a(s_173), .b(gate28inter3), .O(gate28inter10));
  nor2  gate1762(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate1763(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate1764(.a(gate28inter12), .b(gate28inter1), .O(G323));
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate1849(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1850(.a(gate36inter0), .b(s_186), .O(gate36inter1));
  and2  gate1851(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1852(.a(s_186), .O(gate36inter3));
  inv1  gate1853(.a(s_187), .O(gate36inter4));
  nand2 gate1854(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1855(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1856(.a(G26), .O(gate36inter7));
  inv1  gate1857(.a(G30), .O(gate36inter8));
  nand2 gate1858(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1859(.a(s_187), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1860(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1861(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1862(.a(gate36inter12), .b(gate36inter1), .O(G347));

  xor2  gate1793(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate1794(.a(gate37inter0), .b(s_178), .O(gate37inter1));
  and2  gate1795(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate1796(.a(s_178), .O(gate37inter3));
  inv1  gate1797(.a(s_179), .O(gate37inter4));
  nand2 gate1798(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate1799(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate1800(.a(G19), .O(gate37inter7));
  inv1  gate1801(.a(G23), .O(gate37inter8));
  nand2 gate1802(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate1803(.a(s_179), .b(gate37inter3), .O(gate37inter10));
  nor2  gate1804(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate1805(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate1806(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate2507(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate2508(.a(gate39inter0), .b(s_280), .O(gate39inter1));
  and2  gate2509(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate2510(.a(s_280), .O(gate39inter3));
  inv1  gate2511(.a(s_281), .O(gate39inter4));
  nand2 gate2512(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate2513(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate2514(.a(G20), .O(gate39inter7));
  inv1  gate2515(.a(G24), .O(gate39inter8));
  nand2 gate2516(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate2517(.a(s_281), .b(gate39inter3), .O(gate39inter10));
  nor2  gate2518(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate2519(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate2520(.a(gate39inter12), .b(gate39inter1), .O(G356));

  xor2  gate1163(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate1164(.a(gate40inter0), .b(s_88), .O(gate40inter1));
  and2  gate1165(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate1166(.a(s_88), .O(gate40inter3));
  inv1  gate1167(.a(s_89), .O(gate40inter4));
  nand2 gate1168(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate1169(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate1170(.a(G28), .O(gate40inter7));
  inv1  gate1171(.a(G32), .O(gate40inter8));
  nand2 gate1172(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate1173(.a(s_89), .b(gate40inter3), .O(gate40inter10));
  nor2  gate1174(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate1175(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate1176(.a(gate40inter12), .b(gate40inter1), .O(G359));
nand2 gate41( .a(G1), .b(G266), .O(G362) );

  xor2  gate1275(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate1276(.a(gate42inter0), .b(s_104), .O(gate42inter1));
  and2  gate1277(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate1278(.a(s_104), .O(gate42inter3));
  inv1  gate1279(.a(s_105), .O(gate42inter4));
  nand2 gate1280(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate1281(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate1282(.a(G2), .O(gate42inter7));
  inv1  gate1283(.a(G266), .O(gate42inter8));
  nand2 gate1284(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate1285(.a(s_105), .b(gate42inter3), .O(gate42inter10));
  nor2  gate1286(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate1287(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate1288(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate2549(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate2550(.a(gate44inter0), .b(s_286), .O(gate44inter1));
  and2  gate2551(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate2552(.a(s_286), .O(gate44inter3));
  inv1  gate2553(.a(s_287), .O(gate44inter4));
  nand2 gate2554(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate2555(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate2556(.a(G4), .O(gate44inter7));
  inv1  gate2557(.a(G269), .O(gate44inter8));
  nand2 gate2558(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate2559(.a(s_287), .b(gate44inter3), .O(gate44inter10));
  nor2  gate2560(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate2561(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate2562(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );

  xor2  gate1135(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate1136(.a(gate47inter0), .b(s_84), .O(gate47inter1));
  and2  gate1137(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate1138(.a(s_84), .O(gate47inter3));
  inv1  gate1139(.a(s_85), .O(gate47inter4));
  nand2 gate1140(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate1141(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate1142(.a(G7), .O(gate47inter7));
  inv1  gate1143(.a(G275), .O(gate47inter8));
  nand2 gate1144(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate1145(.a(s_85), .b(gate47inter3), .O(gate47inter10));
  nor2  gate1146(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate1147(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate1148(.a(gate47inter12), .b(gate47inter1), .O(G368));
nand2 gate48( .a(G8), .b(G275), .O(G369) );

  xor2  gate1891(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate1892(.a(gate49inter0), .b(s_192), .O(gate49inter1));
  and2  gate1893(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate1894(.a(s_192), .O(gate49inter3));
  inv1  gate1895(.a(s_193), .O(gate49inter4));
  nand2 gate1896(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate1897(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate1898(.a(G9), .O(gate49inter7));
  inv1  gate1899(.a(G278), .O(gate49inter8));
  nand2 gate1900(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate1901(.a(s_193), .b(gate49inter3), .O(gate49inter10));
  nor2  gate1902(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate1903(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate1904(.a(gate49inter12), .b(gate49inter1), .O(G370));
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate2521(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate2522(.a(gate52inter0), .b(s_282), .O(gate52inter1));
  and2  gate2523(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate2524(.a(s_282), .O(gate52inter3));
  inv1  gate2525(.a(s_283), .O(gate52inter4));
  nand2 gate2526(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate2527(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate2528(.a(G12), .O(gate52inter7));
  inv1  gate2529(.a(G281), .O(gate52inter8));
  nand2 gate2530(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate2531(.a(s_283), .b(gate52inter3), .O(gate52inter10));
  nor2  gate2532(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate2533(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate2534(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate2017(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate2018(.a(gate54inter0), .b(s_210), .O(gate54inter1));
  and2  gate2019(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate2020(.a(s_210), .O(gate54inter3));
  inv1  gate2021(.a(s_211), .O(gate54inter4));
  nand2 gate2022(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate2023(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate2024(.a(G14), .O(gate54inter7));
  inv1  gate2025(.a(G284), .O(gate54inter8));
  nand2 gate2026(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate2027(.a(s_211), .b(gate54inter3), .O(gate54inter10));
  nor2  gate2028(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate2029(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate2030(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate995(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate996(.a(gate58inter0), .b(s_64), .O(gate58inter1));
  and2  gate997(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate998(.a(s_64), .O(gate58inter3));
  inv1  gate999(.a(s_65), .O(gate58inter4));
  nand2 gate1000(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate1001(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate1002(.a(G18), .O(gate58inter7));
  inv1  gate1003(.a(G290), .O(gate58inter8));
  nand2 gate1004(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate1005(.a(s_65), .b(gate58inter3), .O(gate58inter10));
  nor2  gate1006(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate1007(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate1008(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );

  xor2  gate2241(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate2242(.a(gate61inter0), .b(s_242), .O(gate61inter1));
  and2  gate2243(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate2244(.a(s_242), .O(gate61inter3));
  inv1  gate2245(.a(s_243), .O(gate61inter4));
  nand2 gate2246(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate2247(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate2248(.a(G21), .O(gate61inter7));
  inv1  gate2249(.a(G296), .O(gate61inter8));
  nand2 gate2250(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate2251(.a(s_243), .b(gate61inter3), .O(gate61inter10));
  nor2  gate2252(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate2253(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate2254(.a(gate61inter12), .b(gate61inter1), .O(G382));

  xor2  gate785(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate786(.a(gate62inter0), .b(s_34), .O(gate62inter1));
  and2  gate787(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate788(.a(s_34), .O(gate62inter3));
  inv1  gate789(.a(s_35), .O(gate62inter4));
  nand2 gate790(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate791(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate792(.a(G22), .O(gate62inter7));
  inv1  gate793(.a(G296), .O(gate62inter8));
  nand2 gate794(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate795(.a(s_35), .b(gate62inter3), .O(gate62inter10));
  nor2  gate796(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate797(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate798(.a(gate62inter12), .b(gate62inter1), .O(G383));

  xor2  gate1975(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate1976(.a(gate63inter0), .b(s_204), .O(gate63inter1));
  and2  gate1977(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate1978(.a(s_204), .O(gate63inter3));
  inv1  gate1979(.a(s_205), .O(gate63inter4));
  nand2 gate1980(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate1981(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate1982(.a(G23), .O(gate63inter7));
  inv1  gate1983(.a(G299), .O(gate63inter8));
  nand2 gate1984(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate1985(.a(s_205), .b(gate63inter3), .O(gate63inter10));
  nor2  gate1986(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate1987(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate1988(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate1331(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate1332(.a(gate65inter0), .b(s_112), .O(gate65inter1));
  and2  gate1333(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate1334(.a(s_112), .O(gate65inter3));
  inv1  gate1335(.a(s_113), .O(gate65inter4));
  nand2 gate1336(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate1337(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate1338(.a(G25), .O(gate65inter7));
  inv1  gate1339(.a(G302), .O(gate65inter8));
  nand2 gate1340(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate1341(.a(s_113), .b(gate65inter3), .O(gate65inter10));
  nor2  gate1342(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate1343(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate1344(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate2563(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate2564(.a(gate67inter0), .b(s_288), .O(gate67inter1));
  and2  gate2565(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate2566(.a(s_288), .O(gate67inter3));
  inv1  gate2567(.a(s_289), .O(gate67inter4));
  nand2 gate2568(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate2569(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate2570(.a(G27), .O(gate67inter7));
  inv1  gate2571(.a(G305), .O(gate67inter8));
  nand2 gate2572(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate2573(.a(s_289), .b(gate67inter3), .O(gate67inter10));
  nor2  gate2574(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate2575(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate2576(.a(gate67inter12), .b(gate67inter1), .O(G388));

  xor2  gate1037(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate1038(.a(gate68inter0), .b(s_70), .O(gate68inter1));
  and2  gate1039(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate1040(.a(s_70), .O(gate68inter3));
  inv1  gate1041(.a(s_71), .O(gate68inter4));
  nand2 gate1042(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate1043(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate1044(.a(G28), .O(gate68inter7));
  inv1  gate1045(.a(G305), .O(gate68inter8));
  nand2 gate1046(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate1047(.a(s_71), .b(gate68inter3), .O(gate68inter10));
  nor2  gate1048(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate1049(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate1050(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate2255(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate2256(.a(gate70inter0), .b(s_244), .O(gate70inter1));
  and2  gate2257(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate2258(.a(s_244), .O(gate70inter3));
  inv1  gate2259(.a(s_245), .O(gate70inter4));
  nand2 gate2260(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate2261(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate2262(.a(G30), .O(gate70inter7));
  inv1  gate2263(.a(G308), .O(gate70inter8));
  nand2 gate2264(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate2265(.a(s_245), .b(gate70inter3), .O(gate70inter10));
  nor2  gate2266(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate2267(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate2268(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );

  xor2  gate631(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate632(.a(gate72inter0), .b(s_12), .O(gate72inter1));
  and2  gate633(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate634(.a(s_12), .O(gate72inter3));
  inv1  gate635(.a(s_13), .O(gate72inter4));
  nand2 gate636(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate637(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate638(.a(G32), .O(gate72inter7));
  inv1  gate639(.a(G311), .O(gate72inter8));
  nand2 gate640(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate641(.a(s_13), .b(gate72inter3), .O(gate72inter10));
  nor2  gate642(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate643(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate644(.a(gate72inter12), .b(gate72inter1), .O(G393));
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate2143(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate2144(.a(gate75inter0), .b(s_228), .O(gate75inter1));
  and2  gate2145(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate2146(.a(s_228), .O(gate75inter3));
  inv1  gate2147(.a(s_229), .O(gate75inter4));
  nand2 gate2148(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate2149(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate2150(.a(G9), .O(gate75inter7));
  inv1  gate2151(.a(G317), .O(gate75inter8));
  nand2 gate2152(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate2153(.a(s_229), .b(gate75inter3), .O(gate75inter10));
  nor2  gate2154(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate2155(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate2156(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate855(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate856(.a(gate78inter0), .b(s_44), .O(gate78inter1));
  and2  gate857(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate858(.a(s_44), .O(gate78inter3));
  inv1  gate859(.a(s_45), .O(gate78inter4));
  nand2 gate860(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate861(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate862(.a(G6), .O(gate78inter7));
  inv1  gate863(.a(G320), .O(gate78inter8));
  nand2 gate864(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate865(.a(s_45), .b(gate78inter3), .O(gate78inter10));
  nor2  gate866(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate867(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate868(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate869(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate870(.a(gate81inter0), .b(s_46), .O(gate81inter1));
  and2  gate871(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate872(.a(s_46), .O(gate81inter3));
  inv1  gate873(.a(s_47), .O(gate81inter4));
  nand2 gate874(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate875(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate876(.a(G3), .O(gate81inter7));
  inv1  gate877(.a(G326), .O(gate81inter8));
  nand2 gate878(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate879(.a(s_47), .b(gate81inter3), .O(gate81inter10));
  nor2  gate880(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate881(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate882(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );

  xor2  gate1485(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate1486(.a(gate83inter0), .b(s_134), .O(gate83inter1));
  and2  gate1487(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate1488(.a(s_134), .O(gate83inter3));
  inv1  gate1489(.a(s_135), .O(gate83inter4));
  nand2 gate1490(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate1491(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate1492(.a(G11), .O(gate83inter7));
  inv1  gate1493(.a(G329), .O(gate83inter8));
  nand2 gate1494(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate1495(.a(s_135), .b(gate83inter3), .O(gate83inter10));
  nor2  gate1496(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate1497(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate1498(.a(gate83inter12), .b(gate83inter1), .O(G404));

  xor2  gate827(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate828(.a(gate84inter0), .b(s_40), .O(gate84inter1));
  and2  gate829(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate830(.a(s_40), .O(gate84inter3));
  inv1  gate831(.a(s_41), .O(gate84inter4));
  nand2 gate832(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate833(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate834(.a(G15), .O(gate84inter7));
  inv1  gate835(.a(G329), .O(gate84inter8));
  nand2 gate836(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate837(.a(s_41), .b(gate84inter3), .O(gate84inter10));
  nor2  gate838(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate839(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate840(.a(gate84inter12), .b(gate84inter1), .O(G405));
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate1863(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate1864(.a(gate86inter0), .b(s_188), .O(gate86inter1));
  and2  gate1865(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate1866(.a(s_188), .O(gate86inter3));
  inv1  gate1867(.a(s_189), .O(gate86inter4));
  nand2 gate1868(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate1869(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate1870(.a(G8), .O(gate86inter7));
  inv1  gate1871(.a(G332), .O(gate86inter8));
  nand2 gate1872(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate1873(.a(s_189), .b(gate86inter3), .O(gate86inter10));
  nor2  gate1874(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate1875(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate1876(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate547(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate548(.a(gate88inter0), .b(s_0), .O(gate88inter1));
  and2  gate549(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate550(.a(s_0), .O(gate88inter3));
  inv1  gate551(.a(s_1), .O(gate88inter4));
  nand2 gate552(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate553(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate554(.a(G16), .O(gate88inter7));
  inv1  gate555(.a(G335), .O(gate88inter8));
  nand2 gate556(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate557(.a(s_1), .b(gate88inter3), .O(gate88inter10));
  nor2  gate558(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate559(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate560(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate2381(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate2382(.a(gate94inter0), .b(s_262), .O(gate94inter1));
  and2  gate2383(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate2384(.a(s_262), .O(gate94inter3));
  inv1  gate2385(.a(s_263), .O(gate94inter4));
  nand2 gate2386(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate2387(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate2388(.a(G22), .O(gate94inter7));
  inv1  gate2389(.a(G344), .O(gate94inter8));
  nand2 gate2390(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate2391(.a(s_263), .b(gate94inter3), .O(gate94inter10));
  nor2  gate2392(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate2393(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate2394(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );

  xor2  gate1765(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate1766(.a(gate97inter0), .b(s_174), .O(gate97inter1));
  and2  gate1767(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate1768(.a(s_174), .O(gate97inter3));
  inv1  gate1769(.a(s_175), .O(gate97inter4));
  nand2 gate1770(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate1771(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate1772(.a(G19), .O(gate97inter7));
  inv1  gate1773(.a(G350), .O(gate97inter8));
  nand2 gate1774(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate1775(.a(s_175), .b(gate97inter3), .O(gate97inter10));
  nor2  gate1776(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate1777(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate1778(.a(gate97inter12), .b(gate97inter1), .O(G418));
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );

  xor2  gate1555(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate1556(.a(gate101inter0), .b(s_144), .O(gate101inter1));
  and2  gate1557(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate1558(.a(s_144), .O(gate101inter3));
  inv1  gate1559(.a(s_145), .O(gate101inter4));
  nand2 gate1560(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate1561(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate1562(.a(G20), .O(gate101inter7));
  inv1  gate1563(.a(G356), .O(gate101inter8));
  nand2 gate1564(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate1565(.a(s_145), .b(gate101inter3), .O(gate101inter10));
  nor2  gate1566(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate1567(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate1568(.a(gate101inter12), .b(gate101inter1), .O(G422));
nand2 gate102( .a(G24), .b(G356), .O(G423) );

  xor2  gate2577(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate2578(.a(gate103inter0), .b(s_290), .O(gate103inter1));
  and2  gate2579(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate2580(.a(s_290), .O(gate103inter3));
  inv1  gate2581(.a(s_291), .O(gate103inter4));
  nand2 gate2582(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate2583(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate2584(.a(G28), .O(gate103inter7));
  inv1  gate2585(.a(G359), .O(gate103inter8));
  nand2 gate2586(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate2587(.a(s_291), .b(gate103inter3), .O(gate103inter10));
  nor2  gate2588(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate2589(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate2590(.a(gate103inter12), .b(gate103inter1), .O(G424));
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate2451(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate2452(.a(gate108inter0), .b(s_272), .O(gate108inter1));
  and2  gate2453(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate2454(.a(s_272), .O(gate108inter3));
  inv1  gate2455(.a(s_273), .O(gate108inter4));
  nand2 gate2456(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate2457(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate2458(.a(G368), .O(gate108inter7));
  inv1  gate2459(.a(G369), .O(gate108inter8));
  nand2 gate2460(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate2461(.a(s_273), .b(gate108inter3), .O(gate108inter10));
  nor2  gate2462(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate2463(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate2464(.a(gate108inter12), .b(gate108inter1), .O(G435));
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );

  xor2  gate2115(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate2116(.a(gate114inter0), .b(s_224), .O(gate114inter1));
  and2  gate2117(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate2118(.a(s_224), .O(gate114inter3));
  inv1  gate2119(.a(s_225), .O(gate114inter4));
  nand2 gate2120(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate2121(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate2122(.a(G380), .O(gate114inter7));
  inv1  gate2123(.a(G381), .O(gate114inter8));
  nand2 gate2124(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate2125(.a(s_225), .b(gate114inter3), .O(gate114inter10));
  nor2  gate2126(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate2127(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate2128(.a(gate114inter12), .b(gate114inter1), .O(G453));

  xor2  gate911(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate912(.a(gate115inter0), .b(s_52), .O(gate115inter1));
  and2  gate913(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate914(.a(s_52), .O(gate115inter3));
  inv1  gate915(.a(s_53), .O(gate115inter4));
  nand2 gate916(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate917(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate918(.a(G382), .O(gate115inter7));
  inv1  gate919(.a(G383), .O(gate115inter8));
  nand2 gate920(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate921(.a(s_53), .b(gate115inter3), .O(gate115inter10));
  nor2  gate922(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate923(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate924(.a(gate115inter12), .b(gate115inter1), .O(G456));

  xor2  gate673(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate674(.a(gate116inter0), .b(s_18), .O(gate116inter1));
  and2  gate675(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate676(.a(s_18), .O(gate116inter3));
  inv1  gate677(.a(s_19), .O(gate116inter4));
  nand2 gate678(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate679(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate680(.a(G384), .O(gate116inter7));
  inv1  gate681(.a(G385), .O(gate116inter8));
  nand2 gate682(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate683(.a(s_19), .b(gate116inter3), .O(gate116inter10));
  nor2  gate684(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate685(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate686(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate2101(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate2102(.a(gate118inter0), .b(s_222), .O(gate118inter1));
  and2  gate2103(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate2104(.a(s_222), .O(gate118inter3));
  inv1  gate2105(.a(s_223), .O(gate118inter4));
  nand2 gate2106(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate2107(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate2108(.a(G388), .O(gate118inter7));
  inv1  gate2109(.a(G389), .O(gate118inter8));
  nand2 gate2110(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate2111(.a(s_223), .b(gate118inter3), .O(gate118inter10));
  nor2  gate2112(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate2113(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate2114(.a(gate118inter12), .b(gate118inter1), .O(G465));
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate1429(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate1430(.a(gate124inter0), .b(s_126), .O(gate124inter1));
  and2  gate1431(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate1432(.a(s_126), .O(gate124inter3));
  inv1  gate1433(.a(s_127), .O(gate124inter4));
  nand2 gate1434(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate1435(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate1436(.a(G400), .O(gate124inter7));
  inv1  gate1437(.a(G401), .O(gate124inter8));
  nand2 gate1438(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate1439(.a(s_127), .b(gate124inter3), .O(gate124inter10));
  nor2  gate1440(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate1441(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate1442(.a(gate124inter12), .b(gate124inter1), .O(G483));

  xor2  gate2199(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate2200(.a(gate125inter0), .b(s_236), .O(gate125inter1));
  and2  gate2201(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate2202(.a(s_236), .O(gate125inter3));
  inv1  gate2203(.a(s_237), .O(gate125inter4));
  nand2 gate2204(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate2205(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate2206(.a(G402), .O(gate125inter7));
  inv1  gate2207(.a(G403), .O(gate125inter8));
  nand2 gate2208(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate2209(.a(s_237), .b(gate125inter3), .O(gate125inter10));
  nor2  gate2210(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate2211(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate2212(.a(gate125inter12), .b(gate125inter1), .O(G486));

  xor2  gate2059(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate2060(.a(gate126inter0), .b(s_216), .O(gate126inter1));
  and2  gate2061(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate2062(.a(s_216), .O(gate126inter3));
  inv1  gate2063(.a(s_217), .O(gate126inter4));
  nand2 gate2064(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate2065(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate2066(.a(G404), .O(gate126inter7));
  inv1  gate2067(.a(G405), .O(gate126inter8));
  nand2 gate2068(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate2069(.a(s_217), .b(gate126inter3), .O(gate126inter10));
  nor2  gate2070(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate2071(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate2072(.a(gate126inter12), .b(gate126inter1), .O(G489));

  xor2  gate953(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate954(.a(gate127inter0), .b(s_58), .O(gate127inter1));
  and2  gate955(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate956(.a(s_58), .O(gate127inter3));
  inv1  gate957(.a(s_59), .O(gate127inter4));
  nand2 gate958(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate959(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate960(.a(G406), .O(gate127inter7));
  inv1  gate961(.a(G407), .O(gate127inter8));
  nand2 gate962(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate963(.a(s_59), .b(gate127inter3), .O(gate127inter10));
  nor2  gate964(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate965(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate966(.a(gate127inter12), .b(gate127inter1), .O(G492));

  xor2  gate2157(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate2158(.a(gate128inter0), .b(s_230), .O(gate128inter1));
  and2  gate2159(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate2160(.a(s_230), .O(gate128inter3));
  inv1  gate2161(.a(s_231), .O(gate128inter4));
  nand2 gate2162(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate2163(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate2164(.a(G408), .O(gate128inter7));
  inv1  gate2165(.a(G409), .O(gate128inter8));
  nand2 gate2166(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate2167(.a(s_231), .b(gate128inter3), .O(gate128inter10));
  nor2  gate2168(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate2169(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate2170(.a(gate128inter12), .b(gate128inter1), .O(G495));
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );

  xor2  gate1121(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate1122(.a(gate133inter0), .b(s_82), .O(gate133inter1));
  and2  gate1123(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate1124(.a(s_82), .O(gate133inter3));
  inv1  gate1125(.a(s_83), .O(gate133inter4));
  nand2 gate1126(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate1127(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate1128(.a(G418), .O(gate133inter7));
  inv1  gate1129(.a(G419), .O(gate133inter8));
  nand2 gate1130(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate1131(.a(s_83), .b(gate133inter3), .O(gate133inter10));
  nor2  gate1132(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate1133(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate1134(.a(gate133inter12), .b(gate133inter1), .O(G510));
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate1569(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate1570(.a(gate136inter0), .b(s_146), .O(gate136inter1));
  and2  gate1571(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate1572(.a(s_146), .O(gate136inter3));
  inv1  gate1573(.a(s_147), .O(gate136inter4));
  nand2 gate1574(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate1575(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate1576(.a(G424), .O(gate136inter7));
  inv1  gate1577(.a(G425), .O(gate136inter8));
  nand2 gate1578(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate1579(.a(s_147), .b(gate136inter3), .O(gate136inter10));
  nor2  gate1580(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate1581(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate1582(.a(gate136inter12), .b(gate136inter1), .O(G519));

  xor2  gate1051(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate1052(.a(gate137inter0), .b(s_72), .O(gate137inter1));
  and2  gate1053(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate1054(.a(s_72), .O(gate137inter3));
  inv1  gate1055(.a(s_73), .O(gate137inter4));
  nand2 gate1056(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate1057(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate1058(.a(G426), .O(gate137inter7));
  inv1  gate1059(.a(G429), .O(gate137inter8));
  nand2 gate1060(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate1061(.a(s_73), .b(gate137inter3), .O(gate137inter10));
  nor2  gate1062(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate1063(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate1064(.a(gate137inter12), .b(gate137inter1), .O(G522));

  xor2  gate771(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate772(.a(gate138inter0), .b(s_32), .O(gate138inter1));
  and2  gate773(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate774(.a(s_32), .O(gate138inter3));
  inv1  gate775(.a(s_33), .O(gate138inter4));
  nand2 gate776(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate777(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate778(.a(G432), .O(gate138inter7));
  inv1  gate779(.a(G435), .O(gate138inter8));
  nand2 gate780(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate781(.a(s_33), .b(gate138inter3), .O(gate138inter10));
  nor2  gate782(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate783(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate784(.a(gate138inter12), .b(gate138inter1), .O(G525));

  xor2  gate2479(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate2480(.a(gate139inter0), .b(s_276), .O(gate139inter1));
  and2  gate2481(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate2482(.a(s_276), .O(gate139inter3));
  inv1  gate2483(.a(s_277), .O(gate139inter4));
  nand2 gate2484(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate2485(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate2486(.a(G438), .O(gate139inter7));
  inv1  gate2487(.a(G441), .O(gate139inter8));
  nand2 gate2488(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate2489(.a(s_277), .b(gate139inter3), .O(gate139inter10));
  nor2  gate2490(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate2491(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate2492(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate1359(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate1360(.a(gate142inter0), .b(s_116), .O(gate142inter1));
  and2  gate1361(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate1362(.a(s_116), .O(gate142inter3));
  inv1  gate1363(.a(s_117), .O(gate142inter4));
  nand2 gate1364(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate1365(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate1366(.a(G456), .O(gate142inter7));
  inv1  gate1367(.a(G459), .O(gate142inter8));
  nand2 gate1368(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate1369(.a(s_117), .b(gate142inter3), .O(gate142inter10));
  nor2  gate1370(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate1371(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate1372(.a(gate142inter12), .b(gate142inter1), .O(G537));
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );

  xor2  gate2031(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate2032(.a(gate145inter0), .b(s_212), .O(gate145inter1));
  and2  gate2033(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate2034(.a(s_212), .O(gate145inter3));
  inv1  gate2035(.a(s_213), .O(gate145inter4));
  nand2 gate2036(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate2037(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate2038(.a(G474), .O(gate145inter7));
  inv1  gate2039(.a(G477), .O(gate145inter8));
  nand2 gate2040(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate2041(.a(s_213), .b(gate145inter3), .O(gate145inter10));
  nor2  gate2042(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate2043(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate2044(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate1191(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate1192(.a(gate153inter0), .b(s_92), .O(gate153inter1));
  and2  gate1193(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate1194(.a(s_92), .O(gate153inter3));
  inv1  gate1195(.a(s_93), .O(gate153inter4));
  nand2 gate1196(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate1197(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate1198(.a(G426), .O(gate153inter7));
  inv1  gate1199(.a(G522), .O(gate153inter8));
  nand2 gate1200(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate1201(.a(s_93), .b(gate153inter3), .O(gate153inter10));
  nor2  gate1202(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate1203(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate1204(.a(gate153inter12), .b(gate153inter1), .O(G570));
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate1065(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate1066(.a(gate156inter0), .b(s_74), .O(gate156inter1));
  and2  gate1067(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate1068(.a(s_74), .O(gate156inter3));
  inv1  gate1069(.a(s_75), .O(gate156inter4));
  nand2 gate1070(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate1071(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate1072(.a(G435), .O(gate156inter7));
  inv1  gate1073(.a(G525), .O(gate156inter8));
  nand2 gate1074(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate1075(.a(s_75), .b(gate156inter3), .O(gate156inter10));
  nor2  gate1076(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate1077(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate1078(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate1989(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate1990(.a(gate159inter0), .b(s_206), .O(gate159inter1));
  and2  gate1991(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate1992(.a(s_206), .O(gate159inter3));
  inv1  gate1993(.a(s_207), .O(gate159inter4));
  nand2 gate1994(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate1995(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate1996(.a(G444), .O(gate159inter7));
  inv1  gate1997(.a(G531), .O(gate159inter8));
  nand2 gate1998(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate1999(.a(s_207), .b(gate159inter3), .O(gate159inter10));
  nor2  gate2000(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate2001(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate2002(.a(gate159inter12), .b(gate159inter1), .O(G576));

  xor2  gate687(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate688(.a(gate160inter0), .b(s_20), .O(gate160inter1));
  and2  gate689(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate690(.a(s_20), .O(gate160inter3));
  inv1  gate691(.a(s_21), .O(gate160inter4));
  nand2 gate692(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate693(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate694(.a(G447), .O(gate160inter7));
  inv1  gate695(.a(G531), .O(gate160inter8));
  nand2 gate696(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate697(.a(s_21), .b(gate160inter3), .O(gate160inter10));
  nor2  gate698(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate699(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate700(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate2171(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate2172(.a(gate162inter0), .b(s_232), .O(gate162inter1));
  and2  gate2173(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate2174(.a(s_232), .O(gate162inter3));
  inv1  gate2175(.a(s_233), .O(gate162inter4));
  nand2 gate2176(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate2177(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate2178(.a(G453), .O(gate162inter7));
  inv1  gate2179(.a(G534), .O(gate162inter8));
  nand2 gate2180(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate2181(.a(s_233), .b(gate162inter3), .O(gate162inter10));
  nor2  gate2182(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate2183(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate2184(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );

  xor2  gate1443(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate1444(.a(gate167inter0), .b(s_128), .O(gate167inter1));
  and2  gate1445(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate1446(.a(s_128), .O(gate167inter3));
  inv1  gate1447(.a(s_129), .O(gate167inter4));
  nand2 gate1448(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate1449(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate1450(.a(G468), .O(gate167inter7));
  inv1  gate1451(.a(G543), .O(gate167inter8));
  nand2 gate1452(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate1453(.a(s_129), .b(gate167inter3), .O(gate167inter10));
  nor2  gate1454(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate1455(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate1456(.a(gate167inter12), .b(gate167inter1), .O(G584));
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate589(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate590(.a(gate172inter0), .b(s_6), .O(gate172inter1));
  and2  gate591(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate592(.a(s_6), .O(gate172inter3));
  inv1  gate593(.a(s_7), .O(gate172inter4));
  nand2 gate594(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate595(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate596(.a(G483), .O(gate172inter7));
  inv1  gate597(.a(G549), .O(gate172inter8));
  nand2 gate598(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate599(.a(s_7), .b(gate172inter3), .O(gate172inter10));
  nor2  gate600(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate601(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate602(.a(gate172inter12), .b(gate172inter1), .O(G589));

  xor2  gate1387(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate1388(.a(gate173inter0), .b(s_120), .O(gate173inter1));
  and2  gate1389(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate1390(.a(s_120), .O(gate173inter3));
  inv1  gate1391(.a(s_121), .O(gate173inter4));
  nand2 gate1392(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate1393(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate1394(.a(G486), .O(gate173inter7));
  inv1  gate1395(.a(G552), .O(gate173inter8));
  nand2 gate1396(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate1397(.a(s_121), .b(gate173inter3), .O(gate173inter10));
  nor2  gate1398(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate1399(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate1400(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );

  xor2  gate1247(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate1248(.a(gate176inter0), .b(s_100), .O(gate176inter1));
  and2  gate1249(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate1250(.a(s_100), .O(gate176inter3));
  inv1  gate1251(.a(s_101), .O(gate176inter4));
  nand2 gate1252(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate1253(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate1254(.a(G495), .O(gate176inter7));
  inv1  gate1255(.a(G555), .O(gate176inter8));
  nand2 gate1256(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate1257(.a(s_101), .b(gate176inter3), .O(gate176inter10));
  nor2  gate1258(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate1259(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate1260(.a(gate176inter12), .b(gate176inter1), .O(G593));

  xor2  gate1695(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate1696(.a(gate177inter0), .b(s_164), .O(gate177inter1));
  and2  gate1697(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate1698(.a(s_164), .O(gate177inter3));
  inv1  gate1699(.a(s_165), .O(gate177inter4));
  nand2 gate1700(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate1701(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate1702(.a(G498), .O(gate177inter7));
  inv1  gate1703(.a(G558), .O(gate177inter8));
  nand2 gate1704(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate1705(.a(s_165), .b(gate177inter3), .O(gate177inter10));
  nor2  gate1706(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate1707(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate1708(.a(gate177inter12), .b(gate177inter1), .O(G594));
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate659(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate660(.a(gate180inter0), .b(s_16), .O(gate180inter1));
  and2  gate661(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate662(.a(s_16), .O(gate180inter3));
  inv1  gate663(.a(s_17), .O(gate180inter4));
  nand2 gate664(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate665(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate666(.a(G507), .O(gate180inter7));
  inv1  gate667(.a(G561), .O(gate180inter8));
  nand2 gate668(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate669(.a(s_17), .b(gate180inter3), .O(gate180inter10));
  nor2  gate670(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate671(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate672(.a(gate180inter12), .b(gate180inter1), .O(G597));

  xor2  gate1541(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate1542(.a(gate181inter0), .b(s_142), .O(gate181inter1));
  and2  gate1543(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate1544(.a(s_142), .O(gate181inter3));
  inv1  gate1545(.a(s_143), .O(gate181inter4));
  nand2 gate1546(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate1547(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate1548(.a(G510), .O(gate181inter7));
  inv1  gate1549(.a(G564), .O(gate181inter8));
  nand2 gate1550(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate1551(.a(s_143), .b(gate181inter3), .O(gate181inter10));
  nor2  gate1552(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate1553(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate1554(.a(gate181inter12), .b(gate181inter1), .O(G598));
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate1289(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1290(.a(gate186inter0), .b(s_106), .O(gate186inter1));
  and2  gate1291(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1292(.a(s_106), .O(gate186inter3));
  inv1  gate1293(.a(s_107), .O(gate186inter4));
  nand2 gate1294(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1295(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1296(.a(G572), .O(gate186inter7));
  inv1  gate1297(.a(G573), .O(gate186inter8));
  nand2 gate1298(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1299(.a(s_107), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1300(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1301(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1302(.a(gate186inter12), .b(gate186inter1), .O(G607));

  xor2  gate1023(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate1024(.a(gate187inter0), .b(s_68), .O(gate187inter1));
  and2  gate1025(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate1026(.a(s_68), .O(gate187inter3));
  inv1  gate1027(.a(s_69), .O(gate187inter4));
  nand2 gate1028(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate1029(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate1030(.a(G574), .O(gate187inter7));
  inv1  gate1031(.a(G575), .O(gate187inter8));
  nand2 gate1032(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate1033(.a(s_69), .b(gate187inter3), .O(gate187inter10));
  nor2  gate1034(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate1035(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate1036(.a(gate187inter12), .b(gate187inter1), .O(G612));
nand2 gate188( .a(G576), .b(G577), .O(G617) );

  xor2  gate2311(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate2312(.a(gate189inter0), .b(s_252), .O(gate189inter1));
  and2  gate2313(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate2314(.a(s_252), .O(gate189inter3));
  inv1  gate2315(.a(s_253), .O(gate189inter4));
  nand2 gate2316(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate2317(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate2318(.a(G578), .O(gate189inter7));
  inv1  gate2319(.a(G579), .O(gate189inter8));
  nand2 gate2320(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate2321(.a(s_253), .b(gate189inter3), .O(gate189inter10));
  nor2  gate2322(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate2323(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate2324(.a(gate189inter12), .b(gate189inter1), .O(G622));

  xor2  gate1177(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate1178(.a(gate190inter0), .b(s_90), .O(gate190inter1));
  and2  gate1179(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate1180(.a(s_90), .O(gate190inter3));
  inv1  gate1181(.a(s_91), .O(gate190inter4));
  nand2 gate1182(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate1183(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate1184(.a(G580), .O(gate190inter7));
  inv1  gate1185(.a(G581), .O(gate190inter8));
  nand2 gate1186(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate1187(.a(s_91), .b(gate190inter3), .O(gate190inter10));
  nor2  gate1188(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate1189(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate1190(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );

  xor2  gate561(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate562(.a(gate192inter0), .b(s_2), .O(gate192inter1));
  and2  gate563(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate564(.a(s_2), .O(gate192inter3));
  inv1  gate565(.a(s_3), .O(gate192inter4));
  nand2 gate566(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate567(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate568(.a(G584), .O(gate192inter7));
  inv1  gate569(.a(G585), .O(gate192inter8));
  nand2 gate570(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate571(.a(s_3), .b(gate192inter3), .O(gate192inter10));
  nor2  gate572(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate573(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate574(.a(gate192inter12), .b(gate192inter1), .O(G637));

  xor2  gate1373(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate1374(.a(gate193inter0), .b(s_118), .O(gate193inter1));
  and2  gate1375(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate1376(.a(s_118), .O(gate193inter3));
  inv1  gate1377(.a(s_119), .O(gate193inter4));
  nand2 gate1378(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate1379(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate1380(.a(G586), .O(gate193inter7));
  inv1  gate1381(.a(G587), .O(gate193inter8));
  nand2 gate1382(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate1383(.a(s_119), .b(gate193inter3), .O(gate193inter10));
  nor2  gate1384(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate1385(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate1386(.a(gate193inter12), .b(gate193inter1), .O(G642));

  xor2  gate1877(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate1878(.a(gate194inter0), .b(s_190), .O(gate194inter1));
  and2  gate1879(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate1880(.a(s_190), .O(gate194inter3));
  inv1  gate1881(.a(s_191), .O(gate194inter4));
  nand2 gate1882(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate1883(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate1884(.a(G588), .O(gate194inter7));
  inv1  gate1885(.a(G589), .O(gate194inter8));
  nand2 gate1886(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate1887(.a(s_191), .b(gate194inter3), .O(gate194inter10));
  nor2  gate1888(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate1889(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate1890(.a(gate194inter12), .b(gate194inter1), .O(G645));
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate575(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate576(.a(gate201inter0), .b(s_4), .O(gate201inter1));
  and2  gate577(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate578(.a(s_4), .O(gate201inter3));
  inv1  gate579(.a(s_5), .O(gate201inter4));
  nand2 gate580(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate581(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate582(.a(G602), .O(gate201inter7));
  inv1  gate583(.a(G607), .O(gate201inter8));
  nand2 gate584(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate585(.a(s_5), .b(gate201inter3), .O(gate201inter10));
  nor2  gate586(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate587(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate588(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );

  xor2  gate2465(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate2466(.a(gate204inter0), .b(s_274), .O(gate204inter1));
  and2  gate2467(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate2468(.a(s_274), .O(gate204inter3));
  inv1  gate2469(.a(s_275), .O(gate204inter4));
  nand2 gate2470(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate2471(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate2472(.a(G607), .O(gate204inter7));
  inv1  gate2473(.a(G617), .O(gate204inter8));
  nand2 gate2474(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate2475(.a(s_275), .b(gate204inter3), .O(gate204inter10));
  nor2  gate2476(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate2477(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate2478(.a(gate204inter12), .b(gate204inter1), .O(G675));
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );

  xor2  gate1919(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate1920(.a(gate207inter0), .b(s_196), .O(gate207inter1));
  and2  gate1921(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate1922(.a(s_196), .O(gate207inter3));
  inv1  gate1923(.a(s_197), .O(gate207inter4));
  nand2 gate1924(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate1925(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate1926(.a(G622), .O(gate207inter7));
  inv1  gate1927(.a(G632), .O(gate207inter8));
  nand2 gate1928(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate1929(.a(s_197), .b(gate207inter3), .O(gate207inter10));
  nor2  gate1930(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate1931(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate1932(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );

  xor2  gate1219(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate1220(.a(gate209inter0), .b(s_96), .O(gate209inter1));
  and2  gate1221(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate1222(.a(s_96), .O(gate209inter3));
  inv1  gate1223(.a(s_97), .O(gate209inter4));
  nand2 gate1224(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate1225(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate1226(.a(G602), .O(gate209inter7));
  inv1  gate1227(.a(G666), .O(gate209inter8));
  nand2 gate1228(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate1229(.a(s_97), .b(gate209inter3), .O(gate209inter10));
  nor2  gate1230(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate1231(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate1232(.a(gate209inter12), .b(gate209inter1), .O(G690));
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate1653(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate1654(.a(gate211inter0), .b(s_158), .O(gate211inter1));
  and2  gate1655(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate1656(.a(s_158), .O(gate211inter3));
  inv1  gate1657(.a(s_159), .O(gate211inter4));
  nand2 gate1658(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate1659(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate1660(.a(G612), .O(gate211inter7));
  inv1  gate1661(.a(G669), .O(gate211inter8));
  nand2 gate1662(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate1663(.a(s_159), .b(gate211inter3), .O(gate211inter10));
  nor2  gate1664(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate1665(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate1666(.a(gate211inter12), .b(gate211inter1), .O(G692));
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate617(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate618(.a(gate213inter0), .b(s_10), .O(gate213inter1));
  and2  gate619(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate620(.a(s_10), .O(gate213inter3));
  inv1  gate621(.a(s_11), .O(gate213inter4));
  nand2 gate622(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate623(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate624(.a(G602), .O(gate213inter7));
  inv1  gate625(.a(G672), .O(gate213inter8));
  nand2 gate626(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate627(.a(s_11), .b(gate213inter3), .O(gate213inter10));
  nor2  gate628(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate629(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate630(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate1961(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate1962(.a(gate215inter0), .b(s_202), .O(gate215inter1));
  and2  gate1963(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate1964(.a(s_202), .O(gate215inter3));
  inv1  gate1965(.a(s_203), .O(gate215inter4));
  nand2 gate1966(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate1967(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate1968(.a(G607), .O(gate215inter7));
  inv1  gate1969(.a(G675), .O(gate215inter8));
  nand2 gate1970(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate1971(.a(s_203), .b(gate215inter3), .O(gate215inter10));
  nor2  gate1972(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate1973(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate1974(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );

  xor2  gate841(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate842(.a(gate217inter0), .b(s_42), .O(gate217inter1));
  and2  gate843(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate844(.a(s_42), .O(gate217inter3));
  inv1  gate845(.a(s_43), .O(gate217inter4));
  nand2 gate846(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate847(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate848(.a(G622), .O(gate217inter7));
  inv1  gate849(.a(G678), .O(gate217inter8));
  nand2 gate850(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate851(.a(s_43), .b(gate217inter3), .O(gate217inter10));
  nor2  gate852(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate853(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate854(.a(gate217inter12), .b(gate217inter1), .O(G698));
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate925(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate926(.a(gate226inter0), .b(s_54), .O(gate226inter1));
  and2  gate927(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate928(.a(s_54), .O(gate226inter3));
  inv1  gate929(.a(s_55), .O(gate226inter4));
  nand2 gate930(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate931(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate932(.a(G692), .O(gate226inter7));
  inv1  gate933(.a(G693), .O(gate226inter8));
  nand2 gate934(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate935(.a(s_55), .b(gate226inter3), .O(gate226inter10));
  nor2  gate936(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate937(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate938(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate2325(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate2326(.a(gate228inter0), .b(s_254), .O(gate228inter1));
  and2  gate2327(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate2328(.a(s_254), .O(gate228inter3));
  inv1  gate2329(.a(s_255), .O(gate228inter4));
  nand2 gate2330(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate2331(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate2332(.a(G696), .O(gate228inter7));
  inv1  gate2333(.a(G697), .O(gate228inter8));
  nand2 gate2334(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate2335(.a(s_255), .b(gate228inter3), .O(gate228inter10));
  nor2  gate2336(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate2337(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate2338(.a(gate228inter12), .b(gate228inter1), .O(G715));

  xor2  gate883(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate884(.a(gate229inter0), .b(s_48), .O(gate229inter1));
  and2  gate885(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate886(.a(s_48), .O(gate229inter3));
  inv1  gate887(.a(s_49), .O(gate229inter4));
  nand2 gate888(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate889(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate890(.a(G698), .O(gate229inter7));
  inv1  gate891(.a(G699), .O(gate229inter8));
  nand2 gate892(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate893(.a(s_49), .b(gate229inter3), .O(gate229inter10));
  nor2  gate894(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate895(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate896(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate799(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate800(.a(gate234inter0), .b(s_36), .O(gate234inter1));
  and2  gate801(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate802(.a(s_36), .O(gate234inter3));
  inv1  gate803(.a(s_37), .O(gate234inter4));
  nand2 gate804(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate805(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate806(.a(G245), .O(gate234inter7));
  inv1  gate807(.a(G721), .O(gate234inter8));
  nand2 gate808(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate809(.a(s_37), .b(gate234inter3), .O(gate234inter10));
  nor2  gate810(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate811(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate812(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate2535(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate2536(.a(gate236inter0), .b(s_284), .O(gate236inter1));
  and2  gate2537(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate2538(.a(s_284), .O(gate236inter3));
  inv1  gate2539(.a(s_285), .O(gate236inter4));
  nand2 gate2540(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate2541(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate2542(.a(G251), .O(gate236inter7));
  inv1  gate2543(.a(G727), .O(gate236inter8));
  nand2 gate2544(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate2545(.a(s_285), .b(gate236inter3), .O(gate236inter10));
  nor2  gate2546(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate2547(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate2548(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );

  xor2  gate1821(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate1822(.a(gate244inter0), .b(s_182), .O(gate244inter1));
  and2  gate1823(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate1824(.a(s_182), .O(gate244inter3));
  inv1  gate1825(.a(s_183), .O(gate244inter4));
  nand2 gate1826(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate1827(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate1828(.a(G721), .O(gate244inter7));
  inv1  gate1829(.a(G733), .O(gate244inter8));
  nand2 gate1830(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate1831(.a(s_183), .b(gate244inter3), .O(gate244inter10));
  nor2  gate1832(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate1833(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate1834(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );

  xor2  gate603(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate604(.a(gate247inter0), .b(s_8), .O(gate247inter1));
  and2  gate605(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate606(.a(s_8), .O(gate247inter3));
  inv1  gate607(.a(s_9), .O(gate247inter4));
  nand2 gate608(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate609(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate610(.a(G251), .O(gate247inter7));
  inv1  gate611(.a(G739), .O(gate247inter8));
  nand2 gate612(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate613(.a(s_9), .b(gate247inter3), .O(gate247inter10));
  nor2  gate614(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate615(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate616(.a(gate247inter12), .b(gate247inter1), .O(G760));
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate2409(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate2410(.a(gate250inter0), .b(s_266), .O(gate250inter1));
  and2  gate2411(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate2412(.a(s_266), .O(gate250inter3));
  inv1  gate2413(.a(s_267), .O(gate250inter4));
  nand2 gate2414(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate2415(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate2416(.a(G706), .O(gate250inter7));
  inv1  gate2417(.a(G742), .O(gate250inter8));
  nand2 gate2418(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate2419(.a(s_267), .b(gate250inter3), .O(gate250inter10));
  nor2  gate2420(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate2421(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate2422(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate715(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate716(.a(gate252inter0), .b(s_24), .O(gate252inter1));
  and2  gate717(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate718(.a(s_24), .O(gate252inter3));
  inv1  gate719(.a(s_25), .O(gate252inter4));
  nand2 gate720(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate721(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate722(.a(G709), .O(gate252inter7));
  inv1  gate723(.a(G745), .O(gate252inter8));
  nand2 gate724(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate725(.a(s_25), .b(gate252inter3), .O(gate252inter10));
  nor2  gate726(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate727(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate728(.a(gate252inter12), .b(gate252inter1), .O(G765));

  xor2  gate939(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate940(.a(gate253inter0), .b(s_56), .O(gate253inter1));
  and2  gate941(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate942(.a(s_56), .O(gate253inter3));
  inv1  gate943(.a(s_57), .O(gate253inter4));
  nand2 gate944(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate945(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate946(.a(G260), .O(gate253inter7));
  inv1  gate947(.a(G748), .O(gate253inter8));
  nand2 gate948(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate949(.a(s_57), .b(gate253inter3), .O(gate253inter10));
  nor2  gate950(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate951(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate952(.a(gate253inter12), .b(gate253inter1), .O(G766));

  xor2  gate701(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate702(.a(gate254inter0), .b(s_22), .O(gate254inter1));
  and2  gate703(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate704(.a(s_22), .O(gate254inter3));
  inv1  gate705(.a(s_23), .O(gate254inter4));
  nand2 gate706(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate707(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate708(.a(G712), .O(gate254inter7));
  inv1  gate709(.a(G748), .O(gate254inter8));
  nand2 gate710(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate711(.a(s_23), .b(gate254inter3), .O(gate254inter10));
  nor2  gate712(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate713(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate714(.a(gate254inter12), .b(gate254inter1), .O(G767));
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate1807(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate1808(.a(gate257inter0), .b(s_180), .O(gate257inter1));
  and2  gate1809(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate1810(.a(s_180), .O(gate257inter3));
  inv1  gate1811(.a(s_181), .O(gate257inter4));
  nand2 gate1812(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate1813(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate1814(.a(G754), .O(gate257inter7));
  inv1  gate1815(.a(G755), .O(gate257inter8));
  nand2 gate1816(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate1817(.a(s_181), .b(gate257inter3), .O(gate257inter10));
  nor2  gate1818(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate1819(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate1820(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate2423(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate2424(.a(gate261inter0), .b(s_268), .O(gate261inter1));
  and2  gate2425(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate2426(.a(s_268), .O(gate261inter3));
  inv1  gate2427(.a(s_269), .O(gate261inter4));
  nand2 gate2428(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate2429(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate2430(.a(G762), .O(gate261inter7));
  inv1  gate2431(.a(G763), .O(gate261inter8));
  nand2 gate2432(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate2433(.a(s_269), .b(gate261inter3), .O(gate261inter10));
  nor2  gate2434(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate2435(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate2436(.a(gate261inter12), .b(gate261inter1), .O(G782));

  xor2  gate1947(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate1948(.a(gate262inter0), .b(s_200), .O(gate262inter1));
  and2  gate1949(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate1950(.a(s_200), .O(gate262inter3));
  inv1  gate1951(.a(s_201), .O(gate262inter4));
  nand2 gate1952(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate1953(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate1954(.a(G764), .O(gate262inter7));
  inv1  gate1955(.a(G765), .O(gate262inter8));
  nand2 gate1956(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate1957(.a(s_201), .b(gate262inter3), .O(gate262inter10));
  nor2  gate1958(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate1959(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate1960(.a(gate262inter12), .b(gate262inter1), .O(G785));

  xor2  gate1681(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate1682(.a(gate263inter0), .b(s_162), .O(gate263inter1));
  and2  gate1683(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate1684(.a(s_162), .O(gate263inter3));
  inv1  gate1685(.a(s_163), .O(gate263inter4));
  nand2 gate1686(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate1687(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate1688(.a(G766), .O(gate263inter7));
  inv1  gate1689(.a(G767), .O(gate263inter8));
  nand2 gate1690(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate1691(.a(s_163), .b(gate263inter3), .O(gate263inter10));
  nor2  gate1692(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate1693(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate1694(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate1261(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate1262(.a(gate266inter0), .b(s_102), .O(gate266inter1));
  and2  gate1263(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate1264(.a(s_102), .O(gate266inter3));
  inv1  gate1265(.a(s_103), .O(gate266inter4));
  nand2 gate1266(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate1267(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate1268(.a(G645), .O(gate266inter7));
  inv1  gate1269(.a(G773), .O(gate266inter8));
  nand2 gate1270(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate1271(.a(s_103), .b(gate266inter3), .O(gate266inter10));
  nor2  gate1272(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate1273(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate1274(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate1303(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate1304(.a(gate268inter0), .b(s_108), .O(gate268inter1));
  and2  gate1305(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate1306(.a(s_108), .O(gate268inter3));
  inv1  gate1307(.a(s_109), .O(gate268inter4));
  nand2 gate1308(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1309(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1310(.a(G651), .O(gate268inter7));
  inv1  gate1311(.a(G779), .O(gate268inter8));
  nand2 gate1312(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1313(.a(s_109), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1314(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1315(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1316(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate1149(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate1150(.a(gate272inter0), .b(s_86), .O(gate272inter1));
  and2  gate1151(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate1152(.a(s_86), .O(gate272inter3));
  inv1  gate1153(.a(s_87), .O(gate272inter4));
  nand2 gate1154(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate1155(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate1156(.a(G663), .O(gate272inter7));
  inv1  gate1157(.a(G791), .O(gate272inter8));
  nand2 gate1158(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate1159(.a(s_87), .b(gate272inter3), .O(gate272inter10));
  nor2  gate1160(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate1161(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate1162(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate2129(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate2130(.a(gate279inter0), .b(s_226), .O(gate279inter1));
  and2  gate2131(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate2132(.a(s_226), .O(gate279inter3));
  inv1  gate2133(.a(s_227), .O(gate279inter4));
  nand2 gate2134(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate2135(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate2136(.a(G651), .O(gate279inter7));
  inv1  gate2137(.a(G803), .O(gate279inter8));
  nand2 gate2138(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate2139(.a(s_227), .b(gate279inter3), .O(gate279inter10));
  nor2  gate2140(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate2141(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate2142(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );

  xor2  gate2213(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate2214(.a(gate281inter0), .b(s_238), .O(gate281inter1));
  and2  gate2215(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate2216(.a(s_238), .O(gate281inter3));
  inv1  gate2217(.a(s_239), .O(gate281inter4));
  nand2 gate2218(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate2219(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate2220(.a(G654), .O(gate281inter7));
  inv1  gate2221(.a(G806), .O(gate281inter8));
  nand2 gate2222(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate2223(.a(s_239), .b(gate281inter3), .O(gate281inter10));
  nor2  gate2224(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate2225(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate2226(.a(gate281inter12), .b(gate281inter1), .O(G826));

  xor2  gate1205(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate1206(.a(gate282inter0), .b(s_94), .O(gate282inter1));
  and2  gate1207(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate1208(.a(s_94), .O(gate282inter3));
  inv1  gate1209(.a(s_95), .O(gate282inter4));
  nand2 gate1210(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate1211(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate1212(.a(G782), .O(gate282inter7));
  inv1  gate1213(.a(G806), .O(gate282inter8));
  nand2 gate1214(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate1215(.a(s_95), .b(gate282inter3), .O(gate282inter10));
  nor2  gate1216(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate1217(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate1218(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate1345(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate1346(.a(gate286inter0), .b(s_114), .O(gate286inter1));
  and2  gate1347(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate1348(.a(s_114), .O(gate286inter3));
  inv1  gate1349(.a(s_115), .O(gate286inter4));
  nand2 gate1350(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate1351(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate1352(.a(G788), .O(gate286inter7));
  inv1  gate1353(.a(G812), .O(gate286inter8));
  nand2 gate1354(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate1355(.a(s_115), .b(gate286inter3), .O(gate286inter10));
  nor2  gate1356(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate1357(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate1358(.a(gate286inter12), .b(gate286inter1), .O(G831));

  xor2  gate1835(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate1836(.a(gate287inter0), .b(s_184), .O(gate287inter1));
  and2  gate1837(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate1838(.a(s_184), .O(gate287inter3));
  inv1  gate1839(.a(s_185), .O(gate287inter4));
  nand2 gate1840(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate1841(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate1842(.a(G663), .O(gate287inter7));
  inv1  gate1843(.a(G815), .O(gate287inter8));
  nand2 gate1844(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate1845(.a(s_185), .b(gate287inter3), .O(gate287inter10));
  nor2  gate1846(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate1847(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate1848(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate1527(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate1528(.a(gate290inter0), .b(s_140), .O(gate290inter1));
  and2  gate1529(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate1530(.a(s_140), .O(gate290inter3));
  inv1  gate1531(.a(s_141), .O(gate290inter4));
  nand2 gate1532(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate1533(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate1534(.a(G820), .O(gate290inter7));
  inv1  gate1535(.a(G821), .O(gate290inter8));
  nand2 gate1536(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate1537(.a(s_141), .b(gate290inter3), .O(gate290inter10));
  nor2  gate1538(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate1539(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate1540(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate2045(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate2046(.a(gate389inter0), .b(s_214), .O(gate389inter1));
  and2  gate2047(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate2048(.a(s_214), .O(gate389inter3));
  inv1  gate2049(.a(s_215), .O(gate389inter4));
  nand2 gate2050(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate2051(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate2052(.a(G3), .O(gate389inter7));
  inv1  gate2053(.a(G1042), .O(gate389inter8));
  nand2 gate2054(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate2055(.a(s_215), .b(gate389inter3), .O(gate389inter10));
  nor2  gate2056(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate2057(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate2058(.a(gate389inter12), .b(gate389inter1), .O(G1138));

  xor2  gate1597(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate1598(.a(gate390inter0), .b(s_150), .O(gate390inter1));
  and2  gate1599(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate1600(.a(s_150), .O(gate390inter3));
  inv1  gate1601(.a(s_151), .O(gate390inter4));
  nand2 gate1602(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate1603(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate1604(.a(G4), .O(gate390inter7));
  inv1  gate1605(.a(G1045), .O(gate390inter8));
  nand2 gate1606(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate1607(.a(s_151), .b(gate390inter3), .O(gate390inter10));
  nor2  gate1608(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate1609(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate1610(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate1667(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate1668(.a(gate393inter0), .b(s_160), .O(gate393inter1));
  and2  gate1669(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate1670(.a(s_160), .O(gate393inter3));
  inv1  gate1671(.a(s_161), .O(gate393inter4));
  nand2 gate1672(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate1673(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate1674(.a(G7), .O(gate393inter7));
  inv1  gate1675(.a(G1054), .O(gate393inter8));
  nand2 gate1676(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate1677(.a(s_161), .b(gate393inter3), .O(gate393inter10));
  nor2  gate1678(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate1679(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate1680(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate645(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate646(.a(gate403inter0), .b(s_14), .O(gate403inter1));
  and2  gate647(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate648(.a(s_14), .O(gate403inter3));
  inv1  gate649(.a(s_15), .O(gate403inter4));
  nand2 gate650(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate651(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate652(.a(G17), .O(gate403inter7));
  inv1  gate653(.a(G1084), .O(gate403inter8));
  nand2 gate654(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate655(.a(s_15), .b(gate403inter3), .O(gate403inter10));
  nor2  gate656(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate657(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate658(.a(gate403inter12), .b(gate403inter1), .O(G1180));
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate1401(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate1402(.a(gate410inter0), .b(s_122), .O(gate410inter1));
  and2  gate1403(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate1404(.a(s_122), .O(gate410inter3));
  inv1  gate1405(.a(s_123), .O(gate410inter4));
  nand2 gate1406(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate1407(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate1408(.a(G24), .O(gate410inter7));
  inv1  gate1409(.a(G1105), .O(gate410inter8));
  nand2 gate1410(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate1411(.a(s_123), .b(gate410inter3), .O(gate410inter10));
  nor2  gate1412(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate1413(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate1414(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate1233(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate1234(.a(gate413inter0), .b(s_98), .O(gate413inter1));
  and2  gate1235(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate1236(.a(s_98), .O(gate413inter3));
  inv1  gate1237(.a(s_99), .O(gate413inter4));
  nand2 gate1238(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1239(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1240(.a(G27), .O(gate413inter7));
  inv1  gate1241(.a(G1114), .O(gate413inter8));
  nand2 gate1242(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1243(.a(s_99), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1244(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1245(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1246(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate2353(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate2354(.a(gate415inter0), .b(s_258), .O(gate415inter1));
  and2  gate2355(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate2356(.a(s_258), .O(gate415inter3));
  inv1  gate2357(.a(s_259), .O(gate415inter4));
  nand2 gate2358(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate2359(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate2360(.a(G29), .O(gate415inter7));
  inv1  gate2361(.a(G1120), .O(gate415inter8));
  nand2 gate2362(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate2363(.a(s_259), .b(gate415inter3), .O(gate415inter10));
  nor2  gate2364(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate2365(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate2366(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );

  xor2  gate813(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate814(.a(gate418inter0), .b(s_38), .O(gate418inter1));
  and2  gate815(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate816(.a(s_38), .O(gate418inter3));
  inv1  gate817(.a(s_39), .O(gate418inter4));
  nand2 gate818(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate819(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate820(.a(G32), .O(gate418inter7));
  inv1  gate821(.a(G1129), .O(gate418inter8));
  nand2 gate822(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate823(.a(s_39), .b(gate418inter3), .O(gate418inter10));
  nor2  gate824(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate825(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate826(.a(gate418inter12), .b(gate418inter1), .O(G1225));

  xor2  gate2339(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate2340(.a(gate419inter0), .b(s_256), .O(gate419inter1));
  and2  gate2341(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate2342(.a(s_256), .O(gate419inter3));
  inv1  gate2343(.a(s_257), .O(gate419inter4));
  nand2 gate2344(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate2345(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate2346(.a(G1), .O(gate419inter7));
  inv1  gate2347(.a(G1132), .O(gate419inter8));
  nand2 gate2348(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate2349(.a(s_257), .b(gate419inter3), .O(gate419inter10));
  nor2  gate2350(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate2351(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate2352(.a(gate419inter12), .b(gate419inter1), .O(G1228));

  xor2  gate2003(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate2004(.a(gate420inter0), .b(s_208), .O(gate420inter1));
  and2  gate2005(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate2006(.a(s_208), .O(gate420inter3));
  inv1  gate2007(.a(s_209), .O(gate420inter4));
  nand2 gate2008(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate2009(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate2010(.a(G1036), .O(gate420inter7));
  inv1  gate2011(.a(G1132), .O(gate420inter8));
  nand2 gate2012(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate2013(.a(s_209), .b(gate420inter3), .O(gate420inter10));
  nor2  gate2014(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate2015(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate2016(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate1457(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate1458(.a(gate428inter0), .b(s_130), .O(gate428inter1));
  and2  gate1459(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate1460(.a(s_130), .O(gate428inter3));
  inv1  gate1461(.a(s_131), .O(gate428inter4));
  nand2 gate1462(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate1463(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate1464(.a(G1048), .O(gate428inter7));
  inv1  gate1465(.a(G1144), .O(gate428inter8));
  nand2 gate1466(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate1467(.a(s_131), .b(gate428inter3), .O(gate428inter10));
  nor2  gate1468(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate1469(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate1470(.a(gate428inter12), .b(gate428inter1), .O(G1237));

  xor2  gate1583(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate1584(.a(gate429inter0), .b(s_148), .O(gate429inter1));
  and2  gate1585(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate1586(.a(s_148), .O(gate429inter3));
  inv1  gate1587(.a(s_149), .O(gate429inter4));
  nand2 gate1588(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate1589(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate1590(.a(G6), .O(gate429inter7));
  inv1  gate1591(.a(G1147), .O(gate429inter8));
  nand2 gate1592(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate1593(.a(s_149), .b(gate429inter3), .O(gate429inter10));
  nor2  gate1594(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate1595(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate1596(.a(gate429inter12), .b(gate429inter1), .O(G1238));
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate1779(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate1780(.a(gate437inter0), .b(s_176), .O(gate437inter1));
  and2  gate1781(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate1782(.a(s_176), .O(gate437inter3));
  inv1  gate1783(.a(s_177), .O(gate437inter4));
  nand2 gate1784(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate1785(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate1786(.a(G10), .O(gate437inter7));
  inv1  gate1787(.a(G1159), .O(gate437inter8));
  nand2 gate1788(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate1789(.a(s_177), .b(gate437inter3), .O(gate437inter10));
  nor2  gate1790(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate1791(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate1792(.a(gate437inter12), .b(gate437inter1), .O(G1246));

  xor2  gate1513(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate1514(.a(gate438inter0), .b(s_138), .O(gate438inter1));
  and2  gate1515(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate1516(.a(s_138), .O(gate438inter3));
  inv1  gate1517(.a(s_139), .O(gate438inter4));
  nand2 gate1518(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate1519(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate1520(.a(G1063), .O(gate438inter7));
  inv1  gate1521(.a(G1159), .O(gate438inter8));
  nand2 gate1522(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate1523(.a(s_139), .b(gate438inter3), .O(gate438inter10));
  nor2  gate1524(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate1525(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate1526(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate2227(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate2228(.a(gate441inter0), .b(s_240), .O(gate441inter1));
  and2  gate2229(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate2230(.a(s_240), .O(gate441inter3));
  inv1  gate2231(.a(s_241), .O(gate441inter4));
  nand2 gate2232(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate2233(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate2234(.a(G12), .O(gate441inter7));
  inv1  gate2235(.a(G1165), .O(gate441inter8));
  nand2 gate2236(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate2237(.a(s_241), .b(gate441inter3), .O(gate441inter10));
  nor2  gate2238(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate2239(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate2240(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate1737(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate1738(.a(gate443inter0), .b(s_170), .O(gate443inter1));
  and2  gate1739(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate1740(.a(s_170), .O(gate443inter3));
  inv1  gate1741(.a(s_171), .O(gate443inter4));
  nand2 gate1742(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate1743(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate1744(.a(G13), .O(gate443inter7));
  inv1  gate1745(.a(G1168), .O(gate443inter8));
  nand2 gate1746(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate1747(.a(s_171), .b(gate443inter3), .O(gate443inter10));
  nor2  gate1748(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate1749(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate1750(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate1093(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate1094(.a(gate445inter0), .b(s_78), .O(gate445inter1));
  and2  gate1095(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate1096(.a(s_78), .O(gate445inter3));
  inv1  gate1097(.a(s_79), .O(gate445inter4));
  nand2 gate1098(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate1099(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate1100(.a(G14), .O(gate445inter7));
  inv1  gate1101(.a(G1171), .O(gate445inter8));
  nand2 gate1102(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate1103(.a(s_79), .b(gate445inter3), .O(gate445inter10));
  nor2  gate1104(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate1105(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate1106(.a(gate445inter12), .b(gate445inter1), .O(G1254));

  xor2  gate1905(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate1906(.a(gate446inter0), .b(s_194), .O(gate446inter1));
  and2  gate1907(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate1908(.a(s_194), .O(gate446inter3));
  inv1  gate1909(.a(s_195), .O(gate446inter4));
  nand2 gate1910(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate1911(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate1912(.a(G1075), .O(gate446inter7));
  inv1  gate1913(.a(G1171), .O(gate446inter8));
  nand2 gate1914(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate1915(.a(s_195), .b(gate446inter3), .O(gate446inter10));
  nor2  gate1916(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate1917(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate1918(.a(gate446inter12), .b(gate446inter1), .O(G1255));
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );

  xor2  gate1009(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate1010(.a(gate450inter0), .b(s_66), .O(gate450inter1));
  and2  gate1011(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate1012(.a(s_66), .O(gate450inter3));
  inv1  gate1013(.a(s_67), .O(gate450inter4));
  nand2 gate1014(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate1015(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate1016(.a(G1081), .O(gate450inter7));
  inv1  gate1017(.a(G1177), .O(gate450inter8));
  nand2 gate1018(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate1019(.a(s_67), .b(gate450inter3), .O(gate450inter10));
  nor2  gate1020(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate1021(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate1022(.a(gate450inter12), .b(gate450inter1), .O(G1259));
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate1471(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate1472(.a(gate461inter0), .b(s_132), .O(gate461inter1));
  and2  gate1473(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate1474(.a(s_132), .O(gate461inter3));
  inv1  gate1475(.a(s_133), .O(gate461inter4));
  nand2 gate1476(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate1477(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate1478(.a(G22), .O(gate461inter7));
  inv1  gate1479(.a(G1195), .O(gate461inter8));
  nand2 gate1480(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate1481(.a(s_133), .b(gate461inter3), .O(gate461inter10));
  nor2  gate1482(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate1483(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate1484(.a(gate461inter12), .b(gate461inter1), .O(G1270));
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );

  xor2  gate2437(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate2438(.a(gate468inter0), .b(s_270), .O(gate468inter1));
  and2  gate2439(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate2440(.a(s_270), .O(gate468inter3));
  inv1  gate2441(.a(s_271), .O(gate468inter4));
  nand2 gate2442(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate2443(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate2444(.a(G1108), .O(gate468inter7));
  inv1  gate2445(.a(G1204), .O(gate468inter8));
  nand2 gate2446(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate2447(.a(s_271), .b(gate468inter3), .O(gate468inter10));
  nor2  gate2448(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate2449(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate2450(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );

  xor2  gate981(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate982(.a(gate470inter0), .b(s_62), .O(gate470inter1));
  and2  gate983(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate984(.a(s_62), .O(gate470inter3));
  inv1  gate985(.a(s_63), .O(gate470inter4));
  nand2 gate986(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate987(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate988(.a(G1111), .O(gate470inter7));
  inv1  gate989(.a(G1207), .O(gate470inter8));
  nand2 gate990(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate991(.a(s_63), .b(gate470inter3), .O(gate470inter10));
  nor2  gate992(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate993(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate994(.a(gate470inter12), .b(gate470inter1), .O(G1279));
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate1723(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate1724(.a(gate472inter0), .b(s_168), .O(gate472inter1));
  and2  gate1725(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate1726(.a(s_168), .O(gate472inter3));
  inv1  gate1727(.a(s_169), .O(gate472inter4));
  nand2 gate1728(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate1729(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate1730(.a(G1114), .O(gate472inter7));
  inv1  gate1731(.a(G1210), .O(gate472inter8));
  nand2 gate1732(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate1733(.a(s_169), .b(gate472inter3), .O(gate472inter10));
  nor2  gate1734(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate1735(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate1736(.a(gate472inter12), .b(gate472inter1), .O(G1281));

  xor2  gate2073(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate2074(.a(gate473inter0), .b(s_218), .O(gate473inter1));
  and2  gate2075(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate2076(.a(s_218), .O(gate473inter3));
  inv1  gate2077(.a(s_219), .O(gate473inter4));
  nand2 gate2078(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate2079(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate2080(.a(G28), .O(gate473inter7));
  inv1  gate2081(.a(G1213), .O(gate473inter8));
  nand2 gate2082(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate2083(.a(s_219), .b(gate473inter3), .O(gate473inter10));
  nor2  gate2084(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate2085(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate2086(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate2367(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate2368(.a(gate480inter0), .b(s_260), .O(gate480inter1));
  and2  gate2369(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate2370(.a(s_260), .O(gate480inter3));
  inv1  gate2371(.a(s_261), .O(gate480inter4));
  nand2 gate2372(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate2373(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate2374(.a(G1126), .O(gate480inter7));
  inv1  gate2375(.a(G1222), .O(gate480inter8));
  nand2 gate2376(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate2377(.a(s_261), .b(gate480inter3), .O(gate480inter10));
  nor2  gate2378(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate2379(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate2380(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate1709(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate1710(.a(gate485inter0), .b(s_166), .O(gate485inter1));
  and2  gate1711(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate1712(.a(s_166), .O(gate485inter3));
  inv1  gate1713(.a(s_167), .O(gate485inter4));
  nand2 gate1714(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate1715(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate1716(.a(G1232), .O(gate485inter7));
  inv1  gate1717(.a(G1233), .O(gate485inter8));
  nand2 gate1718(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate1719(.a(s_167), .b(gate485inter3), .O(gate485inter10));
  nor2  gate1720(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate1721(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate1722(.a(gate485inter12), .b(gate485inter1), .O(G1294));

  xor2  gate1415(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate1416(.a(gate486inter0), .b(s_124), .O(gate486inter1));
  and2  gate1417(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate1418(.a(s_124), .O(gate486inter3));
  inv1  gate1419(.a(s_125), .O(gate486inter4));
  nand2 gate1420(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate1421(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate1422(.a(G1234), .O(gate486inter7));
  inv1  gate1423(.a(G1235), .O(gate486inter8));
  nand2 gate1424(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate1425(.a(s_125), .b(gate486inter3), .O(gate486inter10));
  nor2  gate1426(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate1427(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate1428(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate1639(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate1640(.a(gate490inter0), .b(s_156), .O(gate490inter1));
  and2  gate1641(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate1642(.a(s_156), .O(gate490inter3));
  inv1  gate1643(.a(s_157), .O(gate490inter4));
  nand2 gate1644(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate1645(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate1646(.a(G1242), .O(gate490inter7));
  inv1  gate1647(.a(G1243), .O(gate490inter8));
  nand2 gate1648(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate1649(.a(s_157), .b(gate490inter3), .O(gate490inter10));
  nor2  gate1650(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate1651(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate1652(.a(gate490inter12), .b(gate490inter1), .O(G1299));

  xor2  gate2283(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate2284(.a(gate491inter0), .b(s_248), .O(gate491inter1));
  and2  gate2285(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate2286(.a(s_248), .O(gate491inter3));
  inv1  gate2287(.a(s_249), .O(gate491inter4));
  nand2 gate2288(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate2289(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate2290(.a(G1244), .O(gate491inter7));
  inv1  gate2291(.a(G1245), .O(gate491inter8));
  nand2 gate2292(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate2293(.a(s_249), .b(gate491inter3), .O(gate491inter10));
  nor2  gate2294(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate2295(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate2296(.a(gate491inter12), .b(gate491inter1), .O(G1300));

  xor2  gate1625(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate1626(.a(gate492inter0), .b(s_154), .O(gate492inter1));
  and2  gate1627(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate1628(.a(s_154), .O(gate492inter3));
  inv1  gate1629(.a(s_155), .O(gate492inter4));
  nand2 gate1630(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate1631(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate1632(.a(G1246), .O(gate492inter7));
  inv1  gate1633(.a(G1247), .O(gate492inter8));
  nand2 gate1634(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate1635(.a(s_155), .b(gate492inter3), .O(gate492inter10));
  nor2  gate1636(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate1637(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate1638(.a(gate492inter12), .b(gate492inter1), .O(G1301));

  xor2  gate2087(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate2088(.a(gate493inter0), .b(s_220), .O(gate493inter1));
  and2  gate2089(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate2090(.a(s_220), .O(gate493inter3));
  inv1  gate2091(.a(s_221), .O(gate493inter4));
  nand2 gate2092(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate2093(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate2094(.a(G1248), .O(gate493inter7));
  inv1  gate2095(.a(G1249), .O(gate493inter8));
  nand2 gate2096(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate2097(.a(s_221), .b(gate493inter3), .O(gate493inter10));
  nor2  gate2098(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate2099(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate2100(.a(gate493inter12), .b(gate493inter1), .O(G1302));
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );

  xor2  gate1317(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate1318(.a(gate498inter0), .b(s_110), .O(gate498inter1));
  and2  gate1319(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate1320(.a(s_110), .O(gate498inter3));
  inv1  gate1321(.a(s_111), .O(gate498inter4));
  nand2 gate1322(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate1323(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate1324(.a(G1258), .O(gate498inter7));
  inv1  gate1325(.a(G1259), .O(gate498inter8));
  nand2 gate1326(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate1327(.a(s_111), .b(gate498inter3), .O(gate498inter10));
  nor2  gate1328(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate1329(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate1330(.a(gate498inter12), .b(gate498inter1), .O(G1307));
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate2269(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate2270(.a(gate500inter0), .b(s_246), .O(gate500inter1));
  and2  gate2271(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate2272(.a(s_246), .O(gate500inter3));
  inv1  gate2273(.a(s_247), .O(gate500inter4));
  nand2 gate2274(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate2275(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate2276(.a(G1262), .O(gate500inter7));
  inv1  gate2277(.a(G1263), .O(gate500inter8));
  nand2 gate2278(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate2279(.a(s_247), .b(gate500inter3), .O(gate500inter10));
  nor2  gate2280(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate2281(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate2282(.a(gate500inter12), .b(gate500inter1), .O(G1309));

  xor2  gate897(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate898(.a(gate501inter0), .b(s_50), .O(gate501inter1));
  and2  gate899(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate900(.a(s_50), .O(gate501inter3));
  inv1  gate901(.a(s_51), .O(gate501inter4));
  nand2 gate902(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate903(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate904(.a(G1264), .O(gate501inter7));
  inv1  gate905(.a(G1265), .O(gate501inter8));
  nand2 gate906(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate907(.a(s_51), .b(gate501inter3), .O(gate501inter10));
  nor2  gate908(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate909(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate910(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );

  xor2  gate2297(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate2298(.a(gate505inter0), .b(s_250), .O(gate505inter1));
  and2  gate2299(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate2300(.a(s_250), .O(gate505inter3));
  inv1  gate2301(.a(s_251), .O(gate505inter4));
  nand2 gate2302(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate2303(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate2304(.a(G1272), .O(gate505inter7));
  inv1  gate2305(.a(G1273), .O(gate505inter8));
  nand2 gate2306(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate2307(.a(s_251), .b(gate505inter3), .O(gate505inter10));
  nor2  gate2308(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate2309(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate2310(.a(gate505inter12), .b(gate505inter1), .O(G1314));
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule