module c499 (N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
             N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
             N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
             N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
             N137,N724,N725,N726,N727,N728,N729,N730,N731,N732,
             N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,
             N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,
             N753,N754,N755);
input N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
      N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
      N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
      N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
      N137;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81;
output N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,
       N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
       N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
       N754,N755;
wire N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
     N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
     N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,
     N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,
     N290,N293,N296,N299,N302,N305,N308,N311,N314,N315,
     N316,N317,N318,N319,N320,N321,N338,N339,N340,N341,
     N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,
     N352,N353,N354,N367,N380,N393,N406,N419,N432,N445,
     N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
     N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,
     N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,
     N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,
     N594,N595,N596,N597,N598,N599,N600,N601,N602,N607,
     N620,N625,N630,N635,N640,N645,N650,N655,N692,N693,
     N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,
     N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,
     N714,N715,N716,N717,N718,N719,N720,N721,N722,N723, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate2inter0, gate2inter1, gate2inter2, gate2inter3, gate2inter4, gate2inter5, gate2inter6, gate2inter7, gate2inter8, gate2inter9, gate2inter10, gate2inter11, gate2inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate8inter0, gate8inter1, gate8inter2, gate8inter3, gate8inter4, gate8inter5, gate8inter6, gate8inter7, gate8inter8, gate8inter9, gate8inter10, gate8inter11, gate8inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12;


xor2 gate1( .a(N1), .b(N5), .O(N250) );

  xor2  gate441(.a(N13), .b(N9), .O(gate2inter0));
  nand2 gate442(.a(gate2inter0), .b(s_34), .O(gate2inter1));
  and2  gate443(.a(N13), .b(N9), .O(gate2inter2));
  inv1  gate444(.a(s_34), .O(gate2inter3));
  inv1  gate445(.a(s_35), .O(gate2inter4));
  nand2 gate446(.a(gate2inter4), .b(gate2inter3), .O(gate2inter5));
  nor2  gate447(.a(gate2inter5), .b(gate2inter2), .O(gate2inter6));
  inv1  gate448(.a(N9), .O(gate2inter7));
  inv1  gate449(.a(N13), .O(gate2inter8));
  nand2 gate450(.a(gate2inter8), .b(gate2inter7), .O(gate2inter9));
  nand2 gate451(.a(s_35), .b(gate2inter3), .O(gate2inter10));
  nor2  gate452(.a(gate2inter10), .b(gate2inter9), .O(gate2inter11));
  nor2  gate453(.a(gate2inter11), .b(gate2inter6), .O(gate2inter12));
  nand2 gate454(.a(gate2inter12), .b(gate2inter1), .O(N251));
xor2 gate3( .a(N17), .b(N21), .O(N252) );
xor2 gate4( .a(N25), .b(N29), .O(N253) );
xor2 gate5( .a(N33), .b(N37), .O(N254) );
xor2 gate6( .a(N41), .b(N45), .O(N255) );
xor2 gate7( .a(N49), .b(N53), .O(N256) );

  xor2  gate735(.a(N61), .b(N57), .O(gate8inter0));
  nand2 gate736(.a(gate8inter0), .b(s_76), .O(gate8inter1));
  and2  gate737(.a(N61), .b(N57), .O(gate8inter2));
  inv1  gate738(.a(s_76), .O(gate8inter3));
  inv1  gate739(.a(s_77), .O(gate8inter4));
  nand2 gate740(.a(gate8inter4), .b(gate8inter3), .O(gate8inter5));
  nor2  gate741(.a(gate8inter5), .b(gate8inter2), .O(gate8inter6));
  inv1  gate742(.a(N57), .O(gate8inter7));
  inv1  gate743(.a(N61), .O(gate8inter8));
  nand2 gate744(.a(gate8inter8), .b(gate8inter7), .O(gate8inter9));
  nand2 gate745(.a(s_77), .b(gate8inter3), .O(gate8inter10));
  nor2  gate746(.a(gate8inter10), .b(gate8inter9), .O(gate8inter11));
  nor2  gate747(.a(gate8inter11), .b(gate8inter6), .O(gate8inter12));
  nand2 gate748(.a(gate8inter12), .b(gate8inter1), .O(N257));

  xor2  gate399(.a(N69), .b(N65), .O(gate9inter0));
  nand2 gate400(.a(gate9inter0), .b(s_28), .O(gate9inter1));
  and2  gate401(.a(N69), .b(N65), .O(gate9inter2));
  inv1  gate402(.a(s_28), .O(gate9inter3));
  inv1  gate403(.a(s_29), .O(gate9inter4));
  nand2 gate404(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate405(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate406(.a(N65), .O(gate9inter7));
  inv1  gate407(.a(N69), .O(gate9inter8));
  nand2 gate408(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate409(.a(s_29), .b(gate9inter3), .O(gate9inter10));
  nor2  gate410(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate411(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate412(.a(gate9inter12), .b(gate9inter1), .O(N258));
xor2 gate10( .a(N73), .b(N77), .O(N259) );
xor2 gate11( .a(N81), .b(N85), .O(N260) );
xor2 gate12( .a(N89), .b(N93), .O(N261) );
xor2 gate13( .a(N97), .b(N101), .O(N262) );
xor2 gate14( .a(N105), .b(N109), .O(N263) );

  xor2  gate651(.a(N117), .b(N113), .O(gate15inter0));
  nand2 gate652(.a(gate15inter0), .b(s_64), .O(gate15inter1));
  and2  gate653(.a(N117), .b(N113), .O(gate15inter2));
  inv1  gate654(.a(s_64), .O(gate15inter3));
  inv1  gate655(.a(s_65), .O(gate15inter4));
  nand2 gate656(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate657(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate658(.a(N113), .O(gate15inter7));
  inv1  gate659(.a(N117), .O(gate15inter8));
  nand2 gate660(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate661(.a(s_65), .b(gate15inter3), .O(gate15inter10));
  nor2  gate662(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate663(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate664(.a(gate15inter12), .b(gate15inter1), .O(N264));
xor2 gate16( .a(N121), .b(N125), .O(N265) );
and2 gate17( .a(N129), .b(N137), .O(N266) );
and2 gate18( .a(N130), .b(N137), .O(N267) );
and2 gate19( .a(N131), .b(N137), .O(N268) );
and2 gate20( .a(N132), .b(N137), .O(N269) );
and2 gate21( .a(N133), .b(N137), .O(N270) );
and2 gate22( .a(N134), .b(N137), .O(N271) );
and2 gate23( .a(N135), .b(N137), .O(N272) );
and2 gate24( .a(N136), .b(N137), .O(N273) );
xor2 gate25( .a(N1), .b(N17), .O(N274) );
xor2 gate26( .a(N33), .b(N49), .O(N275) );
xor2 gate27( .a(N5), .b(N21), .O(N276) );
xor2 gate28( .a(N37), .b(N53), .O(N277) );

  xor2  gate413(.a(N25), .b(N9), .O(gate29inter0));
  nand2 gate414(.a(gate29inter0), .b(s_30), .O(gate29inter1));
  and2  gate415(.a(N25), .b(N9), .O(gate29inter2));
  inv1  gate416(.a(s_30), .O(gate29inter3));
  inv1  gate417(.a(s_31), .O(gate29inter4));
  nand2 gate418(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate419(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate420(.a(N9), .O(gate29inter7));
  inv1  gate421(.a(N25), .O(gate29inter8));
  nand2 gate422(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate423(.a(s_31), .b(gate29inter3), .O(gate29inter10));
  nor2  gate424(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate425(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate426(.a(gate29inter12), .b(gate29inter1), .O(N278));

  xor2  gate553(.a(N57), .b(N41), .O(gate30inter0));
  nand2 gate554(.a(gate30inter0), .b(s_50), .O(gate30inter1));
  and2  gate555(.a(N57), .b(N41), .O(gate30inter2));
  inv1  gate556(.a(s_50), .O(gate30inter3));
  inv1  gate557(.a(s_51), .O(gate30inter4));
  nand2 gate558(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate559(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate560(.a(N41), .O(gate30inter7));
  inv1  gate561(.a(N57), .O(gate30inter8));
  nand2 gate562(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate563(.a(s_51), .b(gate30inter3), .O(gate30inter10));
  nor2  gate564(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate565(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate566(.a(gate30inter12), .b(gate30inter1), .O(N279));

  xor2  gate511(.a(N29), .b(N13), .O(gate31inter0));
  nand2 gate512(.a(gate31inter0), .b(s_44), .O(gate31inter1));
  and2  gate513(.a(N29), .b(N13), .O(gate31inter2));
  inv1  gate514(.a(s_44), .O(gate31inter3));
  inv1  gate515(.a(s_45), .O(gate31inter4));
  nand2 gate516(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate517(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate518(.a(N13), .O(gate31inter7));
  inv1  gate519(.a(N29), .O(gate31inter8));
  nand2 gate520(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate521(.a(s_45), .b(gate31inter3), .O(gate31inter10));
  nor2  gate522(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate523(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate524(.a(gate31inter12), .b(gate31inter1), .O(N280));
xor2 gate32( .a(N45), .b(N61), .O(N281) );
xor2 gate33( .a(N65), .b(N81), .O(N282) );

  xor2  gate455(.a(N113), .b(N97), .O(gate34inter0));
  nand2 gate456(.a(gate34inter0), .b(s_36), .O(gate34inter1));
  and2  gate457(.a(N113), .b(N97), .O(gate34inter2));
  inv1  gate458(.a(s_36), .O(gate34inter3));
  inv1  gate459(.a(s_37), .O(gate34inter4));
  nand2 gate460(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate461(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate462(.a(N97), .O(gate34inter7));
  inv1  gate463(.a(N113), .O(gate34inter8));
  nand2 gate464(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate465(.a(s_37), .b(gate34inter3), .O(gate34inter10));
  nor2  gate466(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate467(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate468(.a(gate34inter12), .b(gate34inter1), .O(N283));
xor2 gate35( .a(N69), .b(N85), .O(N284) );

  xor2  gate637(.a(N117), .b(N101), .O(gate36inter0));
  nand2 gate638(.a(gate36inter0), .b(s_62), .O(gate36inter1));
  and2  gate639(.a(N117), .b(N101), .O(gate36inter2));
  inv1  gate640(.a(s_62), .O(gate36inter3));
  inv1  gate641(.a(s_63), .O(gate36inter4));
  nand2 gate642(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate643(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate644(.a(N101), .O(gate36inter7));
  inv1  gate645(.a(N117), .O(gate36inter8));
  nand2 gate646(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate647(.a(s_63), .b(gate36inter3), .O(gate36inter10));
  nor2  gate648(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate649(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate650(.a(gate36inter12), .b(gate36inter1), .O(N285));

  xor2  gate525(.a(N89), .b(N73), .O(gate37inter0));
  nand2 gate526(.a(gate37inter0), .b(s_46), .O(gate37inter1));
  and2  gate527(.a(N89), .b(N73), .O(gate37inter2));
  inv1  gate528(.a(s_46), .O(gate37inter3));
  inv1  gate529(.a(s_47), .O(gate37inter4));
  nand2 gate530(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate531(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate532(.a(N73), .O(gate37inter7));
  inv1  gate533(.a(N89), .O(gate37inter8));
  nand2 gate534(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate535(.a(s_47), .b(gate37inter3), .O(gate37inter10));
  nor2  gate536(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate537(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate538(.a(gate37inter12), .b(gate37inter1), .O(N286));
xor2 gate38( .a(N105), .b(N121), .O(N287) );
xor2 gate39( .a(N77), .b(N93), .O(N288) );
xor2 gate40( .a(N109), .b(N125), .O(N289) );

  xor2  gate707(.a(N251), .b(N250), .O(gate41inter0));
  nand2 gate708(.a(gate41inter0), .b(s_72), .O(gate41inter1));
  and2  gate709(.a(N251), .b(N250), .O(gate41inter2));
  inv1  gate710(.a(s_72), .O(gate41inter3));
  inv1  gate711(.a(s_73), .O(gate41inter4));
  nand2 gate712(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate713(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate714(.a(N250), .O(gate41inter7));
  inv1  gate715(.a(N251), .O(gate41inter8));
  nand2 gate716(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate717(.a(s_73), .b(gate41inter3), .O(gate41inter10));
  nor2  gate718(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate719(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate720(.a(gate41inter12), .b(gate41inter1), .O(N290));

  xor2  gate595(.a(N253), .b(N252), .O(gate42inter0));
  nand2 gate596(.a(gate42inter0), .b(s_56), .O(gate42inter1));
  and2  gate597(.a(N253), .b(N252), .O(gate42inter2));
  inv1  gate598(.a(s_56), .O(gate42inter3));
  inv1  gate599(.a(s_57), .O(gate42inter4));
  nand2 gate600(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate601(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate602(.a(N252), .O(gate42inter7));
  inv1  gate603(.a(N253), .O(gate42inter8));
  nand2 gate604(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate605(.a(s_57), .b(gate42inter3), .O(gate42inter10));
  nor2  gate606(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate607(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate608(.a(gate42inter12), .b(gate42inter1), .O(N293));

  xor2  gate357(.a(N255), .b(N254), .O(gate43inter0));
  nand2 gate358(.a(gate43inter0), .b(s_22), .O(gate43inter1));
  and2  gate359(.a(N255), .b(N254), .O(gate43inter2));
  inv1  gate360(.a(s_22), .O(gate43inter3));
  inv1  gate361(.a(s_23), .O(gate43inter4));
  nand2 gate362(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate363(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate364(.a(N254), .O(gate43inter7));
  inv1  gate365(.a(N255), .O(gate43inter8));
  nand2 gate366(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate367(.a(s_23), .b(gate43inter3), .O(gate43inter10));
  nor2  gate368(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate369(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate370(.a(gate43inter12), .b(gate43inter1), .O(N296));
xor2 gate44( .a(N256), .b(N257), .O(N299) );
xor2 gate45( .a(N258), .b(N259), .O(N302) );
xor2 gate46( .a(N260), .b(N261), .O(N305) );

  xor2  gate287(.a(N263), .b(N262), .O(gate47inter0));
  nand2 gate288(.a(gate47inter0), .b(s_12), .O(gate47inter1));
  and2  gate289(.a(N263), .b(N262), .O(gate47inter2));
  inv1  gate290(.a(s_12), .O(gate47inter3));
  inv1  gate291(.a(s_13), .O(gate47inter4));
  nand2 gate292(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate293(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate294(.a(N262), .O(gate47inter7));
  inv1  gate295(.a(N263), .O(gate47inter8));
  nand2 gate296(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate297(.a(s_13), .b(gate47inter3), .O(gate47inter10));
  nor2  gate298(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate299(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate300(.a(gate47inter12), .b(gate47inter1), .O(N308));
xor2 gate48( .a(N264), .b(N265), .O(N311) );
xor2 gate49( .a(N274), .b(N275), .O(N314) );
xor2 gate50( .a(N276), .b(N277), .O(N315) );

  xor2  gate469(.a(N279), .b(N278), .O(gate51inter0));
  nand2 gate470(.a(gate51inter0), .b(s_38), .O(gate51inter1));
  and2  gate471(.a(N279), .b(N278), .O(gate51inter2));
  inv1  gate472(.a(s_38), .O(gate51inter3));
  inv1  gate473(.a(s_39), .O(gate51inter4));
  nand2 gate474(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate475(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate476(.a(N278), .O(gate51inter7));
  inv1  gate477(.a(N279), .O(gate51inter8));
  nand2 gate478(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate479(.a(s_39), .b(gate51inter3), .O(gate51inter10));
  nor2  gate480(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate481(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate482(.a(gate51inter12), .b(gate51inter1), .O(N316));
xor2 gate52( .a(N280), .b(N281), .O(N317) );
xor2 gate53( .a(N282), .b(N283), .O(N318) );

  xor2  gate567(.a(N285), .b(N284), .O(gate54inter0));
  nand2 gate568(.a(gate54inter0), .b(s_52), .O(gate54inter1));
  and2  gate569(.a(N285), .b(N284), .O(gate54inter2));
  inv1  gate570(.a(s_52), .O(gate54inter3));
  inv1  gate571(.a(s_53), .O(gate54inter4));
  nand2 gate572(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate573(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate574(.a(N284), .O(gate54inter7));
  inv1  gate575(.a(N285), .O(gate54inter8));
  nand2 gate576(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate577(.a(s_53), .b(gate54inter3), .O(gate54inter10));
  nor2  gate578(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate579(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate580(.a(gate54inter12), .b(gate54inter1), .O(N319));
xor2 gate55( .a(N286), .b(N287), .O(N320) );
xor2 gate56( .a(N288), .b(N289), .O(N321) );
xor2 gate57( .a(N290), .b(N293), .O(N338) );
xor2 gate58( .a(N296), .b(N299), .O(N339) );

  xor2  gate245(.a(N296), .b(N290), .O(gate59inter0));
  nand2 gate246(.a(gate59inter0), .b(s_6), .O(gate59inter1));
  and2  gate247(.a(N296), .b(N290), .O(gate59inter2));
  inv1  gate248(.a(s_6), .O(gate59inter3));
  inv1  gate249(.a(s_7), .O(gate59inter4));
  nand2 gate250(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate251(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate252(.a(N290), .O(gate59inter7));
  inv1  gate253(.a(N296), .O(gate59inter8));
  nand2 gate254(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate255(.a(s_7), .b(gate59inter3), .O(gate59inter10));
  nor2  gate256(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate257(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate258(.a(gate59inter12), .b(gate59inter1), .O(N340));

  xor2  gate343(.a(N299), .b(N293), .O(gate60inter0));
  nand2 gate344(.a(gate60inter0), .b(s_20), .O(gate60inter1));
  and2  gate345(.a(N299), .b(N293), .O(gate60inter2));
  inv1  gate346(.a(s_20), .O(gate60inter3));
  inv1  gate347(.a(s_21), .O(gate60inter4));
  nand2 gate348(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate349(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate350(.a(N293), .O(gate60inter7));
  inv1  gate351(.a(N299), .O(gate60inter8));
  nand2 gate352(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate353(.a(s_21), .b(gate60inter3), .O(gate60inter10));
  nor2  gate354(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate355(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate356(.a(gate60inter12), .b(gate60inter1), .O(N341));
xor2 gate61( .a(N302), .b(N305), .O(N342) );

  xor2  gate609(.a(N311), .b(N308), .O(gate62inter0));
  nand2 gate610(.a(gate62inter0), .b(s_58), .O(gate62inter1));
  and2  gate611(.a(N311), .b(N308), .O(gate62inter2));
  inv1  gate612(.a(s_58), .O(gate62inter3));
  inv1  gate613(.a(s_59), .O(gate62inter4));
  nand2 gate614(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate615(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate616(.a(N308), .O(gate62inter7));
  inv1  gate617(.a(N311), .O(gate62inter8));
  nand2 gate618(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate619(.a(s_59), .b(gate62inter3), .O(gate62inter10));
  nor2  gate620(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate621(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate622(.a(gate62inter12), .b(gate62inter1), .O(N343));
xor2 gate63( .a(N302), .b(N308), .O(N344) );
xor2 gate64( .a(N305), .b(N311), .O(N345) );

  xor2  gate217(.a(N342), .b(N266), .O(gate65inter0));
  nand2 gate218(.a(gate65inter0), .b(s_2), .O(gate65inter1));
  and2  gate219(.a(N342), .b(N266), .O(gate65inter2));
  inv1  gate220(.a(s_2), .O(gate65inter3));
  inv1  gate221(.a(s_3), .O(gate65inter4));
  nand2 gate222(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate223(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate224(.a(N266), .O(gate65inter7));
  inv1  gate225(.a(N342), .O(gate65inter8));
  nand2 gate226(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate227(.a(s_3), .b(gate65inter3), .O(gate65inter10));
  nor2  gate228(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate229(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate230(.a(gate65inter12), .b(gate65inter1), .O(N346));
xor2 gate66( .a(N267), .b(N343), .O(N347) );
xor2 gate67( .a(N268), .b(N344), .O(N348) );
xor2 gate68( .a(N269), .b(N345), .O(N349) );

  xor2  gate329(.a(N338), .b(N270), .O(gate69inter0));
  nand2 gate330(.a(gate69inter0), .b(s_18), .O(gate69inter1));
  and2  gate331(.a(N338), .b(N270), .O(gate69inter2));
  inv1  gate332(.a(s_18), .O(gate69inter3));
  inv1  gate333(.a(s_19), .O(gate69inter4));
  nand2 gate334(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate335(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate336(.a(N270), .O(gate69inter7));
  inv1  gate337(.a(N338), .O(gate69inter8));
  nand2 gate338(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate339(.a(s_19), .b(gate69inter3), .O(gate69inter10));
  nor2  gate340(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate341(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate342(.a(gate69inter12), .b(gate69inter1), .O(N350));

  xor2  gate679(.a(N339), .b(N271), .O(gate70inter0));
  nand2 gate680(.a(gate70inter0), .b(s_68), .O(gate70inter1));
  and2  gate681(.a(N339), .b(N271), .O(gate70inter2));
  inv1  gate682(.a(s_68), .O(gate70inter3));
  inv1  gate683(.a(s_69), .O(gate70inter4));
  nand2 gate684(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate685(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate686(.a(N271), .O(gate70inter7));
  inv1  gate687(.a(N339), .O(gate70inter8));
  nand2 gate688(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate689(.a(s_69), .b(gate70inter3), .O(gate70inter10));
  nor2  gate690(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate691(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate692(.a(gate70inter12), .b(gate70inter1), .O(N351));
xor2 gate71( .a(N272), .b(N340), .O(N352) );
xor2 gate72( .a(N273), .b(N341), .O(N353) );
xor2 gate73( .a(N314), .b(N346), .O(N354) );

  xor2  gate749(.a(N347), .b(N315), .O(gate74inter0));
  nand2 gate750(.a(gate74inter0), .b(s_78), .O(gate74inter1));
  and2  gate751(.a(N347), .b(N315), .O(gate74inter2));
  inv1  gate752(.a(s_78), .O(gate74inter3));
  inv1  gate753(.a(s_79), .O(gate74inter4));
  nand2 gate754(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate755(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate756(.a(N315), .O(gate74inter7));
  inv1  gate757(.a(N347), .O(gate74inter8));
  nand2 gate758(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate759(.a(s_79), .b(gate74inter3), .O(gate74inter10));
  nor2  gate760(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate761(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate762(.a(gate74inter12), .b(gate74inter1), .O(N367));
xor2 gate75( .a(N316), .b(N348), .O(N380) );
xor2 gate76( .a(N317), .b(N349), .O(N393) );

  xor2  gate371(.a(N350), .b(N318), .O(gate77inter0));
  nand2 gate372(.a(gate77inter0), .b(s_24), .O(gate77inter1));
  and2  gate373(.a(N350), .b(N318), .O(gate77inter2));
  inv1  gate374(.a(s_24), .O(gate77inter3));
  inv1  gate375(.a(s_25), .O(gate77inter4));
  nand2 gate376(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate377(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate378(.a(N318), .O(gate77inter7));
  inv1  gate379(.a(N350), .O(gate77inter8));
  nand2 gate380(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate381(.a(s_25), .b(gate77inter3), .O(gate77inter10));
  nor2  gate382(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate383(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate384(.a(gate77inter12), .b(gate77inter1), .O(N406));

  xor2  gate231(.a(N351), .b(N319), .O(gate78inter0));
  nand2 gate232(.a(gate78inter0), .b(s_4), .O(gate78inter1));
  and2  gate233(.a(N351), .b(N319), .O(gate78inter2));
  inv1  gate234(.a(s_4), .O(gate78inter3));
  inv1  gate235(.a(s_5), .O(gate78inter4));
  nand2 gate236(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate237(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate238(.a(N319), .O(gate78inter7));
  inv1  gate239(.a(N351), .O(gate78inter8));
  nand2 gate240(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate241(.a(s_5), .b(gate78inter3), .O(gate78inter10));
  nor2  gate242(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate243(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate244(.a(gate78inter12), .b(gate78inter1), .O(N419));
xor2 gate79( .a(N320), .b(N352), .O(N432) );
xor2 gate80( .a(N321), .b(N353), .O(N445) );
inv1 gate81( .a(N354), .O(N554) );
inv1 gate82( .a(N367), .O(N555) );
inv1 gate83( .a(N380), .O(N556) );
inv1 gate84( .a(N354), .O(N557) );
inv1 gate85( .a(N367), .O(N558) );
inv1 gate86( .a(N393), .O(N559) );
inv1 gate87( .a(N354), .O(N560) );
inv1 gate88( .a(N380), .O(N561) );
inv1 gate89( .a(N393), .O(N562) );
inv1 gate90( .a(N367), .O(N563) );
inv1 gate91( .a(N380), .O(N564) );
inv1 gate92( .a(N393), .O(N565) );
inv1 gate93( .a(N419), .O(N566) );
inv1 gate94( .a(N445), .O(N567) );
inv1 gate95( .a(N419), .O(N568) );
inv1 gate96( .a(N432), .O(N569) );
inv1 gate97( .a(N406), .O(N570) );
inv1 gate98( .a(N445), .O(N571) );
inv1 gate99( .a(N406), .O(N572) );
inv1 gate100( .a(N432), .O(N573) );
inv1 gate101( .a(N406), .O(N574) );
inv1 gate102( .a(N419), .O(N575) );
inv1 gate103( .a(N432), .O(N576) );
inv1 gate104( .a(N406), .O(N577) );
inv1 gate105( .a(N419), .O(N578) );
inv1 gate106( .a(N445), .O(N579) );
inv1 gate107( .a(N406), .O(N580) );
inv1 gate108( .a(N432), .O(N581) );
inv1 gate109( .a(N445), .O(N582) );
inv1 gate110( .a(N419), .O(N583) );
inv1 gate111( .a(N432), .O(N584) );
inv1 gate112( .a(N445), .O(N585) );
inv1 gate113( .a(N367), .O(N586) );
inv1 gate114( .a(N393), .O(N587) );
inv1 gate115( .a(N367), .O(N588) );
inv1 gate116( .a(N380), .O(N589) );
inv1 gate117( .a(N354), .O(N590) );
inv1 gate118( .a(N393), .O(N591) );
inv1 gate119( .a(N354), .O(N592) );
inv1 gate120( .a(N380), .O(N593) );
and4 gate121( .a(N554), .b(N555), .c(N556), .d(N393), .O(N594) );
and4 gate122( .a(N557), .b(N558), .c(N380), .d(N559), .O(N595) );
and4 gate123( .a(N560), .b(N367), .c(N561), .d(N562), .O(N596) );
and4 gate124( .a(N354), .b(N563), .c(N564), .d(N565), .O(N597) );
and4 gate125( .a(N574), .b(N575), .c(N576), .d(N445), .O(N598) );
and4 gate126( .a(N577), .b(N578), .c(N432), .d(N579), .O(N599) );
and4 gate127( .a(N580), .b(N419), .c(N581), .d(N582), .O(N600) );
and4 gate128( .a(N406), .b(N583), .c(N584), .d(N585), .O(N601) );
or4 gate129( .a(N594), .b(N595), .c(N596), .d(N597), .O(N602) );
or4 gate130( .a(N598), .b(N599), .c(N600), .d(N601), .O(N607) );
and5 gate131( .a(N406), .b(N566), .c(N432), .d(N567), .e(N602), .O(N620) );
and5 gate132( .a(N406), .b(N568), .c(N569), .d(N445), .e(N602), .O(N625) );
and5 gate133( .a(N570), .b(N419), .c(N432), .d(N571), .e(N602), .O(N630) );
and5 gate134( .a(N572), .b(N419), .c(N573), .d(N445), .e(N602), .O(N635) );
and5 gate135( .a(N354), .b(N586), .c(N380), .d(N587), .e(N607), .O(N640) );
and5 gate136( .a(N354), .b(N588), .c(N589), .d(N393), .e(N607), .O(N645) );
and5 gate137( .a(N590), .b(N367), .c(N380), .d(N591), .e(N607), .O(N650) );
and5 gate138( .a(N592), .b(N367), .c(N593), .d(N393), .e(N607), .O(N655) );
and2 gate139( .a(N354), .b(N620), .O(N692) );
and2 gate140( .a(N367), .b(N620), .O(N693) );
and2 gate141( .a(N380), .b(N620), .O(N694) );
and2 gate142( .a(N393), .b(N620), .O(N695) );
and2 gate143( .a(N354), .b(N625), .O(N696) );
and2 gate144( .a(N367), .b(N625), .O(N697) );
and2 gate145( .a(N380), .b(N625), .O(N698) );
and2 gate146( .a(N393), .b(N625), .O(N699) );
and2 gate147( .a(N354), .b(N630), .O(N700) );
and2 gate148( .a(N367), .b(N630), .O(N701) );
and2 gate149( .a(N380), .b(N630), .O(N702) );
and2 gate150( .a(N393), .b(N630), .O(N703) );
and2 gate151( .a(N354), .b(N635), .O(N704) );
and2 gate152( .a(N367), .b(N635), .O(N705) );
and2 gate153( .a(N380), .b(N635), .O(N706) );
and2 gate154( .a(N393), .b(N635), .O(N707) );
and2 gate155( .a(N406), .b(N640), .O(N708) );
and2 gate156( .a(N419), .b(N640), .O(N709) );
and2 gate157( .a(N432), .b(N640), .O(N710) );
and2 gate158( .a(N445), .b(N640), .O(N711) );
and2 gate159( .a(N406), .b(N645), .O(N712) );
and2 gate160( .a(N419), .b(N645), .O(N713) );
and2 gate161( .a(N432), .b(N645), .O(N714) );
and2 gate162( .a(N445), .b(N645), .O(N715) );
and2 gate163( .a(N406), .b(N650), .O(N716) );
and2 gate164( .a(N419), .b(N650), .O(N717) );
and2 gate165( .a(N432), .b(N650), .O(N718) );
and2 gate166( .a(N445), .b(N650), .O(N719) );
and2 gate167( .a(N406), .b(N655), .O(N720) );
and2 gate168( .a(N419), .b(N655), .O(N721) );
and2 gate169( .a(N432), .b(N655), .O(N722) );
and2 gate170( .a(N445), .b(N655), .O(N723) );
xor2 gate171( .a(N1), .b(N692), .O(N724) );

  xor2  gate581(.a(N693), .b(N5), .O(gate172inter0));
  nand2 gate582(.a(gate172inter0), .b(s_54), .O(gate172inter1));
  and2  gate583(.a(N693), .b(N5), .O(gate172inter2));
  inv1  gate584(.a(s_54), .O(gate172inter3));
  inv1  gate585(.a(s_55), .O(gate172inter4));
  nand2 gate586(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate587(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate588(.a(N5), .O(gate172inter7));
  inv1  gate589(.a(N693), .O(gate172inter8));
  nand2 gate590(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate591(.a(s_55), .b(gate172inter3), .O(gate172inter10));
  nor2  gate592(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate593(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate594(.a(gate172inter12), .b(gate172inter1), .O(N725));

  xor2  gate427(.a(N694), .b(N9), .O(gate173inter0));
  nand2 gate428(.a(gate173inter0), .b(s_32), .O(gate173inter1));
  and2  gate429(.a(N694), .b(N9), .O(gate173inter2));
  inv1  gate430(.a(s_32), .O(gate173inter3));
  inv1  gate431(.a(s_33), .O(gate173inter4));
  nand2 gate432(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate433(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate434(.a(N9), .O(gate173inter7));
  inv1  gate435(.a(N694), .O(gate173inter8));
  nand2 gate436(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate437(.a(s_33), .b(gate173inter3), .O(gate173inter10));
  nor2  gate438(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate439(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate440(.a(gate173inter12), .b(gate173inter1), .O(N726));

  xor2  gate259(.a(N695), .b(N13), .O(gate174inter0));
  nand2 gate260(.a(gate174inter0), .b(s_8), .O(gate174inter1));
  and2  gate261(.a(N695), .b(N13), .O(gate174inter2));
  inv1  gate262(.a(s_8), .O(gate174inter3));
  inv1  gate263(.a(s_9), .O(gate174inter4));
  nand2 gate264(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate265(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate266(.a(N13), .O(gate174inter7));
  inv1  gate267(.a(N695), .O(gate174inter8));
  nand2 gate268(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate269(.a(s_9), .b(gate174inter3), .O(gate174inter10));
  nor2  gate270(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate271(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate272(.a(gate174inter12), .b(gate174inter1), .O(N727));

  xor2  gate665(.a(N696), .b(N17), .O(gate175inter0));
  nand2 gate666(.a(gate175inter0), .b(s_66), .O(gate175inter1));
  and2  gate667(.a(N696), .b(N17), .O(gate175inter2));
  inv1  gate668(.a(s_66), .O(gate175inter3));
  inv1  gate669(.a(s_67), .O(gate175inter4));
  nand2 gate670(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate671(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate672(.a(N17), .O(gate175inter7));
  inv1  gate673(.a(N696), .O(gate175inter8));
  nand2 gate674(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate675(.a(s_67), .b(gate175inter3), .O(gate175inter10));
  nor2  gate676(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate677(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate678(.a(gate175inter12), .b(gate175inter1), .O(N728));
xor2 gate176( .a(N21), .b(N697), .O(N729) );
xor2 gate177( .a(N25), .b(N698), .O(N730) );

  xor2  gate273(.a(N699), .b(N29), .O(gate178inter0));
  nand2 gate274(.a(gate178inter0), .b(s_10), .O(gate178inter1));
  and2  gate275(.a(N699), .b(N29), .O(gate178inter2));
  inv1  gate276(.a(s_10), .O(gate178inter3));
  inv1  gate277(.a(s_11), .O(gate178inter4));
  nand2 gate278(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate279(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate280(.a(N29), .O(gate178inter7));
  inv1  gate281(.a(N699), .O(gate178inter8));
  nand2 gate282(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate283(.a(s_11), .b(gate178inter3), .O(gate178inter10));
  nor2  gate284(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate285(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate286(.a(gate178inter12), .b(gate178inter1), .O(N731));

  xor2  gate763(.a(N700), .b(N33), .O(gate179inter0));
  nand2 gate764(.a(gate179inter0), .b(s_80), .O(gate179inter1));
  and2  gate765(.a(N700), .b(N33), .O(gate179inter2));
  inv1  gate766(.a(s_80), .O(gate179inter3));
  inv1  gate767(.a(s_81), .O(gate179inter4));
  nand2 gate768(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate769(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate770(.a(N33), .O(gate179inter7));
  inv1  gate771(.a(N700), .O(gate179inter8));
  nand2 gate772(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate773(.a(s_81), .b(gate179inter3), .O(gate179inter10));
  nor2  gate774(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate775(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate776(.a(gate179inter12), .b(gate179inter1), .O(N732));
xor2 gate180( .a(N37), .b(N701), .O(N733) );
xor2 gate181( .a(N41), .b(N702), .O(N734) );
xor2 gate182( .a(N45), .b(N703), .O(N735) );

  xor2  gate721(.a(N704), .b(N49), .O(gate183inter0));
  nand2 gate722(.a(gate183inter0), .b(s_74), .O(gate183inter1));
  and2  gate723(.a(N704), .b(N49), .O(gate183inter2));
  inv1  gate724(.a(s_74), .O(gate183inter3));
  inv1  gate725(.a(s_75), .O(gate183inter4));
  nand2 gate726(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate727(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate728(.a(N49), .O(gate183inter7));
  inv1  gate729(.a(N704), .O(gate183inter8));
  nand2 gate730(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate731(.a(s_75), .b(gate183inter3), .O(gate183inter10));
  nor2  gate732(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate733(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate734(.a(gate183inter12), .b(gate183inter1), .O(N736));
xor2 gate184( .a(N53), .b(N705), .O(N737) );

  xor2  gate483(.a(N706), .b(N57), .O(gate185inter0));
  nand2 gate484(.a(gate185inter0), .b(s_40), .O(gate185inter1));
  and2  gate485(.a(N706), .b(N57), .O(gate185inter2));
  inv1  gate486(.a(s_40), .O(gate185inter3));
  inv1  gate487(.a(s_41), .O(gate185inter4));
  nand2 gate488(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate489(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate490(.a(N57), .O(gate185inter7));
  inv1  gate491(.a(N706), .O(gate185inter8));
  nand2 gate492(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate493(.a(s_41), .b(gate185inter3), .O(gate185inter10));
  nor2  gate494(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate495(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate496(.a(gate185inter12), .b(gate185inter1), .O(N738));

  xor2  gate203(.a(N707), .b(N61), .O(gate186inter0));
  nand2 gate204(.a(gate186inter0), .b(s_0), .O(gate186inter1));
  and2  gate205(.a(N707), .b(N61), .O(gate186inter2));
  inv1  gate206(.a(s_0), .O(gate186inter3));
  inv1  gate207(.a(s_1), .O(gate186inter4));
  nand2 gate208(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate209(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate210(.a(N61), .O(gate186inter7));
  inv1  gate211(.a(N707), .O(gate186inter8));
  nand2 gate212(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate213(.a(s_1), .b(gate186inter3), .O(gate186inter10));
  nor2  gate214(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate215(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate216(.a(gate186inter12), .b(gate186inter1), .O(N739));

  xor2  gate315(.a(N708), .b(N65), .O(gate187inter0));
  nand2 gate316(.a(gate187inter0), .b(s_16), .O(gate187inter1));
  and2  gate317(.a(N708), .b(N65), .O(gate187inter2));
  inv1  gate318(.a(s_16), .O(gate187inter3));
  inv1  gate319(.a(s_17), .O(gate187inter4));
  nand2 gate320(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate321(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate322(.a(N65), .O(gate187inter7));
  inv1  gate323(.a(N708), .O(gate187inter8));
  nand2 gate324(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate325(.a(s_17), .b(gate187inter3), .O(gate187inter10));
  nor2  gate326(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate327(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate328(.a(gate187inter12), .b(gate187inter1), .O(N740));
xor2 gate188( .a(N69), .b(N709), .O(N741) );

  xor2  gate301(.a(N710), .b(N73), .O(gate189inter0));
  nand2 gate302(.a(gate189inter0), .b(s_14), .O(gate189inter1));
  and2  gate303(.a(N710), .b(N73), .O(gate189inter2));
  inv1  gate304(.a(s_14), .O(gate189inter3));
  inv1  gate305(.a(s_15), .O(gate189inter4));
  nand2 gate306(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate307(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate308(.a(N73), .O(gate189inter7));
  inv1  gate309(.a(N710), .O(gate189inter8));
  nand2 gate310(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate311(.a(s_15), .b(gate189inter3), .O(gate189inter10));
  nor2  gate312(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate313(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate314(.a(gate189inter12), .b(gate189inter1), .O(N742));

  xor2  gate693(.a(N711), .b(N77), .O(gate190inter0));
  nand2 gate694(.a(gate190inter0), .b(s_70), .O(gate190inter1));
  and2  gate695(.a(N711), .b(N77), .O(gate190inter2));
  inv1  gate696(.a(s_70), .O(gate190inter3));
  inv1  gate697(.a(s_71), .O(gate190inter4));
  nand2 gate698(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate699(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate700(.a(N77), .O(gate190inter7));
  inv1  gate701(.a(N711), .O(gate190inter8));
  nand2 gate702(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate703(.a(s_71), .b(gate190inter3), .O(gate190inter10));
  nor2  gate704(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate705(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate706(.a(gate190inter12), .b(gate190inter1), .O(N743));
xor2 gate191( .a(N81), .b(N712), .O(N744) );
xor2 gate192( .a(N85), .b(N713), .O(N745) );
xor2 gate193( .a(N89), .b(N714), .O(N746) );
xor2 gate194( .a(N93), .b(N715), .O(N747) );

  xor2  gate623(.a(N716), .b(N97), .O(gate195inter0));
  nand2 gate624(.a(gate195inter0), .b(s_60), .O(gate195inter1));
  and2  gate625(.a(N716), .b(N97), .O(gate195inter2));
  inv1  gate626(.a(s_60), .O(gate195inter3));
  inv1  gate627(.a(s_61), .O(gate195inter4));
  nand2 gate628(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate629(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate630(.a(N97), .O(gate195inter7));
  inv1  gate631(.a(N716), .O(gate195inter8));
  nand2 gate632(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate633(.a(s_61), .b(gate195inter3), .O(gate195inter10));
  nor2  gate634(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate635(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate636(.a(gate195inter12), .b(gate195inter1), .O(N748));

  xor2  gate497(.a(N717), .b(N101), .O(gate196inter0));
  nand2 gate498(.a(gate196inter0), .b(s_42), .O(gate196inter1));
  and2  gate499(.a(N717), .b(N101), .O(gate196inter2));
  inv1  gate500(.a(s_42), .O(gate196inter3));
  inv1  gate501(.a(s_43), .O(gate196inter4));
  nand2 gate502(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate503(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate504(.a(N101), .O(gate196inter7));
  inv1  gate505(.a(N717), .O(gate196inter8));
  nand2 gate506(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate507(.a(s_43), .b(gate196inter3), .O(gate196inter10));
  nor2  gate508(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate509(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate510(.a(gate196inter12), .b(gate196inter1), .O(N749));

  xor2  gate385(.a(N718), .b(N105), .O(gate197inter0));
  nand2 gate386(.a(gate197inter0), .b(s_26), .O(gate197inter1));
  and2  gate387(.a(N718), .b(N105), .O(gate197inter2));
  inv1  gate388(.a(s_26), .O(gate197inter3));
  inv1  gate389(.a(s_27), .O(gate197inter4));
  nand2 gate390(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate391(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate392(.a(N105), .O(gate197inter7));
  inv1  gate393(.a(N718), .O(gate197inter8));
  nand2 gate394(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate395(.a(s_27), .b(gate197inter3), .O(gate197inter10));
  nor2  gate396(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate397(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate398(.a(gate197inter12), .b(gate197inter1), .O(N750));
xor2 gate198( .a(N109), .b(N719), .O(N751) );
xor2 gate199( .a(N113), .b(N720), .O(N752) );
xor2 gate200( .a(N117), .b(N721), .O(N753) );

  xor2  gate539(.a(N722), .b(N121), .O(gate201inter0));
  nand2 gate540(.a(gate201inter0), .b(s_48), .O(gate201inter1));
  and2  gate541(.a(N722), .b(N121), .O(gate201inter2));
  inv1  gate542(.a(s_48), .O(gate201inter3));
  inv1  gate543(.a(s_49), .O(gate201inter4));
  nand2 gate544(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate545(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate546(.a(N121), .O(gate201inter7));
  inv1  gate547(.a(N722), .O(gate201inter8));
  nand2 gate548(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate549(.a(s_49), .b(gate201inter3), .O(gate201inter10));
  nor2  gate550(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate551(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate552(.a(gate201inter12), .b(gate201inter1), .O(N754));
xor2 gate202( .a(N125), .b(N723), .O(N755) );

endmodule