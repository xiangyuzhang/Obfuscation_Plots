module c432 (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
             N430,N431,N432);
input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
      N99,N102,N105,N108,N112,N115;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61;
output N223,N329,N370,N421,N430,N431,N432;
wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12;


inv1 gate1( .a(N1), .O(N118) );
inv1 gate2( .a(N4), .O(N119) );
inv1 gate3( .a(N11), .O(N122) );
inv1 gate4( .a(N17), .O(N123) );
inv1 gate5( .a(N24), .O(N126) );
inv1 gate6( .a(N30), .O(N127) );
inv1 gate7( .a(N37), .O(N130) );
inv1 gate8( .a(N43), .O(N131) );
inv1 gate9( .a(N50), .O(N134) );
inv1 gate10( .a(N56), .O(N135) );
inv1 gate11( .a(N63), .O(N138) );
inv1 gate12( .a(N69), .O(N139) );
inv1 gate13( .a(N76), .O(N142) );
inv1 gate14( .a(N82), .O(N143) );
inv1 gate15( .a(N89), .O(N146) );
inv1 gate16( .a(N95), .O(N147) );
inv1 gate17( .a(N102), .O(N150) );
inv1 gate18( .a(N108), .O(N151) );

  xor2  gate245(.a(N4), .b(N118), .O(gate19inter0));
  nand2 gate246(.a(gate19inter0), .b(s_12), .O(gate19inter1));
  and2  gate247(.a(N4), .b(N118), .O(gate19inter2));
  inv1  gate248(.a(s_12), .O(gate19inter3));
  inv1  gate249(.a(s_13), .O(gate19inter4));
  nand2 gate250(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate251(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate252(.a(N118), .O(gate19inter7));
  inv1  gate253(.a(N4), .O(gate19inter8));
  nand2 gate254(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate255(.a(s_13), .b(gate19inter3), .O(gate19inter10));
  nor2  gate256(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate257(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate258(.a(gate19inter12), .b(gate19inter1), .O(N154));

  xor2  gate329(.a(N119), .b(N8), .O(gate20inter0));
  nand2 gate330(.a(gate20inter0), .b(s_24), .O(gate20inter1));
  and2  gate331(.a(N119), .b(N8), .O(gate20inter2));
  inv1  gate332(.a(s_24), .O(gate20inter3));
  inv1  gate333(.a(s_25), .O(gate20inter4));
  nand2 gate334(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate335(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate336(.a(N8), .O(gate20inter7));
  inv1  gate337(.a(N119), .O(gate20inter8));
  nand2 gate338(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate339(.a(s_25), .b(gate20inter3), .O(gate20inter10));
  nor2  gate340(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate341(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate342(.a(gate20inter12), .b(gate20inter1), .O(N157));
nor2 gate21( .a(N14), .b(N119), .O(N158) );
nand2 gate22( .a(N122), .b(N17), .O(N159) );

  xor2  gate441(.a(N30), .b(N126), .O(gate23inter0));
  nand2 gate442(.a(gate23inter0), .b(s_40), .O(gate23inter1));
  and2  gate443(.a(N30), .b(N126), .O(gate23inter2));
  inv1  gate444(.a(s_40), .O(gate23inter3));
  inv1  gate445(.a(s_41), .O(gate23inter4));
  nand2 gate446(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate447(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate448(.a(N126), .O(gate23inter7));
  inv1  gate449(.a(N30), .O(gate23inter8));
  nand2 gate450(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate451(.a(s_41), .b(gate23inter3), .O(gate23inter10));
  nor2  gate452(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate453(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate454(.a(gate23inter12), .b(gate23inter1), .O(N162));
nand2 gate24( .a(N130), .b(N43), .O(N165) );
nand2 gate25( .a(N134), .b(N56), .O(N168) );
nand2 gate26( .a(N138), .b(N69), .O(N171) );

  xor2  gate427(.a(N82), .b(N142), .O(gate27inter0));
  nand2 gate428(.a(gate27inter0), .b(s_38), .O(gate27inter1));
  and2  gate429(.a(N82), .b(N142), .O(gate27inter2));
  inv1  gate430(.a(s_38), .O(gate27inter3));
  inv1  gate431(.a(s_39), .O(gate27inter4));
  nand2 gate432(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate433(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate434(.a(N142), .O(gate27inter7));
  inv1  gate435(.a(N82), .O(gate27inter8));
  nand2 gate436(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate437(.a(s_39), .b(gate27inter3), .O(gate27inter10));
  nor2  gate438(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate439(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate440(.a(gate27inter12), .b(gate27inter1), .O(N174));
nand2 gate28( .a(N146), .b(N95), .O(N177) );
nand2 gate29( .a(N150), .b(N108), .O(N180) );

  xor2  gate539(.a(N123), .b(N21), .O(gate30inter0));
  nand2 gate540(.a(gate30inter0), .b(s_54), .O(gate30inter1));
  and2  gate541(.a(N123), .b(N21), .O(gate30inter2));
  inv1  gate542(.a(s_54), .O(gate30inter3));
  inv1  gate543(.a(s_55), .O(gate30inter4));
  nand2 gate544(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate545(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate546(.a(N21), .O(gate30inter7));
  inv1  gate547(.a(N123), .O(gate30inter8));
  nand2 gate548(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate549(.a(s_55), .b(gate30inter3), .O(gate30inter10));
  nor2  gate550(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate551(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate552(.a(gate30inter12), .b(gate30inter1), .O(N183));
nor2 gate31( .a(N27), .b(N123), .O(N184) );
nor2 gate32( .a(N34), .b(N127), .O(N185) );
nor2 gate33( .a(N40), .b(N127), .O(N186) );

  xor2  gate497(.a(N131), .b(N47), .O(gate34inter0));
  nand2 gate498(.a(gate34inter0), .b(s_48), .O(gate34inter1));
  and2  gate499(.a(N131), .b(N47), .O(gate34inter2));
  inv1  gate500(.a(s_48), .O(gate34inter3));
  inv1  gate501(.a(s_49), .O(gate34inter4));
  nand2 gate502(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate503(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate504(.a(N47), .O(gate34inter7));
  inv1  gate505(.a(N131), .O(gate34inter8));
  nand2 gate506(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate507(.a(s_49), .b(gate34inter3), .O(gate34inter10));
  nor2  gate508(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate509(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate510(.a(gate34inter12), .b(gate34inter1), .O(N187));

  xor2  gate483(.a(N131), .b(N53), .O(gate35inter0));
  nand2 gate484(.a(gate35inter0), .b(s_46), .O(gate35inter1));
  and2  gate485(.a(N131), .b(N53), .O(gate35inter2));
  inv1  gate486(.a(s_46), .O(gate35inter3));
  inv1  gate487(.a(s_47), .O(gate35inter4));
  nand2 gate488(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate489(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate490(.a(N53), .O(gate35inter7));
  inv1  gate491(.a(N131), .O(gate35inter8));
  nand2 gate492(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate493(.a(s_47), .b(gate35inter3), .O(gate35inter10));
  nor2  gate494(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate495(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate496(.a(gate35inter12), .b(gate35inter1), .O(N188));
nor2 gate36( .a(N60), .b(N135), .O(N189) );
nor2 gate37( .a(N66), .b(N135), .O(N190) );
nor2 gate38( .a(N73), .b(N139), .O(N191) );
nor2 gate39( .a(N79), .b(N139), .O(N192) );

  xor2  gate469(.a(N143), .b(N86), .O(gate40inter0));
  nand2 gate470(.a(gate40inter0), .b(s_44), .O(gate40inter1));
  and2  gate471(.a(N143), .b(N86), .O(gate40inter2));
  inv1  gate472(.a(s_44), .O(gate40inter3));
  inv1  gate473(.a(s_45), .O(gate40inter4));
  nand2 gate474(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate475(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate476(.a(N86), .O(gate40inter7));
  inv1  gate477(.a(N143), .O(gate40inter8));
  nand2 gate478(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate479(.a(s_45), .b(gate40inter3), .O(gate40inter10));
  nor2  gate480(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate481(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate482(.a(gate40inter12), .b(gate40inter1), .O(N193));
nor2 gate41( .a(N92), .b(N143), .O(N194) );
nor2 gate42( .a(N99), .b(N147), .O(N195) );

  xor2  gate287(.a(N147), .b(N105), .O(gate43inter0));
  nand2 gate288(.a(gate43inter0), .b(s_18), .O(gate43inter1));
  and2  gate289(.a(N147), .b(N105), .O(gate43inter2));
  inv1  gate290(.a(s_18), .O(gate43inter3));
  inv1  gate291(.a(s_19), .O(gate43inter4));
  nand2 gate292(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate293(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate294(.a(N105), .O(gate43inter7));
  inv1  gate295(.a(N147), .O(gate43inter8));
  nand2 gate296(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate297(.a(s_19), .b(gate43inter3), .O(gate43inter10));
  nor2  gate298(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate299(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate300(.a(gate43inter12), .b(gate43inter1), .O(N196));
nor2 gate44( .a(N112), .b(N151), .O(N197) );
nor2 gate45( .a(N115), .b(N151), .O(N198) );
and9 gate46( .a(N154), .b(N159), .c(N162), .d(N165), .e(N168), .f(N171), .g(N174), .h(N177), .i(N180), .O(N199) );
inv1 gate47( .a(N199), .O(N203) );
inv1 gate48( .a(N199), .O(N213) );
inv1 gate49( .a(N199), .O(N223) );
xor2 gate50( .a(N203), .b(N154), .O(N224) );
xor2 gate51( .a(N203), .b(N159), .O(N227) );
xor2 gate52( .a(N203), .b(N162), .O(N230) );
xor2 gate53( .a(N203), .b(N165), .O(N233) );
xor2 gate54( .a(N203), .b(N168), .O(N236) );

  xor2  gate371(.a(N171), .b(N203), .O(gate55inter0));
  nand2 gate372(.a(gate55inter0), .b(s_30), .O(gate55inter1));
  and2  gate373(.a(N171), .b(N203), .O(gate55inter2));
  inv1  gate374(.a(s_30), .O(gate55inter3));
  inv1  gate375(.a(s_31), .O(gate55inter4));
  nand2 gate376(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate377(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate378(.a(N203), .O(gate55inter7));
  inv1  gate379(.a(N171), .O(gate55inter8));
  nand2 gate380(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate381(.a(s_31), .b(gate55inter3), .O(gate55inter10));
  nor2  gate382(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate383(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate384(.a(gate55inter12), .b(gate55inter1), .O(N239));

  xor2  gate343(.a(N213), .b(N1), .O(gate56inter0));
  nand2 gate344(.a(gate56inter0), .b(s_26), .O(gate56inter1));
  and2  gate345(.a(N213), .b(N1), .O(gate56inter2));
  inv1  gate346(.a(s_26), .O(gate56inter3));
  inv1  gate347(.a(s_27), .O(gate56inter4));
  nand2 gate348(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate349(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate350(.a(N1), .O(gate56inter7));
  inv1  gate351(.a(N213), .O(gate56inter8));
  nand2 gate352(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate353(.a(s_27), .b(gate56inter3), .O(gate56inter10));
  nor2  gate354(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate355(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate356(.a(gate56inter12), .b(gate56inter1), .O(N242));

  xor2  gate189(.a(N174), .b(N203), .O(gate57inter0));
  nand2 gate190(.a(gate57inter0), .b(s_4), .O(gate57inter1));
  and2  gate191(.a(N174), .b(N203), .O(gate57inter2));
  inv1  gate192(.a(s_4), .O(gate57inter3));
  inv1  gate193(.a(s_5), .O(gate57inter4));
  nand2 gate194(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate195(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate196(.a(N203), .O(gate57inter7));
  inv1  gate197(.a(N174), .O(gate57inter8));
  nand2 gate198(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate199(.a(s_5), .b(gate57inter3), .O(gate57inter10));
  nor2  gate200(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate201(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate202(.a(gate57inter12), .b(gate57inter1), .O(N243));

  xor2  gate357(.a(N11), .b(N213), .O(gate58inter0));
  nand2 gate358(.a(gate58inter0), .b(s_28), .O(gate58inter1));
  and2  gate359(.a(N11), .b(N213), .O(gate58inter2));
  inv1  gate360(.a(s_28), .O(gate58inter3));
  inv1  gate361(.a(s_29), .O(gate58inter4));
  nand2 gate362(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate363(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate364(.a(N213), .O(gate58inter7));
  inv1  gate365(.a(N11), .O(gate58inter8));
  nand2 gate366(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate367(.a(s_29), .b(gate58inter3), .O(gate58inter10));
  nor2  gate368(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate369(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate370(.a(gate58inter12), .b(gate58inter1), .O(N246));
xor2 gate59( .a(N203), .b(N177), .O(N247) );
nand2 gate60( .a(N213), .b(N24), .O(N250) );
xor2 gate61( .a(N203), .b(N180), .O(N251) );
nand2 gate62( .a(N213), .b(N37), .O(N254) );
nand2 gate63( .a(N213), .b(N50), .O(N255) );
nand2 gate64( .a(N213), .b(N63), .O(N256) );
nand2 gate65( .a(N213), .b(N76), .O(N257) );
nand2 gate66( .a(N213), .b(N89), .O(N258) );
nand2 gate67( .a(N213), .b(N102), .O(N259) );
nand2 gate68( .a(N224), .b(N157), .O(N260) );
nand2 gate69( .a(N224), .b(N158), .O(N263) );
nand2 gate70( .a(N227), .b(N183), .O(N264) );
nand2 gate71( .a(N230), .b(N185), .O(N267) );

  xor2  gate553(.a(N187), .b(N233), .O(gate72inter0));
  nand2 gate554(.a(gate72inter0), .b(s_56), .O(gate72inter1));
  and2  gate555(.a(N187), .b(N233), .O(gate72inter2));
  inv1  gate556(.a(s_56), .O(gate72inter3));
  inv1  gate557(.a(s_57), .O(gate72inter4));
  nand2 gate558(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate559(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate560(.a(N233), .O(gate72inter7));
  inv1  gate561(.a(N187), .O(gate72inter8));
  nand2 gate562(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate563(.a(s_57), .b(gate72inter3), .O(gate72inter10));
  nor2  gate564(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate565(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate566(.a(gate72inter12), .b(gate72inter1), .O(N270));
nand2 gate73( .a(N236), .b(N189), .O(N273) );
nand2 gate74( .a(N239), .b(N191), .O(N276) );

  xor2  gate231(.a(N193), .b(N243), .O(gate75inter0));
  nand2 gate232(.a(gate75inter0), .b(s_10), .O(gate75inter1));
  and2  gate233(.a(N193), .b(N243), .O(gate75inter2));
  inv1  gate234(.a(s_10), .O(gate75inter3));
  inv1  gate235(.a(s_11), .O(gate75inter4));
  nand2 gate236(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate237(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate238(.a(N243), .O(gate75inter7));
  inv1  gate239(.a(N193), .O(gate75inter8));
  nand2 gate240(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate241(.a(s_11), .b(gate75inter3), .O(gate75inter10));
  nor2  gate242(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate243(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate244(.a(gate75inter12), .b(gate75inter1), .O(N279));
nand2 gate76( .a(N247), .b(N195), .O(N282) );

  xor2  gate525(.a(N197), .b(N251), .O(gate77inter0));
  nand2 gate526(.a(gate77inter0), .b(s_52), .O(gate77inter1));
  and2  gate527(.a(N197), .b(N251), .O(gate77inter2));
  inv1  gate528(.a(s_52), .O(gate77inter3));
  inv1  gate529(.a(s_53), .O(gate77inter4));
  nand2 gate530(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate531(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate532(.a(N251), .O(gate77inter7));
  inv1  gate533(.a(N197), .O(gate77inter8));
  nand2 gate534(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate535(.a(s_53), .b(gate77inter3), .O(gate77inter10));
  nor2  gate536(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate537(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate538(.a(gate77inter12), .b(gate77inter1), .O(N285));

  xor2  gate567(.a(N184), .b(N227), .O(gate78inter0));
  nand2 gate568(.a(gate78inter0), .b(s_58), .O(gate78inter1));
  and2  gate569(.a(N184), .b(N227), .O(gate78inter2));
  inv1  gate570(.a(s_58), .O(gate78inter3));
  inv1  gate571(.a(s_59), .O(gate78inter4));
  nand2 gate572(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate573(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate574(.a(N227), .O(gate78inter7));
  inv1  gate575(.a(N184), .O(gate78inter8));
  nand2 gate576(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate577(.a(s_59), .b(gate78inter3), .O(gate78inter10));
  nor2  gate578(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate579(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate580(.a(gate78inter12), .b(gate78inter1), .O(N288));
nand2 gate79( .a(N230), .b(N186), .O(N289) );
nand2 gate80( .a(N233), .b(N188), .O(N290) );

  xor2  gate455(.a(N190), .b(N236), .O(gate81inter0));
  nand2 gate456(.a(gate81inter0), .b(s_42), .O(gate81inter1));
  and2  gate457(.a(N190), .b(N236), .O(gate81inter2));
  inv1  gate458(.a(s_42), .O(gate81inter3));
  inv1  gate459(.a(s_43), .O(gate81inter4));
  nand2 gate460(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate461(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate462(.a(N236), .O(gate81inter7));
  inv1  gate463(.a(N190), .O(gate81inter8));
  nand2 gate464(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate465(.a(s_43), .b(gate81inter3), .O(gate81inter10));
  nor2  gate466(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate467(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate468(.a(gate81inter12), .b(gate81inter1), .O(N291));
nand2 gate82( .a(N239), .b(N192), .O(N292) );

  xor2  gate301(.a(N194), .b(N243), .O(gate83inter0));
  nand2 gate302(.a(gate83inter0), .b(s_20), .O(gate83inter1));
  and2  gate303(.a(N194), .b(N243), .O(gate83inter2));
  inv1  gate304(.a(s_20), .O(gate83inter3));
  inv1  gate305(.a(s_21), .O(gate83inter4));
  nand2 gate306(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate307(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate308(.a(N243), .O(gate83inter7));
  inv1  gate309(.a(N194), .O(gate83inter8));
  nand2 gate310(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate311(.a(s_21), .b(gate83inter3), .O(gate83inter10));
  nor2  gate312(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate313(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate314(.a(gate83inter12), .b(gate83inter1), .O(N293));

  xor2  gate217(.a(N196), .b(N247), .O(gate84inter0));
  nand2 gate218(.a(gate84inter0), .b(s_8), .O(gate84inter1));
  and2  gate219(.a(N196), .b(N247), .O(gate84inter2));
  inv1  gate220(.a(s_8), .O(gate84inter3));
  inv1  gate221(.a(s_9), .O(gate84inter4));
  nand2 gate222(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate223(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate224(.a(N247), .O(gate84inter7));
  inv1  gate225(.a(N196), .O(gate84inter8));
  nand2 gate226(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate227(.a(s_9), .b(gate84inter3), .O(gate84inter10));
  nor2  gate228(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate229(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate230(.a(gate84inter12), .b(gate84inter1), .O(N294));
nand2 gate85( .a(N251), .b(N198), .O(N295) );
and9 gate86( .a(N260), .b(N264), .c(N267), .d(N270), .e(N273), .f(N276), .g(N279), .h(N282), .i(N285), .O(N296) );
inv1 gate87( .a(N263), .O(N300) );
inv1 gate88( .a(N288), .O(N301) );
inv1 gate89( .a(N289), .O(N302) );
inv1 gate90( .a(N290), .O(N303) );
inv1 gate91( .a(N291), .O(N304) );
inv1 gate92( .a(N292), .O(N305) );
inv1 gate93( .a(N293), .O(N306) );
inv1 gate94( .a(N294), .O(N307) );
inv1 gate95( .a(N295), .O(N308) );
inv1 gate96( .a(N296), .O(N309) );
inv1 gate97( .a(N296), .O(N319) );
inv1 gate98( .a(N296), .O(N329) );
xor2 gate99( .a(N309), .b(N260), .O(N330) );
xor2 gate100( .a(N309), .b(N264), .O(N331) );
xor2 gate101( .a(N309), .b(N267), .O(N332) );
xor2 gate102( .a(N309), .b(N270), .O(N333) );

  xor2  gate273(.a(N319), .b(N8), .O(gate103inter0));
  nand2 gate274(.a(gate103inter0), .b(s_16), .O(gate103inter1));
  and2  gate275(.a(N319), .b(N8), .O(gate103inter2));
  inv1  gate276(.a(s_16), .O(gate103inter3));
  inv1  gate277(.a(s_17), .O(gate103inter4));
  nand2 gate278(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate279(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate280(.a(N8), .O(gate103inter7));
  inv1  gate281(.a(N319), .O(gate103inter8));
  nand2 gate282(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate283(.a(s_17), .b(gate103inter3), .O(gate103inter10));
  nor2  gate284(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate285(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate286(.a(gate103inter12), .b(gate103inter1), .O(N334));
xor2 gate104( .a(N309), .b(N273), .O(N335) );
nand2 gate105( .a(N319), .b(N21), .O(N336) );
xor2 gate106( .a(N309), .b(N276), .O(N337) );
nand2 gate107( .a(N319), .b(N34), .O(N338) );
xor2 gate108( .a(N309), .b(N279), .O(N339) );
nand2 gate109( .a(N319), .b(N47), .O(N340) );
xor2 gate110( .a(N309), .b(N282), .O(N341) );
nand2 gate111( .a(N319), .b(N60), .O(N342) );
xor2 gate112( .a(N309), .b(N285), .O(N343) );
nand2 gate113( .a(N319), .b(N73), .O(N344) );
nand2 gate114( .a(N319), .b(N86), .O(N345) );

  xor2  gate315(.a(N99), .b(N319), .O(gate115inter0));
  nand2 gate316(.a(gate115inter0), .b(s_22), .O(gate115inter1));
  and2  gate317(.a(N99), .b(N319), .O(gate115inter2));
  inv1  gate318(.a(s_22), .O(gate115inter3));
  inv1  gate319(.a(s_23), .O(gate115inter4));
  nand2 gate320(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate321(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate322(.a(N319), .O(gate115inter7));
  inv1  gate323(.a(N99), .O(gate115inter8));
  nand2 gate324(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate325(.a(s_23), .b(gate115inter3), .O(gate115inter10));
  nor2  gate326(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate327(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate328(.a(gate115inter12), .b(gate115inter1), .O(N346));
nand2 gate116( .a(N319), .b(N112), .O(N347) );
nand2 gate117( .a(N330), .b(N300), .O(N348) );

  xor2  gate399(.a(N301), .b(N331), .O(gate118inter0));
  nand2 gate400(.a(gate118inter0), .b(s_34), .O(gate118inter1));
  and2  gate401(.a(N301), .b(N331), .O(gate118inter2));
  inv1  gate402(.a(s_34), .O(gate118inter3));
  inv1  gate403(.a(s_35), .O(gate118inter4));
  nand2 gate404(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate405(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate406(.a(N331), .O(gate118inter7));
  inv1  gate407(.a(N301), .O(gate118inter8));
  nand2 gate408(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate409(.a(s_35), .b(gate118inter3), .O(gate118inter10));
  nor2  gate410(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate411(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate412(.a(gate118inter12), .b(gate118inter1), .O(N349));
nand2 gate119( .a(N332), .b(N302), .O(N350) );
nand2 gate120( .a(N333), .b(N303), .O(N351) );

  xor2  gate413(.a(N304), .b(N335), .O(gate121inter0));
  nand2 gate414(.a(gate121inter0), .b(s_36), .O(gate121inter1));
  and2  gate415(.a(N304), .b(N335), .O(gate121inter2));
  inv1  gate416(.a(s_36), .O(gate121inter3));
  inv1  gate417(.a(s_37), .O(gate121inter4));
  nand2 gate418(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate419(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate420(.a(N335), .O(gate121inter7));
  inv1  gate421(.a(N304), .O(gate121inter8));
  nand2 gate422(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate423(.a(s_37), .b(gate121inter3), .O(gate121inter10));
  nor2  gate424(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate425(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate426(.a(gate121inter12), .b(gate121inter1), .O(N352));

  xor2  gate581(.a(N305), .b(N337), .O(gate122inter0));
  nand2 gate582(.a(gate122inter0), .b(s_60), .O(gate122inter1));
  and2  gate583(.a(N305), .b(N337), .O(gate122inter2));
  inv1  gate584(.a(s_60), .O(gate122inter3));
  inv1  gate585(.a(s_61), .O(gate122inter4));
  nand2 gate586(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate587(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate588(.a(N337), .O(gate122inter7));
  inv1  gate589(.a(N305), .O(gate122inter8));
  nand2 gate590(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate591(.a(s_61), .b(gate122inter3), .O(gate122inter10));
  nor2  gate592(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate593(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate594(.a(gate122inter12), .b(gate122inter1), .O(N353));

  xor2  gate385(.a(N306), .b(N339), .O(gate123inter0));
  nand2 gate386(.a(gate123inter0), .b(s_32), .O(gate123inter1));
  and2  gate387(.a(N306), .b(N339), .O(gate123inter2));
  inv1  gate388(.a(s_32), .O(gate123inter3));
  inv1  gate389(.a(s_33), .O(gate123inter4));
  nand2 gate390(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate391(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate392(.a(N339), .O(gate123inter7));
  inv1  gate393(.a(N306), .O(gate123inter8));
  nand2 gate394(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate395(.a(s_33), .b(gate123inter3), .O(gate123inter10));
  nor2  gate396(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate397(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate398(.a(gate123inter12), .b(gate123inter1), .O(N354));

  xor2  gate175(.a(N307), .b(N341), .O(gate124inter0));
  nand2 gate176(.a(gate124inter0), .b(s_2), .O(gate124inter1));
  and2  gate177(.a(N307), .b(N341), .O(gate124inter2));
  inv1  gate178(.a(s_2), .O(gate124inter3));
  inv1  gate179(.a(s_3), .O(gate124inter4));
  nand2 gate180(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate181(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate182(.a(N341), .O(gate124inter7));
  inv1  gate183(.a(N307), .O(gate124inter8));
  nand2 gate184(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate185(.a(s_3), .b(gate124inter3), .O(gate124inter10));
  nor2  gate186(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate187(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate188(.a(gate124inter12), .b(gate124inter1), .O(N355));

  xor2  gate511(.a(N308), .b(N343), .O(gate125inter0));
  nand2 gate512(.a(gate125inter0), .b(s_50), .O(gate125inter1));
  and2  gate513(.a(N308), .b(N343), .O(gate125inter2));
  inv1  gate514(.a(s_50), .O(gate125inter3));
  inv1  gate515(.a(s_51), .O(gate125inter4));
  nand2 gate516(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate517(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate518(.a(N343), .O(gate125inter7));
  inv1  gate519(.a(N308), .O(gate125inter8));
  nand2 gate520(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate521(.a(s_51), .b(gate125inter3), .O(gate125inter10));
  nor2  gate522(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate523(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate524(.a(gate125inter12), .b(gate125inter1), .O(N356));
and9 gate126( .a(N348), .b(N349), .c(N350), .d(N351), .e(N352), .f(N353), .g(N354), .h(N355), .i(N356), .O(N357) );
inv1 gate127( .a(N357), .O(N360) );
inv1 gate128( .a(N357), .O(N370) );
nand2 gate129( .a(N14), .b(N360), .O(N371) );

  xor2  gate203(.a(N27), .b(N360), .O(gate130inter0));
  nand2 gate204(.a(gate130inter0), .b(s_6), .O(gate130inter1));
  and2  gate205(.a(N27), .b(N360), .O(gate130inter2));
  inv1  gate206(.a(s_6), .O(gate130inter3));
  inv1  gate207(.a(s_7), .O(gate130inter4));
  nand2 gate208(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate209(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate210(.a(N360), .O(gate130inter7));
  inv1  gate211(.a(N27), .O(gate130inter8));
  nand2 gate212(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate213(.a(s_7), .b(gate130inter3), .O(gate130inter10));
  nor2  gate214(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate215(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate216(.a(gate130inter12), .b(gate130inter1), .O(N372));
nand2 gate131( .a(N360), .b(N40), .O(N373) );
nand2 gate132( .a(N360), .b(N53), .O(N374) );
nand2 gate133( .a(N360), .b(N66), .O(N375) );

  xor2  gate161(.a(N79), .b(N360), .O(gate134inter0));
  nand2 gate162(.a(gate134inter0), .b(s_0), .O(gate134inter1));
  and2  gate163(.a(N79), .b(N360), .O(gate134inter2));
  inv1  gate164(.a(s_0), .O(gate134inter3));
  inv1  gate165(.a(s_1), .O(gate134inter4));
  nand2 gate166(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate167(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate168(.a(N360), .O(gate134inter7));
  inv1  gate169(.a(N79), .O(gate134inter8));
  nand2 gate170(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate171(.a(s_1), .b(gate134inter3), .O(gate134inter10));
  nor2  gate172(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate173(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate174(.a(gate134inter12), .b(gate134inter1), .O(N376));
nand2 gate135( .a(N360), .b(N92), .O(N377) );

  xor2  gate259(.a(N105), .b(N360), .O(gate136inter0));
  nand2 gate260(.a(gate136inter0), .b(s_14), .O(gate136inter1));
  and2  gate261(.a(N105), .b(N360), .O(gate136inter2));
  inv1  gate262(.a(s_14), .O(gate136inter3));
  inv1  gate263(.a(s_15), .O(gate136inter4));
  nand2 gate264(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate265(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate266(.a(N360), .O(gate136inter7));
  inv1  gate267(.a(N105), .O(gate136inter8));
  nand2 gate268(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate269(.a(s_15), .b(gate136inter3), .O(gate136inter10));
  nor2  gate270(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate271(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate272(.a(gate136inter12), .b(gate136inter1), .O(N378));
nand2 gate137( .a(N360), .b(N115), .O(N379) );
nand4 gate138( .a(N4), .b(N242), .c(N334), .d(N371), .O(N380) );
nand4 gate139( .a(N246), .b(N336), .c(N372), .d(N17), .O(N381) );
nand4 gate140( .a(N250), .b(N338), .c(N373), .d(N30), .O(N386) );
nand4 gate141( .a(N254), .b(N340), .c(N374), .d(N43), .O(N393) );
nand4 gate142( .a(N255), .b(N342), .c(N375), .d(N56), .O(N399) );
nand4 gate143( .a(N256), .b(N344), .c(N376), .d(N69), .O(N404) );
nand4 gate144( .a(N257), .b(N345), .c(N377), .d(N82), .O(N407) );
nand4 gate145( .a(N258), .b(N346), .c(N378), .d(N95), .O(N411) );
nand4 gate146( .a(N259), .b(N347), .c(N379), .d(N108), .O(N414) );
inv1 gate147( .a(N380), .O(N415) );
and8 gate148( .a(N381), .b(N386), .c(N393), .d(N399), .e(N404), .f(N407), .g(N411), .h(N414), .O(N416) );
inv1 gate149( .a(N393), .O(N417) );
inv1 gate150( .a(N404), .O(N418) );
inv1 gate151( .a(N407), .O(N419) );
inv1 gate152( .a(N411), .O(N420) );
nor2 gate153( .a(N415), .b(N416), .O(N421) );
nand2 gate154( .a(N386), .b(N417), .O(N422) );
nand4 gate155( .a(N386), .b(N393), .c(N418), .d(N399), .O(N425) );
nand3 gate156( .a(N399), .b(N393), .c(N419), .O(N428) );
nand4 gate157( .a(N386), .b(N393), .c(N407), .d(N420), .O(N429) );
nand4 gate158( .a(N381), .b(N386), .c(N422), .d(N399), .O(N430) );
nand4 gate159( .a(N381), .b(N386), .c(N425), .d(N428), .O(N431) );
nand4 gate160( .a(N381), .b(N422), .c(N425), .d(N429), .O(N432) );

endmodule