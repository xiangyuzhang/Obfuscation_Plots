module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate841(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate842(.a(gate15inter0), .b(s_42), .O(gate15inter1));
  and2  gate843(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate844(.a(s_42), .O(gate15inter3));
  inv1  gate845(.a(s_43), .O(gate15inter4));
  nand2 gate846(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate847(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate848(.a(G13), .O(gate15inter7));
  inv1  gate849(.a(G14), .O(gate15inter8));
  nand2 gate850(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate851(.a(s_43), .b(gate15inter3), .O(gate15inter10));
  nor2  gate852(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate853(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate854(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate1023(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate1024(.a(gate21inter0), .b(s_68), .O(gate21inter1));
  and2  gate1025(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate1026(.a(s_68), .O(gate21inter3));
  inv1  gate1027(.a(s_69), .O(gate21inter4));
  nand2 gate1028(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate1029(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate1030(.a(G25), .O(gate21inter7));
  inv1  gate1031(.a(G26), .O(gate21inter8));
  nand2 gate1032(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate1033(.a(s_69), .b(gate21inter3), .O(gate21inter10));
  nor2  gate1034(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate1035(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate1036(.a(gate21inter12), .b(gate21inter1), .O(G302));

  xor2  gate897(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate898(.a(gate22inter0), .b(s_50), .O(gate22inter1));
  and2  gate899(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate900(.a(s_50), .O(gate22inter3));
  inv1  gate901(.a(s_51), .O(gate22inter4));
  nand2 gate902(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate903(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate904(.a(G27), .O(gate22inter7));
  inv1  gate905(.a(G28), .O(gate22inter8));
  nand2 gate906(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate907(.a(s_51), .b(gate22inter3), .O(gate22inter10));
  nor2  gate908(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate909(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate910(.a(gate22inter12), .b(gate22inter1), .O(G305));
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate1317(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate1318(.a(gate27inter0), .b(s_110), .O(gate27inter1));
  and2  gate1319(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate1320(.a(s_110), .O(gate27inter3));
  inv1  gate1321(.a(s_111), .O(gate27inter4));
  nand2 gate1322(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate1323(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate1324(.a(G2), .O(gate27inter7));
  inv1  gate1325(.a(G6), .O(gate27inter8));
  nand2 gate1326(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate1327(.a(s_111), .b(gate27inter3), .O(gate27inter10));
  nor2  gate1328(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate1329(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate1330(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate981(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate982(.a(gate29inter0), .b(s_62), .O(gate29inter1));
  and2  gate983(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate984(.a(s_62), .O(gate29inter3));
  inv1  gate985(.a(s_63), .O(gate29inter4));
  nand2 gate986(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate987(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate988(.a(G3), .O(gate29inter7));
  inv1  gate989(.a(G7), .O(gate29inter8));
  nand2 gate990(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate991(.a(s_63), .b(gate29inter3), .O(gate29inter10));
  nor2  gate992(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate993(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate994(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate785(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate786(.a(gate33inter0), .b(s_34), .O(gate33inter1));
  and2  gate787(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate788(.a(s_34), .O(gate33inter3));
  inv1  gate789(.a(s_35), .O(gate33inter4));
  nand2 gate790(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate791(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate792(.a(G17), .O(gate33inter7));
  inv1  gate793(.a(G21), .O(gate33inter8));
  nand2 gate794(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate795(.a(s_35), .b(gate33inter3), .O(gate33inter10));
  nor2  gate796(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate797(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate798(.a(gate33inter12), .b(gate33inter1), .O(G338));
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate1191(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate1192(.a(gate37inter0), .b(s_92), .O(gate37inter1));
  and2  gate1193(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate1194(.a(s_92), .O(gate37inter3));
  inv1  gate1195(.a(s_93), .O(gate37inter4));
  nand2 gate1196(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate1197(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate1198(.a(G19), .O(gate37inter7));
  inv1  gate1199(.a(G23), .O(gate37inter8));
  nand2 gate1200(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate1201(.a(s_93), .b(gate37inter3), .O(gate37inter10));
  nor2  gate1202(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate1203(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate1204(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate1051(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate1052(.a(gate44inter0), .b(s_72), .O(gate44inter1));
  and2  gate1053(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate1054(.a(s_72), .O(gate44inter3));
  inv1  gate1055(.a(s_73), .O(gate44inter4));
  nand2 gate1056(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate1057(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate1058(.a(G4), .O(gate44inter7));
  inv1  gate1059(.a(G269), .O(gate44inter8));
  nand2 gate1060(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate1061(.a(s_73), .b(gate44inter3), .O(gate44inter10));
  nor2  gate1062(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate1063(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate1064(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate645(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate646(.a(gate71inter0), .b(s_14), .O(gate71inter1));
  and2  gate647(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate648(.a(s_14), .O(gate71inter3));
  inv1  gate649(.a(s_15), .O(gate71inter4));
  nand2 gate650(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate651(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate652(.a(G31), .O(gate71inter7));
  inv1  gate653(.a(G311), .O(gate71inter8));
  nand2 gate654(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate655(.a(s_15), .b(gate71inter3), .O(gate71inter10));
  nor2  gate656(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate657(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate658(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );

  xor2  gate911(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate912(.a(gate76inter0), .b(s_52), .O(gate76inter1));
  and2  gate913(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate914(.a(s_52), .O(gate76inter3));
  inv1  gate915(.a(s_53), .O(gate76inter4));
  nand2 gate916(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate917(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate918(.a(G13), .O(gate76inter7));
  inv1  gate919(.a(G317), .O(gate76inter8));
  nand2 gate920(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate921(.a(s_53), .b(gate76inter3), .O(gate76inter10));
  nor2  gate922(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate923(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate924(.a(gate76inter12), .b(gate76inter1), .O(G397));

  xor2  gate771(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate772(.a(gate77inter0), .b(s_32), .O(gate77inter1));
  and2  gate773(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate774(.a(s_32), .O(gate77inter3));
  inv1  gate775(.a(s_33), .O(gate77inter4));
  nand2 gate776(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate777(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate778(.a(G2), .O(gate77inter7));
  inv1  gate779(.a(G320), .O(gate77inter8));
  nand2 gate780(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate781(.a(s_33), .b(gate77inter3), .O(gate77inter10));
  nor2  gate782(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate783(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate784(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate1205(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate1206(.a(gate82inter0), .b(s_94), .O(gate82inter1));
  and2  gate1207(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate1208(.a(s_94), .O(gate82inter3));
  inv1  gate1209(.a(s_95), .O(gate82inter4));
  nand2 gate1210(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate1211(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate1212(.a(G7), .O(gate82inter7));
  inv1  gate1213(.a(G326), .O(gate82inter8));
  nand2 gate1214(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate1215(.a(s_95), .b(gate82inter3), .O(gate82inter10));
  nor2  gate1216(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate1217(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate1218(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate687(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate688(.a(gate85inter0), .b(s_20), .O(gate85inter1));
  and2  gate689(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate690(.a(s_20), .O(gate85inter3));
  inv1  gate691(.a(s_21), .O(gate85inter4));
  nand2 gate692(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate693(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate694(.a(G4), .O(gate85inter7));
  inv1  gate695(.a(G332), .O(gate85inter8));
  nand2 gate696(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate697(.a(s_21), .b(gate85inter3), .O(gate85inter10));
  nor2  gate698(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate699(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate700(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate1149(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate1150(.a(gate88inter0), .b(s_86), .O(gate88inter1));
  and2  gate1151(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate1152(.a(s_86), .O(gate88inter3));
  inv1  gate1153(.a(s_87), .O(gate88inter4));
  nand2 gate1154(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate1155(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate1156(.a(G16), .O(gate88inter7));
  inv1  gate1157(.a(G335), .O(gate88inter8));
  nand2 gate1158(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate1159(.a(s_87), .b(gate88inter3), .O(gate88inter10));
  nor2  gate1160(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate1161(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate1162(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate603(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate604(.a(gate91inter0), .b(s_8), .O(gate91inter1));
  and2  gate605(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate606(.a(s_8), .O(gate91inter3));
  inv1  gate607(.a(s_9), .O(gate91inter4));
  nand2 gate608(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate609(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate610(.a(G25), .O(gate91inter7));
  inv1  gate611(.a(G341), .O(gate91inter8));
  nand2 gate612(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate613(.a(s_9), .b(gate91inter3), .O(gate91inter10));
  nor2  gate614(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate615(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate616(.a(gate91inter12), .b(gate91inter1), .O(G412));

  xor2  gate1079(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate1080(.a(gate92inter0), .b(s_76), .O(gate92inter1));
  and2  gate1081(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate1082(.a(s_76), .O(gate92inter3));
  inv1  gate1083(.a(s_77), .O(gate92inter4));
  nand2 gate1084(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate1085(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate1086(.a(G29), .O(gate92inter7));
  inv1  gate1087(.a(G341), .O(gate92inter8));
  nand2 gate1088(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate1089(.a(s_77), .b(gate92inter3), .O(gate92inter10));
  nor2  gate1090(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate1091(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate1092(.a(gate92inter12), .b(gate92inter1), .O(G413));

  xor2  gate1135(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate1136(.a(gate93inter0), .b(s_84), .O(gate93inter1));
  and2  gate1137(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate1138(.a(s_84), .O(gate93inter3));
  inv1  gate1139(.a(s_85), .O(gate93inter4));
  nand2 gate1140(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate1141(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate1142(.a(G18), .O(gate93inter7));
  inv1  gate1143(.a(G344), .O(gate93inter8));
  nand2 gate1144(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate1145(.a(s_85), .b(gate93inter3), .O(gate93inter10));
  nor2  gate1146(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate1147(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate1148(.a(gate93inter12), .b(gate93inter1), .O(G414));
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate757(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate758(.a(gate106inter0), .b(s_30), .O(gate106inter1));
  and2  gate759(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate760(.a(s_30), .O(gate106inter3));
  inv1  gate761(.a(s_31), .O(gate106inter4));
  nand2 gate762(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate763(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate764(.a(G364), .O(gate106inter7));
  inv1  gate765(.a(G365), .O(gate106inter8));
  nand2 gate766(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate767(.a(s_31), .b(gate106inter3), .O(gate106inter10));
  nor2  gate768(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate769(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate770(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );

  xor2  gate1121(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate1122(.a(gate134inter0), .b(s_82), .O(gate134inter1));
  and2  gate1123(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate1124(.a(s_82), .O(gate134inter3));
  inv1  gate1125(.a(s_83), .O(gate134inter4));
  nand2 gate1126(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate1127(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate1128(.a(G420), .O(gate134inter7));
  inv1  gate1129(.a(G421), .O(gate134inter8));
  nand2 gate1130(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate1131(.a(s_83), .b(gate134inter3), .O(gate134inter10));
  nor2  gate1132(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate1133(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate1134(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );

  xor2  gate855(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate856(.a(gate139inter0), .b(s_44), .O(gate139inter1));
  and2  gate857(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate858(.a(s_44), .O(gate139inter3));
  inv1  gate859(.a(s_45), .O(gate139inter4));
  nand2 gate860(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate861(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate862(.a(G438), .O(gate139inter7));
  inv1  gate863(.a(G441), .O(gate139inter8));
  nand2 gate864(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate865(.a(s_45), .b(gate139inter3), .O(gate139inter10));
  nor2  gate866(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate867(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate868(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate1065(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1066(.a(gate148inter0), .b(s_74), .O(gate148inter1));
  and2  gate1067(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1068(.a(s_74), .O(gate148inter3));
  inv1  gate1069(.a(s_75), .O(gate148inter4));
  nand2 gate1070(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1071(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1072(.a(G492), .O(gate148inter7));
  inv1  gate1073(.a(G495), .O(gate148inter8));
  nand2 gate1074(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1075(.a(s_75), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1076(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1077(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1078(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );

  xor2  gate673(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate674(.a(gate152inter0), .b(s_18), .O(gate152inter1));
  and2  gate675(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate676(.a(s_18), .O(gate152inter3));
  inv1  gate677(.a(s_19), .O(gate152inter4));
  nand2 gate678(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate679(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate680(.a(G516), .O(gate152inter7));
  inv1  gate681(.a(G519), .O(gate152inter8));
  nand2 gate682(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate683(.a(s_19), .b(gate152inter3), .O(gate152inter10));
  nor2  gate684(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate685(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate686(.a(gate152inter12), .b(gate152inter1), .O(G567));

  xor2  gate561(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate562(.a(gate153inter0), .b(s_2), .O(gate153inter1));
  and2  gate563(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate564(.a(s_2), .O(gate153inter3));
  inv1  gate565(.a(s_3), .O(gate153inter4));
  nand2 gate566(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate567(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate568(.a(G426), .O(gate153inter7));
  inv1  gate569(.a(G522), .O(gate153inter8));
  nand2 gate570(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate571(.a(s_3), .b(gate153inter3), .O(gate153inter10));
  nor2  gate572(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate573(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate574(.a(gate153inter12), .b(gate153inter1), .O(G570));
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate547(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate548(.a(gate161inter0), .b(s_0), .O(gate161inter1));
  and2  gate549(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate550(.a(s_0), .O(gate161inter3));
  inv1  gate551(.a(s_1), .O(gate161inter4));
  nand2 gate552(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate553(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate554(.a(G450), .O(gate161inter7));
  inv1  gate555(.a(G534), .O(gate161inter8));
  nand2 gate556(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate557(.a(s_1), .b(gate161inter3), .O(gate161inter10));
  nor2  gate558(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate559(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate560(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );

  xor2  gate729(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate730(.a(gate163inter0), .b(s_26), .O(gate163inter1));
  and2  gate731(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate732(.a(s_26), .O(gate163inter3));
  inv1  gate733(.a(s_27), .O(gate163inter4));
  nand2 gate734(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate735(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate736(.a(G456), .O(gate163inter7));
  inv1  gate737(.a(G537), .O(gate163inter8));
  nand2 gate738(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate739(.a(s_27), .b(gate163inter3), .O(gate163inter10));
  nor2  gate740(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate741(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate742(.a(gate163inter12), .b(gate163inter1), .O(G580));
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );

  xor2  gate1261(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate1262(.a(gate168inter0), .b(s_102), .O(gate168inter1));
  and2  gate1263(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate1264(.a(s_102), .O(gate168inter3));
  inv1  gate1265(.a(s_103), .O(gate168inter4));
  nand2 gate1266(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate1267(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate1268(.a(G471), .O(gate168inter7));
  inv1  gate1269(.a(G543), .O(gate168inter8));
  nand2 gate1270(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate1271(.a(s_103), .b(gate168inter3), .O(gate168inter10));
  nor2  gate1272(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate1273(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate1274(.a(gate168inter12), .b(gate168inter1), .O(G585));
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate827(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate828(.a(gate170inter0), .b(s_40), .O(gate170inter1));
  and2  gate829(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate830(.a(s_40), .O(gate170inter3));
  inv1  gate831(.a(s_41), .O(gate170inter4));
  nand2 gate832(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate833(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate834(.a(G477), .O(gate170inter7));
  inv1  gate835(.a(G546), .O(gate170inter8));
  nand2 gate836(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate837(.a(s_41), .b(gate170inter3), .O(gate170inter10));
  nor2  gate838(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate839(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate840(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate1247(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate1248(.a(gate174inter0), .b(s_100), .O(gate174inter1));
  and2  gate1249(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate1250(.a(s_100), .O(gate174inter3));
  inv1  gate1251(.a(s_101), .O(gate174inter4));
  nand2 gate1252(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate1253(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate1254(.a(G489), .O(gate174inter7));
  inv1  gate1255(.a(G552), .O(gate174inter8));
  nand2 gate1256(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate1257(.a(s_101), .b(gate174inter3), .O(gate174inter10));
  nor2  gate1258(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate1259(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate1260(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );

  xor2  gate617(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate618(.a(gate189inter0), .b(s_10), .O(gate189inter1));
  and2  gate619(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate620(.a(s_10), .O(gate189inter3));
  inv1  gate621(.a(s_11), .O(gate189inter4));
  nand2 gate622(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate623(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate624(.a(G578), .O(gate189inter7));
  inv1  gate625(.a(G579), .O(gate189inter8));
  nand2 gate626(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate627(.a(s_11), .b(gate189inter3), .O(gate189inter10));
  nor2  gate628(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate629(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate630(.a(gate189inter12), .b(gate189inter1), .O(G622));
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate1093(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate1094(.a(gate200inter0), .b(s_78), .O(gate200inter1));
  and2  gate1095(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate1096(.a(s_78), .O(gate200inter3));
  inv1  gate1097(.a(s_79), .O(gate200inter4));
  nand2 gate1098(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate1099(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate1100(.a(G600), .O(gate200inter7));
  inv1  gate1101(.a(G601), .O(gate200inter8));
  nand2 gate1102(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate1103(.a(s_79), .b(gate200inter3), .O(gate200inter10));
  nor2  gate1104(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate1105(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate1106(.a(gate200inter12), .b(gate200inter1), .O(G663));

  xor2  gate939(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate940(.a(gate201inter0), .b(s_56), .O(gate201inter1));
  and2  gate941(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate942(.a(s_56), .O(gate201inter3));
  inv1  gate943(.a(s_57), .O(gate201inter4));
  nand2 gate944(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate945(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate946(.a(G602), .O(gate201inter7));
  inv1  gate947(.a(G607), .O(gate201inter8));
  nand2 gate948(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate949(.a(s_57), .b(gate201inter3), .O(gate201inter10));
  nor2  gate950(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate951(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate952(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate1107(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate1108(.a(gate206inter0), .b(s_80), .O(gate206inter1));
  and2  gate1109(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate1110(.a(s_80), .O(gate206inter3));
  inv1  gate1111(.a(s_81), .O(gate206inter4));
  nand2 gate1112(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate1113(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate1114(.a(G632), .O(gate206inter7));
  inv1  gate1115(.a(G637), .O(gate206inter8));
  nand2 gate1116(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate1117(.a(s_81), .b(gate206inter3), .O(gate206inter10));
  nor2  gate1118(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate1119(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate1120(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );

  xor2  gate967(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate968(.a(gate208inter0), .b(s_60), .O(gate208inter1));
  and2  gate969(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate970(.a(s_60), .O(gate208inter3));
  inv1  gate971(.a(s_61), .O(gate208inter4));
  nand2 gate972(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate973(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate974(.a(G627), .O(gate208inter7));
  inv1  gate975(.a(G637), .O(gate208inter8));
  nand2 gate976(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate977(.a(s_61), .b(gate208inter3), .O(gate208inter10));
  nor2  gate978(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate979(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate980(.a(gate208inter12), .b(gate208inter1), .O(G687));
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate1303(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate1304(.a(gate211inter0), .b(s_108), .O(gate211inter1));
  and2  gate1305(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate1306(.a(s_108), .O(gate211inter3));
  inv1  gate1307(.a(s_109), .O(gate211inter4));
  nand2 gate1308(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate1309(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate1310(.a(G612), .O(gate211inter7));
  inv1  gate1311(.a(G669), .O(gate211inter8));
  nand2 gate1312(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate1313(.a(s_109), .b(gate211inter3), .O(gate211inter10));
  nor2  gate1314(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate1315(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate1316(.a(gate211inter12), .b(gate211inter1), .O(G692));

  xor2  gate1009(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate1010(.a(gate212inter0), .b(s_66), .O(gate212inter1));
  and2  gate1011(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate1012(.a(s_66), .O(gate212inter3));
  inv1  gate1013(.a(s_67), .O(gate212inter4));
  nand2 gate1014(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate1015(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate1016(.a(G617), .O(gate212inter7));
  inv1  gate1017(.a(G669), .O(gate212inter8));
  nand2 gate1018(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate1019(.a(s_67), .b(gate212inter3), .O(gate212inter10));
  nor2  gate1020(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate1021(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate1022(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate995(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate996(.a(gate231inter0), .b(s_64), .O(gate231inter1));
  and2  gate997(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate998(.a(s_64), .O(gate231inter3));
  inv1  gate999(.a(s_65), .O(gate231inter4));
  nand2 gate1000(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate1001(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate1002(.a(G702), .O(gate231inter7));
  inv1  gate1003(.a(G703), .O(gate231inter8));
  nand2 gate1004(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate1005(.a(s_65), .b(gate231inter3), .O(gate231inter10));
  nor2  gate1006(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate1007(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate1008(.a(gate231inter12), .b(gate231inter1), .O(G724));

  xor2  gate1177(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate1178(.a(gate232inter0), .b(s_90), .O(gate232inter1));
  and2  gate1179(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate1180(.a(s_90), .O(gate232inter3));
  inv1  gate1181(.a(s_91), .O(gate232inter4));
  nand2 gate1182(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate1183(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate1184(.a(G704), .O(gate232inter7));
  inv1  gate1185(.a(G705), .O(gate232inter8));
  nand2 gate1186(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate1187(.a(s_91), .b(gate232inter3), .O(gate232inter10));
  nor2  gate1188(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate1189(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate1190(.a(gate232inter12), .b(gate232inter1), .O(G727));
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate1275(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate1276(.a(gate248inter0), .b(s_104), .O(gate248inter1));
  and2  gate1277(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate1278(.a(s_104), .O(gate248inter3));
  inv1  gate1279(.a(s_105), .O(gate248inter4));
  nand2 gate1280(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate1281(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate1282(.a(G727), .O(gate248inter7));
  inv1  gate1283(.a(G739), .O(gate248inter8));
  nand2 gate1284(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate1285(.a(s_105), .b(gate248inter3), .O(gate248inter10));
  nor2  gate1286(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate1287(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate1288(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate1037(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate1038(.a(gate252inter0), .b(s_70), .O(gate252inter1));
  and2  gate1039(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate1040(.a(s_70), .O(gate252inter3));
  inv1  gate1041(.a(s_71), .O(gate252inter4));
  nand2 gate1042(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate1043(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate1044(.a(G709), .O(gate252inter7));
  inv1  gate1045(.a(G745), .O(gate252inter8));
  nand2 gate1046(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate1047(.a(s_71), .b(gate252inter3), .O(gate252inter10));
  nor2  gate1048(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate1049(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate1050(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate715(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate716(.a(gate256inter0), .b(s_24), .O(gate256inter1));
  and2  gate717(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate718(.a(s_24), .O(gate256inter3));
  inv1  gate719(.a(s_25), .O(gate256inter4));
  nand2 gate720(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate721(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate722(.a(G715), .O(gate256inter7));
  inv1  gate723(.a(G751), .O(gate256inter8));
  nand2 gate724(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate725(.a(s_25), .b(gate256inter3), .O(gate256inter10));
  nor2  gate726(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate727(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate728(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate743(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate744(.a(gate269inter0), .b(s_28), .O(gate269inter1));
  and2  gate745(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate746(.a(s_28), .O(gate269inter3));
  inv1  gate747(.a(s_29), .O(gate269inter4));
  nand2 gate748(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate749(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate750(.a(G654), .O(gate269inter7));
  inv1  gate751(.a(G782), .O(gate269inter8));
  nand2 gate752(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate753(.a(s_29), .b(gate269inter3), .O(gate269inter10));
  nor2  gate754(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate755(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate756(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate869(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate870(.a(gate272inter0), .b(s_46), .O(gate272inter1));
  and2  gate871(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate872(.a(s_46), .O(gate272inter3));
  inv1  gate873(.a(s_47), .O(gate272inter4));
  nand2 gate874(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate875(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate876(.a(G663), .O(gate272inter7));
  inv1  gate877(.a(G791), .O(gate272inter8));
  nand2 gate878(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate879(.a(s_47), .b(gate272inter3), .O(gate272inter10));
  nor2  gate880(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate881(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate882(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate1163(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate1164(.a(gate274inter0), .b(s_88), .O(gate274inter1));
  and2  gate1165(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate1166(.a(s_88), .O(gate274inter3));
  inv1  gate1167(.a(s_89), .O(gate274inter4));
  nand2 gate1168(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate1169(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate1170(.a(G770), .O(gate274inter7));
  inv1  gate1171(.a(G794), .O(gate274inter8));
  nand2 gate1172(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate1173(.a(s_89), .b(gate274inter3), .O(gate274inter10));
  nor2  gate1174(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate1175(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate1176(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate701(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate702(.a(gate279inter0), .b(s_22), .O(gate279inter1));
  and2  gate703(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate704(.a(s_22), .O(gate279inter3));
  inv1  gate705(.a(s_23), .O(gate279inter4));
  nand2 gate706(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate707(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate708(.a(G651), .O(gate279inter7));
  inv1  gate709(.a(G803), .O(gate279inter8));
  nand2 gate710(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate711(.a(s_23), .b(gate279inter3), .O(gate279inter10));
  nor2  gate712(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate713(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate714(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate589(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate590(.a(gate296inter0), .b(s_6), .O(gate296inter1));
  and2  gate591(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate592(.a(s_6), .O(gate296inter3));
  inv1  gate593(.a(s_7), .O(gate296inter4));
  nand2 gate594(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate595(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate596(.a(G826), .O(gate296inter7));
  inv1  gate597(.a(G827), .O(gate296inter8));
  nand2 gate598(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate599(.a(s_7), .b(gate296inter3), .O(gate296inter10));
  nor2  gate600(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate601(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate602(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate659(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate660(.a(gate390inter0), .b(s_16), .O(gate390inter1));
  and2  gate661(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate662(.a(s_16), .O(gate390inter3));
  inv1  gate663(.a(s_17), .O(gate390inter4));
  nand2 gate664(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate665(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate666(.a(G4), .O(gate390inter7));
  inv1  gate667(.a(G1045), .O(gate390inter8));
  nand2 gate668(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate669(.a(s_17), .b(gate390inter3), .O(gate390inter10));
  nor2  gate670(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate671(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate672(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );

  xor2  gate813(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate814(.a(gate396inter0), .b(s_38), .O(gate396inter1));
  and2  gate815(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate816(.a(s_38), .O(gate396inter3));
  inv1  gate817(.a(s_39), .O(gate396inter4));
  nand2 gate818(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate819(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate820(.a(G10), .O(gate396inter7));
  inv1  gate821(.a(G1063), .O(gate396inter8));
  nand2 gate822(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate823(.a(s_39), .b(gate396inter3), .O(gate396inter10));
  nor2  gate824(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate825(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate826(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate1233(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1234(.a(gate420inter0), .b(s_98), .O(gate420inter1));
  and2  gate1235(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1236(.a(s_98), .O(gate420inter3));
  inv1  gate1237(.a(s_99), .O(gate420inter4));
  nand2 gate1238(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1239(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1240(.a(G1036), .O(gate420inter7));
  inv1  gate1241(.a(G1132), .O(gate420inter8));
  nand2 gate1242(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1243(.a(s_99), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1244(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1245(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1246(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );

  xor2  gate925(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate926(.a(gate423inter0), .b(s_54), .O(gate423inter1));
  and2  gate927(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate928(.a(s_54), .O(gate423inter3));
  inv1  gate929(.a(s_55), .O(gate423inter4));
  nand2 gate930(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate931(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate932(.a(G3), .O(gate423inter7));
  inv1  gate933(.a(G1138), .O(gate423inter8));
  nand2 gate934(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate935(.a(s_55), .b(gate423inter3), .O(gate423inter10));
  nor2  gate936(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate937(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate938(.a(gate423inter12), .b(gate423inter1), .O(G1232));
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate575(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate576(.a(gate430inter0), .b(s_4), .O(gate430inter1));
  and2  gate577(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate578(.a(s_4), .O(gate430inter3));
  inv1  gate579(.a(s_5), .O(gate430inter4));
  nand2 gate580(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate581(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate582(.a(G1051), .O(gate430inter7));
  inv1  gate583(.a(G1147), .O(gate430inter8));
  nand2 gate584(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate585(.a(s_5), .b(gate430inter3), .O(gate430inter10));
  nor2  gate586(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate587(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate588(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate953(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate954(.a(gate441inter0), .b(s_58), .O(gate441inter1));
  and2  gate955(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate956(.a(s_58), .O(gate441inter3));
  inv1  gate957(.a(s_59), .O(gate441inter4));
  nand2 gate958(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate959(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate960(.a(G12), .O(gate441inter7));
  inv1  gate961(.a(G1165), .O(gate441inter8));
  nand2 gate962(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate963(.a(s_59), .b(gate441inter3), .O(gate441inter10));
  nor2  gate964(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate965(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate966(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate631(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate632(.a(gate443inter0), .b(s_12), .O(gate443inter1));
  and2  gate633(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate634(.a(s_12), .O(gate443inter3));
  inv1  gate635(.a(s_13), .O(gate443inter4));
  nand2 gate636(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate637(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate638(.a(G13), .O(gate443inter7));
  inv1  gate639(.a(G1168), .O(gate443inter8));
  nand2 gate640(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate641(.a(s_13), .b(gate443inter3), .O(gate443inter10));
  nor2  gate642(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate643(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate644(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate883(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate884(.a(gate465inter0), .b(s_48), .O(gate465inter1));
  and2  gate885(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate886(.a(s_48), .O(gate465inter3));
  inv1  gate887(.a(s_49), .O(gate465inter4));
  nand2 gate888(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate889(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate890(.a(G24), .O(gate465inter7));
  inv1  gate891(.a(G1201), .O(gate465inter8));
  nand2 gate892(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate893(.a(s_49), .b(gate465inter3), .O(gate465inter10));
  nor2  gate894(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate895(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate896(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate1289(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate1290(.a(gate492inter0), .b(s_106), .O(gate492inter1));
  and2  gate1291(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate1292(.a(s_106), .O(gate492inter3));
  inv1  gate1293(.a(s_107), .O(gate492inter4));
  nand2 gate1294(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate1295(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate1296(.a(G1246), .O(gate492inter7));
  inv1  gate1297(.a(G1247), .O(gate492inter8));
  nand2 gate1298(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate1299(.a(s_107), .b(gate492inter3), .O(gate492inter10));
  nor2  gate1300(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate1301(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate1302(.a(gate492inter12), .b(gate492inter1), .O(G1301));
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );

  xor2  gate799(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate800(.a(gate495inter0), .b(s_36), .O(gate495inter1));
  and2  gate801(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate802(.a(s_36), .O(gate495inter3));
  inv1  gate803(.a(s_37), .O(gate495inter4));
  nand2 gate804(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate805(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate806(.a(G1252), .O(gate495inter7));
  inv1  gate807(.a(G1253), .O(gate495inter8));
  nand2 gate808(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate809(.a(s_37), .b(gate495inter3), .O(gate495inter10));
  nor2  gate810(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate811(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate812(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate1219(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate1220(.a(gate503inter0), .b(s_96), .O(gate503inter1));
  and2  gate1221(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate1222(.a(s_96), .O(gate503inter3));
  inv1  gate1223(.a(s_97), .O(gate503inter4));
  nand2 gate1224(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate1225(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate1226(.a(G1268), .O(gate503inter7));
  inv1  gate1227(.a(G1269), .O(gate503inter8));
  nand2 gate1228(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate1229(.a(s_97), .b(gate503inter3), .O(gate503inter10));
  nor2  gate1230(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate1231(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate1232(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule