module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );

  xor2  gate897(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate898(.a(gate10inter0), .b(s_50), .O(gate10inter1));
  and2  gate899(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate900(.a(s_50), .O(gate10inter3));
  inv1  gate901(.a(s_51), .O(gate10inter4));
  nand2 gate902(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate903(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate904(.a(G3), .O(gate10inter7));
  inv1  gate905(.a(G4), .O(gate10inter8));
  nand2 gate906(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate907(.a(s_51), .b(gate10inter3), .O(gate10inter10));
  nor2  gate908(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate909(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate910(.a(gate10inter12), .b(gate10inter1), .O(G269));

  xor2  gate799(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate800(.a(gate11inter0), .b(s_36), .O(gate11inter1));
  and2  gate801(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate802(.a(s_36), .O(gate11inter3));
  inv1  gate803(.a(s_37), .O(gate11inter4));
  nand2 gate804(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate805(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate806(.a(G5), .O(gate11inter7));
  inv1  gate807(.a(G6), .O(gate11inter8));
  nand2 gate808(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate809(.a(s_37), .b(gate11inter3), .O(gate11inter10));
  nor2  gate810(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate811(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate812(.a(gate11inter12), .b(gate11inter1), .O(G272));

  xor2  gate1485(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate1486(.a(gate12inter0), .b(s_134), .O(gate12inter1));
  and2  gate1487(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate1488(.a(s_134), .O(gate12inter3));
  inv1  gate1489(.a(s_135), .O(gate12inter4));
  nand2 gate1490(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate1491(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate1492(.a(G7), .O(gate12inter7));
  inv1  gate1493(.a(G8), .O(gate12inter8));
  nand2 gate1494(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate1495(.a(s_135), .b(gate12inter3), .O(gate12inter10));
  nor2  gate1496(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate1497(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate1498(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );

  xor2  gate1835(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate1836(.a(gate14inter0), .b(s_184), .O(gate14inter1));
  and2  gate1837(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate1838(.a(s_184), .O(gate14inter3));
  inv1  gate1839(.a(s_185), .O(gate14inter4));
  nand2 gate1840(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate1841(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate1842(.a(G11), .O(gate14inter7));
  inv1  gate1843(.a(G12), .O(gate14inter8));
  nand2 gate1844(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate1845(.a(s_185), .b(gate14inter3), .O(gate14inter10));
  nor2  gate1846(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate1847(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate1848(.a(gate14inter12), .b(gate14inter1), .O(G281));

  xor2  gate953(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate954(.a(gate15inter0), .b(s_58), .O(gate15inter1));
  and2  gate955(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate956(.a(s_58), .O(gate15inter3));
  inv1  gate957(.a(s_59), .O(gate15inter4));
  nand2 gate958(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate959(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate960(.a(G13), .O(gate15inter7));
  inv1  gate961(.a(G14), .O(gate15inter8));
  nand2 gate962(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate963(.a(s_59), .b(gate15inter3), .O(gate15inter10));
  nor2  gate964(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate965(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate966(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate743(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate744(.a(gate17inter0), .b(s_28), .O(gate17inter1));
  and2  gate745(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate746(.a(s_28), .O(gate17inter3));
  inv1  gate747(.a(s_29), .O(gate17inter4));
  nand2 gate748(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate749(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate750(.a(G17), .O(gate17inter7));
  inv1  gate751(.a(G18), .O(gate17inter8));
  nand2 gate752(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate753(.a(s_29), .b(gate17inter3), .O(gate17inter10));
  nor2  gate754(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate755(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate756(.a(gate17inter12), .b(gate17inter1), .O(G290));

  xor2  gate883(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate884(.a(gate18inter0), .b(s_48), .O(gate18inter1));
  and2  gate885(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate886(.a(s_48), .O(gate18inter3));
  inv1  gate887(.a(s_49), .O(gate18inter4));
  nand2 gate888(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate889(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate890(.a(G19), .O(gate18inter7));
  inv1  gate891(.a(G20), .O(gate18inter8));
  nand2 gate892(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate893(.a(s_49), .b(gate18inter3), .O(gate18inter10));
  nor2  gate894(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate895(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate896(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate617(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate618(.a(gate29inter0), .b(s_10), .O(gate29inter1));
  and2  gate619(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate620(.a(s_10), .O(gate29inter3));
  inv1  gate621(.a(s_11), .O(gate29inter4));
  nand2 gate622(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate623(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate624(.a(G3), .O(gate29inter7));
  inv1  gate625(.a(G7), .O(gate29inter8));
  nand2 gate626(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate627(.a(s_11), .b(gate29inter3), .O(gate29inter10));
  nor2  gate628(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate629(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate630(.a(gate29inter12), .b(gate29inter1), .O(G326));

  xor2  gate1037(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate1038(.a(gate30inter0), .b(s_70), .O(gate30inter1));
  and2  gate1039(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate1040(.a(s_70), .O(gate30inter3));
  inv1  gate1041(.a(s_71), .O(gate30inter4));
  nand2 gate1042(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate1043(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate1044(.a(G11), .O(gate30inter7));
  inv1  gate1045(.a(G15), .O(gate30inter8));
  nand2 gate1046(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate1047(.a(s_71), .b(gate30inter3), .O(gate30inter10));
  nor2  gate1048(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate1049(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate1050(.a(gate30inter12), .b(gate30inter1), .O(G329));
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate1415(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate1416(.a(gate41inter0), .b(s_124), .O(gate41inter1));
  and2  gate1417(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate1418(.a(s_124), .O(gate41inter3));
  inv1  gate1419(.a(s_125), .O(gate41inter4));
  nand2 gate1420(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate1421(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate1422(.a(G1), .O(gate41inter7));
  inv1  gate1423(.a(G266), .O(gate41inter8));
  nand2 gate1424(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate1425(.a(s_125), .b(gate41inter3), .O(gate41inter10));
  nor2  gate1426(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate1427(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate1428(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate925(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate926(.a(gate46inter0), .b(s_54), .O(gate46inter1));
  and2  gate927(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate928(.a(s_54), .O(gate46inter3));
  inv1  gate929(.a(s_55), .O(gate46inter4));
  nand2 gate930(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate931(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate932(.a(G6), .O(gate46inter7));
  inv1  gate933(.a(G272), .O(gate46inter8));
  nand2 gate934(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate935(.a(s_55), .b(gate46inter3), .O(gate46inter10));
  nor2  gate936(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate937(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate938(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );

  xor2  gate1751(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate1752(.a(gate50inter0), .b(s_172), .O(gate50inter1));
  and2  gate1753(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate1754(.a(s_172), .O(gate50inter3));
  inv1  gate1755(.a(s_173), .O(gate50inter4));
  nand2 gate1756(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate1757(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate1758(.a(G10), .O(gate50inter7));
  inv1  gate1759(.a(G278), .O(gate50inter8));
  nand2 gate1760(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate1761(.a(s_173), .b(gate50inter3), .O(gate50inter10));
  nor2  gate1762(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate1763(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate1764(.a(gate50inter12), .b(gate50inter1), .O(G371));
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );

  xor2  gate1527(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate1528(.a(gate56inter0), .b(s_140), .O(gate56inter1));
  and2  gate1529(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate1530(.a(s_140), .O(gate56inter3));
  inv1  gate1531(.a(s_141), .O(gate56inter4));
  nand2 gate1532(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate1533(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate1534(.a(G16), .O(gate56inter7));
  inv1  gate1535(.a(G287), .O(gate56inter8));
  nand2 gate1536(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate1537(.a(s_141), .b(gate56inter3), .O(gate56inter10));
  nor2  gate1538(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate1539(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate1540(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate1387(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate1388(.a(gate59inter0), .b(s_120), .O(gate59inter1));
  and2  gate1389(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate1390(.a(s_120), .O(gate59inter3));
  inv1  gate1391(.a(s_121), .O(gate59inter4));
  nand2 gate1392(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate1393(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate1394(.a(G19), .O(gate59inter7));
  inv1  gate1395(.a(G293), .O(gate59inter8));
  nand2 gate1396(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate1397(.a(s_121), .b(gate59inter3), .O(gate59inter10));
  nor2  gate1398(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate1399(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate1400(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );

  xor2  gate1317(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate1318(.a(gate61inter0), .b(s_110), .O(gate61inter1));
  and2  gate1319(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate1320(.a(s_110), .O(gate61inter3));
  inv1  gate1321(.a(s_111), .O(gate61inter4));
  nand2 gate1322(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate1323(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate1324(.a(G21), .O(gate61inter7));
  inv1  gate1325(.a(G296), .O(gate61inter8));
  nand2 gate1326(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate1327(.a(s_111), .b(gate61inter3), .O(gate61inter10));
  nor2  gate1328(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate1329(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate1330(.a(gate61inter12), .b(gate61inter1), .O(G382));
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );

  xor2  gate1625(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate1626(.a(gate68inter0), .b(s_154), .O(gate68inter1));
  and2  gate1627(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate1628(.a(s_154), .O(gate68inter3));
  inv1  gate1629(.a(s_155), .O(gate68inter4));
  nand2 gate1630(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate1631(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate1632(.a(G28), .O(gate68inter7));
  inv1  gate1633(.a(G305), .O(gate68inter8));
  nand2 gate1634(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate1635(.a(s_155), .b(gate68inter3), .O(gate68inter10));
  nor2  gate1636(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate1637(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate1638(.a(gate68inter12), .b(gate68inter1), .O(G389));

  xor2  gate575(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate576(.a(gate69inter0), .b(s_4), .O(gate69inter1));
  and2  gate577(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate578(.a(s_4), .O(gate69inter3));
  inv1  gate579(.a(s_5), .O(gate69inter4));
  nand2 gate580(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate581(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate582(.a(G29), .O(gate69inter7));
  inv1  gate583(.a(G308), .O(gate69inter8));
  nand2 gate584(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate585(.a(s_5), .b(gate69inter3), .O(gate69inter10));
  nor2  gate586(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate587(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate588(.a(gate69inter12), .b(gate69inter1), .O(G390));
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate1191(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate1192(.a(gate71inter0), .b(s_92), .O(gate71inter1));
  and2  gate1193(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate1194(.a(s_92), .O(gate71inter3));
  inv1  gate1195(.a(s_93), .O(gate71inter4));
  nand2 gate1196(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate1197(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate1198(.a(G31), .O(gate71inter7));
  inv1  gate1199(.a(G311), .O(gate71inter8));
  nand2 gate1200(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate1201(.a(s_93), .b(gate71inter3), .O(gate71inter10));
  nor2  gate1202(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate1203(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate1204(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );

  xor2  gate1597(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate1598(.a(gate79inter0), .b(s_150), .O(gate79inter1));
  and2  gate1599(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate1600(.a(s_150), .O(gate79inter3));
  inv1  gate1601(.a(s_151), .O(gate79inter4));
  nand2 gate1602(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate1603(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate1604(.a(G10), .O(gate79inter7));
  inv1  gate1605(.a(G323), .O(gate79inter8));
  nand2 gate1606(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate1607(.a(s_151), .b(gate79inter3), .O(gate79inter10));
  nor2  gate1608(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate1609(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate1610(.a(gate79inter12), .b(gate79inter1), .O(G400));
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate1919(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate1920(.a(gate85inter0), .b(s_196), .O(gate85inter1));
  and2  gate1921(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate1922(.a(s_196), .O(gate85inter3));
  inv1  gate1923(.a(s_197), .O(gate85inter4));
  nand2 gate1924(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate1925(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate1926(.a(G4), .O(gate85inter7));
  inv1  gate1927(.a(G332), .O(gate85inter8));
  nand2 gate1928(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate1929(.a(s_197), .b(gate85inter3), .O(gate85inter10));
  nor2  gate1930(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate1931(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate1932(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate1219(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate1220(.a(gate88inter0), .b(s_96), .O(gate88inter1));
  and2  gate1221(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate1222(.a(s_96), .O(gate88inter3));
  inv1  gate1223(.a(s_97), .O(gate88inter4));
  nand2 gate1224(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate1225(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate1226(.a(G16), .O(gate88inter7));
  inv1  gate1227(.a(G335), .O(gate88inter8));
  nand2 gate1228(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate1229(.a(s_97), .b(gate88inter3), .O(gate88inter10));
  nor2  gate1230(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate1231(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate1232(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );

  xor2  gate1555(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate1556(.a(gate92inter0), .b(s_144), .O(gate92inter1));
  and2  gate1557(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate1558(.a(s_144), .O(gate92inter3));
  inv1  gate1559(.a(s_145), .O(gate92inter4));
  nand2 gate1560(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate1561(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate1562(.a(G29), .O(gate92inter7));
  inv1  gate1563(.a(G341), .O(gate92inter8));
  nand2 gate1564(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate1565(.a(s_145), .b(gate92inter3), .O(gate92inter10));
  nor2  gate1566(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate1567(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate1568(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate589(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate590(.a(gate100inter0), .b(s_6), .O(gate100inter1));
  and2  gate591(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate592(.a(s_6), .O(gate100inter3));
  inv1  gate593(.a(s_7), .O(gate100inter4));
  nand2 gate594(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate595(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate596(.a(G31), .O(gate100inter7));
  inv1  gate597(.a(G353), .O(gate100inter8));
  nand2 gate598(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate599(.a(s_7), .b(gate100inter3), .O(gate100inter10));
  nor2  gate600(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate601(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate602(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );

  xor2  gate1569(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate1570(.a(gate103inter0), .b(s_146), .O(gate103inter1));
  and2  gate1571(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate1572(.a(s_146), .O(gate103inter3));
  inv1  gate1573(.a(s_147), .O(gate103inter4));
  nand2 gate1574(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate1575(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate1576(.a(G28), .O(gate103inter7));
  inv1  gate1577(.a(G359), .O(gate103inter8));
  nand2 gate1578(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate1579(.a(s_147), .b(gate103inter3), .O(gate103inter10));
  nor2  gate1580(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate1581(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate1582(.a(gate103inter12), .b(gate103inter1), .O(G424));
nand2 gate104( .a(G32), .b(G359), .O(G425) );

  xor2  gate1401(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate1402(.a(gate105inter0), .b(s_122), .O(gate105inter1));
  and2  gate1403(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate1404(.a(s_122), .O(gate105inter3));
  inv1  gate1405(.a(s_123), .O(gate105inter4));
  nand2 gate1406(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate1407(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate1408(.a(G362), .O(gate105inter7));
  inv1  gate1409(.a(G363), .O(gate105inter8));
  nand2 gate1410(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate1411(.a(s_123), .b(gate105inter3), .O(gate105inter10));
  nor2  gate1412(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate1413(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate1414(.a(gate105inter12), .b(gate105inter1), .O(G426));
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate757(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate758(.a(gate110inter0), .b(s_30), .O(gate110inter1));
  and2  gate759(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate760(.a(s_30), .O(gate110inter3));
  inv1  gate761(.a(s_31), .O(gate110inter4));
  nand2 gate762(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate763(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate764(.a(G372), .O(gate110inter7));
  inv1  gate765(.a(G373), .O(gate110inter8));
  nand2 gate766(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate767(.a(s_31), .b(gate110inter3), .O(gate110inter10));
  nor2  gate768(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate769(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate770(.a(gate110inter12), .b(gate110inter1), .O(G441));

  xor2  gate1807(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate1808(.a(gate111inter0), .b(s_180), .O(gate111inter1));
  and2  gate1809(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate1810(.a(s_180), .O(gate111inter3));
  inv1  gate1811(.a(s_181), .O(gate111inter4));
  nand2 gate1812(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate1813(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate1814(.a(G374), .O(gate111inter7));
  inv1  gate1815(.a(G375), .O(gate111inter8));
  nand2 gate1816(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate1817(.a(s_181), .b(gate111inter3), .O(gate111inter10));
  nor2  gate1818(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate1819(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate1820(.a(gate111inter12), .b(gate111inter1), .O(G444));
nand2 gate112( .a(G376), .b(G377), .O(G447) );

  xor2  gate1961(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate1962(.a(gate113inter0), .b(s_202), .O(gate113inter1));
  and2  gate1963(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate1964(.a(s_202), .O(gate113inter3));
  inv1  gate1965(.a(s_203), .O(gate113inter4));
  nand2 gate1966(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate1967(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate1968(.a(G378), .O(gate113inter7));
  inv1  gate1969(.a(G379), .O(gate113inter8));
  nand2 gate1970(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate1971(.a(s_203), .b(gate113inter3), .O(gate113inter10));
  nor2  gate1972(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate1973(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate1974(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );

  xor2  gate1289(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate1290(.a(gate122inter0), .b(s_106), .O(gate122inter1));
  and2  gate1291(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate1292(.a(s_106), .O(gate122inter3));
  inv1  gate1293(.a(s_107), .O(gate122inter4));
  nand2 gate1294(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate1295(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate1296(.a(G396), .O(gate122inter7));
  inv1  gate1297(.a(G397), .O(gate122inter8));
  nand2 gate1298(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate1299(.a(s_107), .b(gate122inter3), .O(gate122inter10));
  nor2  gate1300(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate1301(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate1302(.a(gate122inter12), .b(gate122inter1), .O(G477));

  xor2  gate1765(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate1766(.a(gate123inter0), .b(s_174), .O(gate123inter1));
  and2  gate1767(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate1768(.a(s_174), .O(gate123inter3));
  inv1  gate1769(.a(s_175), .O(gate123inter4));
  nand2 gate1770(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate1771(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate1772(.a(G398), .O(gate123inter7));
  inv1  gate1773(.a(G399), .O(gate123inter8));
  nand2 gate1774(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate1775(.a(s_175), .b(gate123inter3), .O(gate123inter10));
  nor2  gate1776(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate1777(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate1778(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );

  xor2  gate1429(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate1430(.a(gate127inter0), .b(s_126), .O(gate127inter1));
  and2  gate1431(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate1432(.a(s_126), .O(gate127inter3));
  inv1  gate1433(.a(s_127), .O(gate127inter4));
  nand2 gate1434(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate1435(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate1436(.a(G406), .O(gate127inter7));
  inv1  gate1437(.a(G407), .O(gate127inter8));
  nand2 gate1438(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate1439(.a(s_127), .b(gate127inter3), .O(gate127inter10));
  nor2  gate1440(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate1441(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate1442(.a(gate127inter12), .b(gate127inter1), .O(G492));

  xor2  gate1275(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate1276(.a(gate128inter0), .b(s_104), .O(gate128inter1));
  and2  gate1277(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate1278(.a(s_104), .O(gate128inter3));
  inv1  gate1279(.a(s_105), .O(gate128inter4));
  nand2 gate1280(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate1281(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate1282(.a(G408), .O(gate128inter7));
  inv1  gate1283(.a(G409), .O(gate128inter8));
  nand2 gate1284(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate1285(.a(s_105), .b(gate128inter3), .O(gate128inter10));
  nor2  gate1286(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate1287(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate1288(.a(gate128inter12), .b(gate128inter1), .O(G495));
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate785(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate786(.a(gate131inter0), .b(s_34), .O(gate131inter1));
  and2  gate787(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate788(.a(s_34), .O(gate131inter3));
  inv1  gate789(.a(s_35), .O(gate131inter4));
  nand2 gate790(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate791(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate792(.a(G414), .O(gate131inter7));
  inv1  gate793(.a(G415), .O(gate131inter8));
  nand2 gate794(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate795(.a(s_35), .b(gate131inter3), .O(gate131inter10));
  nor2  gate796(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate797(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate798(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );

  xor2  gate1261(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate1262(.a(gate133inter0), .b(s_102), .O(gate133inter1));
  and2  gate1263(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate1264(.a(s_102), .O(gate133inter3));
  inv1  gate1265(.a(s_103), .O(gate133inter4));
  nand2 gate1266(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate1267(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate1268(.a(G418), .O(gate133inter7));
  inv1  gate1269(.a(G419), .O(gate133inter8));
  nand2 gate1270(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate1271(.a(s_103), .b(gate133inter3), .O(gate133inter10));
  nor2  gate1272(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate1273(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate1274(.a(gate133inter12), .b(gate133inter1), .O(G510));
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate1891(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate1892(.a(gate141inter0), .b(s_192), .O(gate141inter1));
  and2  gate1893(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate1894(.a(s_192), .O(gate141inter3));
  inv1  gate1895(.a(s_193), .O(gate141inter4));
  nand2 gate1896(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate1897(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate1898(.a(G450), .O(gate141inter7));
  inv1  gate1899(.a(G453), .O(gate141inter8));
  nand2 gate1900(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate1901(.a(s_193), .b(gate141inter3), .O(gate141inter10));
  nor2  gate1902(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate1903(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate1904(.a(gate141inter12), .b(gate141inter1), .O(G534));

  xor2  gate1513(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate1514(.a(gate142inter0), .b(s_138), .O(gate142inter1));
  and2  gate1515(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate1516(.a(s_138), .O(gate142inter3));
  inv1  gate1517(.a(s_139), .O(gate142inter4));
  nand2 gate1518(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate1519(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate1520(.a(G456), .O(gate142inter7));
  inv1  gate1521(.a(G459), .O(gate142inter8));
  nand2 gate1522(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate1523(.a(s_139), .b(gate142inter3), .O(gate142inter10));
  nor2  gate1524(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate1525(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate1526(.a(gate142inter12), .b(gate142inter1), .O(G537));
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );

  xor2  gate1023(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate1024(.a(gate163inter0), .b(s_68), .O(gate163inter1));
  and2  gate1025(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate1026(.a(s_68), .O(gate163inter3));
  inv1  gate1027(.a(s_69), .O(gate163inter4));
  nand2 gate1028(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate1029(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate1030(.a(G456), .O(gate163inter7));
  inv1  gate1031(.a(G537), .O(gate163inter8));
  nand2 gate1032(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate1033(.a(s_69), .b(gate163inter3), .O(gate163inter10));
  nor2  gate1034(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate1035(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate1036(.a(gate163inter12), .b(gate163inter1), .O(G580));

  xor2  gate2017(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate2018(.a(gate164inter0), .b(s_210), .O(gate164inter1));
  and2  gate2019(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate2020(.a(s_210), .O(gate164inter3));
  inv1  gate2021(.a(s_211), .O(gate164inter4));
  nand2 gate2022(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate2023(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate2024(.a(G459), .O(gate164inter7));
  inv1  gate2025(.a(G537), .O(gate164inter8));
  nand2 gate2026(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate2027(.a(s_211), .b(gate164inter3), .O(gate164inter10));
  nor2  gate2028(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate2029(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate2030(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate1947(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate1948(.a(gate175inter0), .b(s_200), .O(gate175inter1));
  and2  gate1949(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate1950(.a(s_200), .O(gate175inter3));
  inv1  gate1951(.a(s_201), .O(gate175inter4));
  nand2 gate1952(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1953(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1954(.a(G492), .O(gate175inter7));
  inv1  gate1955(.a(G555), .O(gate175inter8));
  nand2 gate1956(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1957(.a(s_201), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1958(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1959(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1960(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate1877(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate1878(.a(gate180inter0), .b(s_190), .O(gate180inter1));
  and2  gate1879(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate1880(.a(s_190), .O(gate180inter3));
  inv1  gate1881(.a(s_191), .O(gate180inter4));
  nand2 gate1882(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate1883(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate1884(.a(G507), .O(gate180inter7));
  inv1  gate1885(.a(G561), .O(gate180inter8));
  nand2 gate1886(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate1887(.a(s_191), .b(gate180inter3), .O(gate180inter10));
  nor2  gate1888(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate1889(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate1890(.a(gate180inter12), .b(gate180inter1), .O(G597));
nand2 gate181( .a(G510), .b(G564), .O(G598) );

  xor2  gate1975(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate1976(.a(gate182inter0), .b(s_204), .O(gate182inter1));
  and2  gate1977(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate1978(.a(s_204), .O(gate182inter3));
  inv1  gate1979(.a(s_205), .O(gate182inter4));
  nand2 gate1980(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate1981(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate1982(.a(G513), .O(gate182inter7));
  inv1  gate1983(.a(G564), .O(gate182inter8));
  nand2 gate1984(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate1985(.a(s_205), .b(gate182inter3), .O(gate182inter10));
  nor2  gate1986(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate1987(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate1988(.a(gate182inter12), .b(gate182inter1), .O(G599));

  xor2  gate1639(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate1640(.a(gate183inter0), .b(s_156), .O(gate183inter1));
  and2  gate1641(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate1642(.a(s_156), .O(gate183inter3));
  inv1  gate1643(.a(s_157), .O(gate183inter4));
  nand2 gate1644(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate1645(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate1646(.a(G516), .O(gate183inter7));
  inv1  gate1647(.a(G567), .O(gate183inter8));
  nand2 gate1648(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate1649(.a(s_157), .b(gate183inter3), .O(gate183inter10));
  nor2  gate1650(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate1651(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate1652(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate1821(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1822(.a(gate186inter0), .b(s_182), .O(gate186inter1));
  and2  gate1823(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1824(.a(s_182), .O(gate186inter3));
  inv1  gate1825(.a(s_183), .O(gate186inter4));
  nand2 gate1826(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1827(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1828(.a(G572), .O(gate186inter7));
  inv1  gate1829(.a(G573), .O(gate186inter8));
  nand2 gate1830(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1831(.a(s_183), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1832(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1833(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1834(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );

  xor2  gate1737(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate1738(.a(gate189inter0), .b(s_170), .O(gate189inter1));
  and2  gate1739(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate1740(.a(s_170), .O(gate189inter3));
  inv1  gate1741(.a(s_171), .O(gate189inter4));
  nand2 gate1742(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate1743(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate1744(.a(G578), .O(gate189inter7));
  inv1  gate1745(.a(G579), .O(gate189inter8));
  nand2 gate1746(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate1747(.a(s_171), .b(gate189inter3), .O(gate189inter10));
  nor2  gate1748(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate1749(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate1750(.a(gate189inter12), .b(gate189inter1), .O(G622));

  xor2  gate561(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate562(.a(gate190inter0), .b(s_2), .O(gate190inter1));
  and2  gate563(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate564(.a(s_2), .O(gate190inter3));
  inv1  gate565(.a(s_3), .O(gate190inter4));
  nand2 gate566(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate567(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate568(.a(G580), .O(gate190inter7));
  inv1  gate569(.a(G581), .O(gate190inter8));
  nand2 gate570(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate571(.a(s_3), .b(gate190inter3), .O(gate190inter10));
  nor2  gate572(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate573(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate574(.a(gate190inter12), .b(gate190inter1), .O(G627));
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate1541(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate1542(.a(gate196inter0), .b(s_142), .O(gate196inter1));
  and2  gate1543(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate1544(.a(s_142), .O(gate196inter3));
  inv1  gate1545(.a(s_143), .O(gate196inter4));
  nand2 gate1546(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate1547(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate1548(.a(G592), .O(gate196inter7));
  inv1  gate1549(.a(G593), .O(gate196inter8));
  nand2 gate1550(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate1551(.a(s_143), .b(gate196inter3), .O(gate196inter10));
  nor2  gate1552(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate1553(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate1554(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate855(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate856(.a(gate206inter0), .b(s_44), .O(gate206inter1));
  and2  gate857(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate858(.a(s_44), .O(gate206inter3));
  inv1  gate859(.a(s_45), .O(gate206inter4));
  nand2 gate860(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate861(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate862(.a(G632), .O(gate206inter7));
  inv1  gate863(.a(G637), .O(gate206inter8));
  nand2 gate864(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate865(.a(s_45), .b(gate206inter3), .O(gate206inter10));
  nor2  gate866(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate867(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate868(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );

  xor2  gate1093(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate1094(.a(gate209inter0), .b(s_78), .O(gate209inter1));
  and2  gate1095(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate1096(.a(s_78), .O(gate209inter3));
  inv1  gate1097(.a(s_79), .O(gate209inter4));
  nand2 gate1098(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate1099(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate1100(.a(G602), .O(gate209inter7));
  inv1  gate1101(.a(G666), .O(gate209inter8));
  nand2 gate1102(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate1103(.a(s_79), .b(gate209inter3), .O(gate209inter10));
  nor2  gate1104(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate1105(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate1106(.a(gate209inter12), .b(gate209inter1), .O(G690));
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );

  xor2  gate715(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate716(.a(gate221inter0), .b(s_24), .O(gate221inter1));
  and2  gate717(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate718(.a(s_24), .O(gate221inter3));
  inv1  gate719(.a(s_25), .O(gate221inter4));
  nand2 gate720(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate721(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate722(.a(G622), .O(gate221inter7));
  inv1  gate723(.a(G684), .O(gate221inter8));
  nand2 gate724(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate725(.a(s_25), .b(gate221inter3), .O(gate221inter10));
  nor2  gate726(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate727(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate728(.a(gate221inter12), .b(gate221inter1), .O(G702));

  xor2  gate1009(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate1010(.a(gate222inter0), .b(s_66), .O(gate222inter1));
  and2  gate1011(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate1012(.a(s_66), .O(gate222inter3));
  inv1  gate1013(.a(s_67), .O(gate222inter4));
  nand2 gate1014(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate1015(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate1016(.a(G632), .O(gate222inter7));
  inv1  gate1017(.a(G684), .O(gate222inter8));
  nand2 gate1018(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate1019(.a(s_67), .b(gate222inter3), .O(gate222inter10));
  nor2  gate1020(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate1021(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate1022(.a(gate222inter12), .b(gate222inter1), .O(G703));
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate687(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate688(.a(gate226inter0), .b(s_20), .O(gate226inter1));
  and2  gate689(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate690(.a(s_20), .O(gate226inter3));
  inv1  gate691(.a(s_21), .O(gate226inter4));
  nand2 gate692(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate693(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate694(.a(G692), .O(gate226inter7));
  inv1  gate695(.a(G693), .O(gate226inter8));
  nand2 gate696(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate697(.a(s_21), .b(gate226inter3), .O(gate226inter10));
  nor2  gate698(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate699(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate700(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );

  xor2  gate1499(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate1500(.a(gate230inter0), .b(s_136), .O(gate230inter1));
  and2  gate1501(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate1502(.a(s_136), .O(gate230inter3));
  inv1  gate1503(.a(s_137), .O(gate230inter4));
  nand2 gate1504(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate1505(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate1506(.a(G700), .O(gate230inter7));
  inv1  gate1507(.a(G701), .O(gate230inter8));
  nand2 gate1508(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate1509(.a(s_137), .b(gate230inter3), .O(gate230inter10));
  nor2  gate1510(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate1511(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate1512(.a(gate230inter12), .b(gate230inter1), .O(G721));
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate1233(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate1234(.a(gate233inter0), .b(s_98), .O(gate233inter1));
  and2  gate1235(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate1236(.a(s_98), .O(gate233inter3));
  inv1  gate1237(.a(s_99), .O(gate233inter4));
  nand2 gate1238(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1239(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1240(.a(G242), .O(gate233inter7));
  inv1  gate1241(.a(G718), .O(gate233inter8));
  nand2 gate1242(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1243(.a(s_99), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1244(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1245(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1246(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );

  xor2  gate1247(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate1248(.a(gate238inter0), .b(s_100), .O(gate238inter1));
  and2  gate1249(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate1250(.a(s_100), .O(gate238inter3));
  inv1  gate1251(.a(s_101), .O(gate238inter4));
  nand2 gate1252(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate1253(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate1254(.a(G257), .O(gate238inter7));
  inv1  gate1255(.a(G709), .O(gate238inter8));
  nand2 gate1256(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate1257(.a(s_101), .b(gate238inter3), .O(gate238inter10));
  nor2  gate1258(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate1259(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate1260(.a(gate238inter12), .b(gate238inter1), .O(G745));

  xor2  gate1177(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate1178(.a(gate239inter0), .b(s_90), .O(gate239inter1));
  and2  gate1179(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate1180(.a(s_90), .O(gate239inter3));
  inv1  gate1181(.a(s_91), .O(gate239inter4));
  nand2 gate1182(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate1183(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate1184(.a(G260), .O(gate239inter7));
  inv1  gate1185(.a(G712), .O(gate239inter8));
  nand2 gate1186(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate1187(.a(s_91), .b(gate239inter3), .O(gate239inter10));
  nor2  gate1188(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate1189(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate1190(.a(gate239inter12), .b(gate239inter1), .O(G748));
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );

  xor2  gate1611(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate1612(.a(gate242inter0), .b(s_152), .O(gate242inter1));
  and2  gate1613(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate1614(.a(s_152), .O(gate242inter3));
  inv1  gate1615(.a(s_153), .O(gate242inter4));
  nand2 gate1616(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate1617(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate1618(.a(G718), .O(gate242inter7));
  inv1  gate1619(.a(G730), .O(gate242inter8));
  nand2 gate1620(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate1621(.a(s_153), .b(gate242inter3), .O(gate242inter10));
  nor2  gate1622(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate1623(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate1624(.a(gate242inter12), .b(gate242inter1), .O(G755));
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate673(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate674(.a(gate245inter0), .b(s_18), .O(gate245inter1));
  and2  gate675(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate676(.a(s_18), .O(gate245inter3));
  inv1  gate677(.a(s_19), .O(gate245inter4));
  nand2 gate678(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate679(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate680(.a(G248), .O(gate245inter7));
  inv1  gate681(.a(G736), .O(gate245inter8));
  nand2 gate682(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate683(.a(s_19), .b(gate245inter3), .O(gate245inter10));
  nor2  gate684(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate685(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate686(.a(gate245inter12), .b(gate245inter1), .O(G758));

  xor2  gate911(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate912(.a(gate246inter0), .b(s_52), .O(gate246inter1));
  and2  gate913(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate914(.a(s_52), .O(gate246inter3));
  inv1  gate915(.a(s_53), .O(gate246inter4));
  nand2 gate916(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate917(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate918(.a(G724), .O(gate246inter7));
  inv1  gate919(.a(G736), .O(gate246inter8));
  nand2 gate920(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate921(.a(s_53), .b(gate246inter3), .O(gate246inter10));
  nor2  gate922(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate923(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate924(.a(gate246inter12), .b(gate246inter1), .O(G759));
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate645(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate646(.a(gate250inter0), .b(s_14), .O(gate250inter1));
  and2  gate647(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate648(.a(s_14), .O(gate250inter3));
  inv1  gate649(.a(s_15), .O(gate250inter4));
  nand2 gate650(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate651(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate652(.a(G706), .O(gate250inter7));
  inv1  gate653(.a(G742), .O(gate250inter8));
  nand2 gate654(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate655(.a(s_15), .b(gate250inter3), .O(gate250inter10));
  nor2  gate656(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate657(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate658(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate1849(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate1850(.a(gate261inter0), .b(s_186), .O(gate261inter1));
  and2  gate1851(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate1852(.a(s_186), .O(gate261inter3));
  inv1  gate1853(.a(s_187), .O(gate261inter4));
  nand2 gate1854(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate1855(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate1856(.a(G762), .O(gate261inter7));
  inv1  gate1857(.a(G763), .O(gate261inter8));
  nand2 gate1858(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate1859(.a(s_187), .b(gate261inter3), .O(gate261inter10));
  nor2  gate1860(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate1861(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate1862(.a(gate261inter12), .b(gate261inter1), .O(G782));
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );

  xor2  gate1065(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate1066(.a(gate275inter0), .b(s_74), .O(gate275inter1));
  and2  gate1067(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate1068(.a(s_74), .O(gate275inter3));
  inv1  gate1069(.a(s_75), .O(gate275inter4));
  nand2 gate1070(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate1071(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate1072(.a(G645), .O(gate275inter7));
  inv1  gate1073(.a(G797), .O(gate275inter8));
  nand2 gate1074(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate1075(.a(s_75), .b(gate275inter3), .O(gate275inter10));
  nor2  gate1076(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate1077(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate1078(.a(gate275inter12), .b(gate275inter1), .O(G820));
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate659(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate660(.a(gate279inter0), .b(s_16), .O(gate279inter1));
  and2  gate661(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate662(.a(s_16), .O(gate279inter3));
  inv1  gate663(.a(s_17), .O(gate279inter4));
  nand2 gate664(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate665(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate666(.a(G651), .O(gate279inter7));
  inv1  gate667(.a(G803), .O(gate279inter8));
  nand2 gate668(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate669(.a(s_17), .b(gate279inter3), .O(gate279inter10));
  nor2  gate670(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate671(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate672(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate1373(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate1374(.a(gate283inter0), .b(s_118), .O(gate283inter1));
  and2  gate1375(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate1376(.a(s_118), .O(gate283inter3));
  inv1  gate1377(.a(s_119), .O(gate283inter4));
  nand2 gate1378(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate1379(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate1380(.a(G657), .O(gate283inter7));
  inv1  gate1381(.a(G809), .O(gate283inter8));
  nand2 gate1382(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate1383(.a(s_119), .b(gate283inter3), .O(gate283inter10));
  nor2  gate1384(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate1385(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate1386(.a(gate283inter12), .b(gate283inter1), .O(G828));

  xor2  gate1863(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate1864(.a(gate284inter0), .b(s_188), .O(gate284inter1));
  and2  gate1865(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate1866(.a(s_188), .O(gate284inter3));
  inv1  gate1867(.a(s_189), .O(gate284inter4));
  nand2 gate1868(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate1869(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate1870(.a(G785), .O(gate284inter7));
  inv1  gate1871(.a(G809), .O(gate284inter8));
  nand2 gate1872(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate1873(.a(s_189), .b(gate284inter3), .O(gate284inter10));
  nor2  gate1874(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate1875(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate1876(.a(gate284inter12), .b(gate284inter1), .O(G829));

  xor2  gate1933(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate1934(.a(gate285inter0), .b(s_198), .O(gate285inter1));
  and2  gate1935(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate1936(.a(s_198), .O(gate285inter3));
  inv1  gate1937(.a(s_199), .O(gate285inter4));
  nand2 gate1938(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate1939(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate1940(.a(G660), .O(gate285inter7));
  inv1  gate1941(.a(G812), .O(gate285inter8));
  nand2 gate1942(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate1943(.a(s_199), .b(gate285inter3), .O(gate285inter10));
  nor2  gate1944(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate1945(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate1946(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate1723(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate1724(.a(gate287inter0), .b(s_168), .O(gate287inter1));
  and2  gate1725(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate1726(.a(s_168), .O(gate287inter3));
  inv1  gate1727(.a(s_169), .O(gate287inter4));
  nand2 gate1728(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate1729(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate1730(.a(G663), .O(gate287inter7));
  inv1  gate1731(.a(G815), .O(gate287inter8));
  nand2 gate1732(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate1733(.a(s_169), .b(gate287inter3), .O(gate287inter10));
  nor2  gate1734(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate1735(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate1736(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate1653(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate1654(.a(gate289inter0), .b(s_158), .O(gate289inter1));
  and2  gate1655(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate1656(.a(s_158), .O(gate289inter3));
  inv1  gate1657(.a(s_159), .O(gate289inter4));
  nand2 gate1658(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate1659(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate1660(.a(G818), .O(gate289inter7));
  inv1  gate1661(.a(G819), .O(gate289inter8));
  nand2 gate1662(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate1663(.a(s_159), .b(gate289inter3), .O(gate289inter10));
  nor2  gate1664(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate1665(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate1666(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate1205(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate1206(.a(gate291inter0), .b(s_94), .O(gate291inter1));
  and2  gate1207(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate1208(.a(s_94), .O(gate291inter3));
  inv1  gate1209(.a(s_95), .O(gate291inter4));
  nand2 gate1210(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate1211(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate1212(.a(G822), .O(gate291inter7));
  inv1  gate1213(.a(G823), .O(gate291inter8));
  nand2 gate1214(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate1215(.a(s_95), .b(gate291inter3), .O(gate291inter10));
  nor2  gate1216(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate1217(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate1218(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate1457(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate1458(.a(gate293inter0), .b(s_130), .O(gate293inter1));
  and2  gate1459(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate1460(.a(s_130), .O(gate293inter3));
  inv1  gate1461(.a(s_131), .O(gate293inter4));
  nand2 gate1462(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate1463(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate1464(.a(G828), .O(gate293inter7));
  inv1  gate1465(.a(G829), .O(gate293inter8));
  nand2 gate1466(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate1467(.a(s_131), .b(gate293inter3), .O(gate293inter10));
  nor2  gate1468(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate1469(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate1470(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate1359(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate1360(.a(gate388inter0), .b(s_116), .O(gate388inter1));
  and2  gate1361(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate1362(.a(s_116), .O(gate388inter3));
  inv1  gate1363(.a(s_117), .O(gate388inter4));
  nand2 gate1364(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate1365(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate1366(.a(G2), .O(gate388inter7));
  inv1  gate1367(.a(G1039), .O(gate388inter8));
  nand2 gate1368(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate1369(.a(s_117), .b(gate388inter3), .O(gate388inter10));
  nor2  gate1370(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate1371(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate1372(.a(gate388inter12), .b(gate388inter1), .O(G1135));
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate1793(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate1794(.a(gate390inter0), .b(s_178), .O(gate390inter1));
  and2  gate1795(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate1796(.a(s_178), .O(gate390inter3));
  inv1  gate1797(.a(s_179), .O(gate390inter4));
  nand2 gate1798(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate1799(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate1800(.a(G4), .O(gate390inter7));
  inv1  gate1801(.a(G1045), .O(gate390inter8));
  nand2 gate1802(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate1803(.a(s_179), .b(gate390inter3), .O(gate390inter10));
  nor2  gate1804(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate1805(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate1806(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate2003(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate2004(.a(gate395inter0), .b(s_208), .O(gate395inter1));
  and2  gate2005(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate2006(.a(s_208), .O(gate395inter3));
  inv1  gate2007(.a(s_209), .O(gate395inter4));
  nand2 gate2008(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate2009(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate2010(.a(G9), .O(gate395inter7));
  inv1  gate2011(.a(G1060), .O(gate395inter8));
  nand2 gate2012(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate2013(.a(s_209), .b(gate395inter3), .O(gate395inter10));
  nor2  gate2014(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate2015(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate2016(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate1779(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate1780(.a(gate398inter0), .b(s_176), .O(gate398inter1));
  and2  gate1781(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate1782(.a(s_176), .O(gate398inter3));
  inv1  gate1783(.a(s_177), .O(gate398inter4));
  nand2 gate1784(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate1785(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate1786(.a(G12), .O(gate398inter7));
  inv1  gate1787(.a(G1069), .O(gate398inter8));
  nand2 gate1788(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate1789(.a(s_177), .b(gate398inter3), .O(gate398inter10));
  nor2  gate1790(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate1791(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate1792(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate547(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate548(.a(gate403inter0), .b(s_0), .O(gate403inter1));
  and2  gate549(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate550(.a(s_0), .O(gate403inter3));
  inv1  gate551(.a(s_1), .O(gate403inter4));
  nand2 gate552(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate553(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate554(.a(G17), .O(gate403inter7));
  inv1  gate555(.a(G1084), .O(gate403inter8));
  nand2 gate556(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate557(.a(s_1), .b(gate403inter3), .O(gate403inter10));
  nor2  gate558(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate559(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate560(.a(gate403inter12), .b(gate403inter1), .O(G1180));

  xor2  gate631(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate632(.a(gate404inter0), .b(s_12), .O(gate404inter1));
  and2  gate633(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate634(.a(s_12), .O(gate404inter3));
  inv1  gate635(.a(s_13), .O(gate404inter4));
  nand2 gate636(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate637(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate638(.a(G18), .O(gate404inter7));
  inv1  gate639(.a(G1087), .O(gate404inter8));
  nand2 gate640(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate641(.a(s_13), .b(gate404inter3), .O(gate404inter10));
  nor2  gate642(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate643(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate644(.a(gate404inter12), .b(gate404inter1), .O(G1183));

  xor2  gate1107(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate1108(.a(gate405inter0), .b(s_80), .O(gate405inter1));
  and2  gate1109(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate1110(.a(s_80), .O(gate405inter3));
  inv1  gate1111(.a(s_81), .O(gate405inter4));
  nand2 gate1112(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate1113(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate1114(.a(G19), .O(gate405inter7));
  inv1  gate1115(.a(G1090), .O(gate405inter8));
  nand2 gate1116(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate1117(.a(s_81), .b(gate405inter3), .O(gate405inter10));
  nor2  gate1118(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate1119(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate1120(.a(gate405inter12), .b(gate405inter1), .O(G1186));

  xor2  gate1695(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate1696(.a(gate406inter0), .b(s_164), .O(gate406inter1));
  and2  gate1697(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate1698(.a(s_164), .O(gate406inter3));
  inv1  gate1699(.a(s_165), .O(gate406inter4));
  nand2 gate1700(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate1701(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate1702(.a(G20), .O(gate406inter7));
  inv1  gate1703(.a(G1093), .O(gate406inter8));
  nand2 gate1704(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate1705(.a(s_165), .b(gate406inter3), .O(gate406inter10));
  nor2  gate1706(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate1707(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate1708(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate1303(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate1304(.a(gate410inter0), .b(s_108), .O(gate410inter1));
  and2  gate1305(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate1306(.a(s_108), .O(gate410inter3));
  inv1  gate1307(.a(s_109), .O(gate410inter4));
  nand2 gate1308(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate1309(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate1310(.a(G24), .O(gate410inter7));
  inv1  gate1311(.a(G1105), .O(gate410inter8));
  nand2 gate1312(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate1313(.a(s_109), .b(gate410inter3), .O(gate410inter10));
  nor2  gate1314(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate1315(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate1316(.a(gate410inter12), .b(gate410inter1), .O(G1201));

  xor2  gate1905(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate1906(.a(gate411inter0), .b(s_194), .O(gate411inter1));
  and2  gate1907(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate1908(.a(s_194), .O(gate411inter3));
  inv1  gate1909(.a(s_195), .O(gate411inter4));
  nand2 gate1910(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate1911(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate1912(.a(G25), .O(gate411inter7));
  inv1  gate1913(.a(G1108), .O(gate411inter8));
  nand2 gate1914(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate1915(.a(s_195), .b(gate411inter3), .O(gate411inter10));
  nor2  gate1916(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate1917(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate1918(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );

  xor2  gate603(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate604(.a(gate414inter0), .b(s_8), .O(gate414inter1));
  and2  gate605(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate606(.a(s_8), .O(gate414inter3));
  inv1  gate607(.a(s_9), .O(gate414inter4));
  nand2 gate608(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate609(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate610(.a(G28), .O(gate414inter7));
  inv1  gate611(.a(G1117), .O(gate414inter8));
  nand2 gate612(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate613(.a(s_9), .b(gate414inter3), .O(gate414inter10));
  nor2  gate614(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate615(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate616(.a(gate414inter12), .b(gate414inter1), .O(G1213));
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate869(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate870(.a(gate417inter0), .b(s_46), .O(gate417inter1));
  and2  gate871(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate872(.a(s_46), .O(gate417inter3));
  inv1  gate873(.a(s_47), .O(gate417inter4));
  nand2 gate874(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate875(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate876(.a(G31), .O(gate417inter7));
  inv1  gate877(.a(G1126), .O(gate417inter8));
  nand2 gate878(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate879(.a(s_47), .b(gate417inter3), .O(gate417inter10));
  nor2  gate880(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate881(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate882(.a(gate417inter12), .b(gate417inter1), .O(G1222));

  xor2  gate813(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate814(.a(gate418inter0), .b(s_38), .O(gate418inter1));
  and2  gate815(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate816(.a(s_38), .O(gate418inter3));
  inv1  gate817(.a(s_39), .O(gate418inter4));
  nand2 gate818(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate819(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate820(.a(G32), .O(gate418inter7));
  inv1  gate821(.a(G1129), .O(gate418inter8));
  nand2 gate822(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate823(.a(s_39), .b(gate418inter3), .O(gate418inter10));
  nor2  gate824(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate825(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate826(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate995(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate996(.a(gate421inter0), .b(s_64), .O(gate421inter1));
  and2  gate997(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate998(.a(s_64), .O(gate421inter3));
  inv1  gate999(.a(s_65), .O(gate421inter4));
  nand2 gate1000(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate1001(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate1002(.a(G2), .O(gate421inter7));
  inv1  gate1003(.a(G1135), .O(gate421inter8));
  nand2 gate1004(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate1005(.a(s_65), .b(gate421inter3), .O(gate421inter10));
  nor2  gate1006(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate1007(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate1008(.a(gate421inter12), .b(gate421inter1), .O(G1230));

  xor2  gate827(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate828(.a(gate422inter0), .b(s_40), .O(gate422inter1));
  and2  gate829(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate830(.a(s_40), .O(gate422inter3));
  inv1  gate831(.a(s_41), .O(gate422inter4));
  nand2 gate832(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate833(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate834(.a(G1039), .O(gate422inter7));
  inv1  gate835(.a(G1135), .O(gate422inter8));
  nand2 gate836(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate837(.a(s_41), .b(gate422inter3), .O(gate422inter10));
  nor2  gate838(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate839(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate840(.a(gate422inter12), .b(gate422inter1), .O(G1231));

  xor2  gate1471(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate1472(.a(gate423inter0), .b(s_132), .O(gate423inter1));
  and2  gate1473(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate1474(.a(s_132), .O(gate423inter3));
  inv1  gate1475(.a(s_133), .O(gate423inter4));
  nand2 gate1476(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate1477(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate1478(.a(G3), .O(gate423inter7));
  inv1  gate1479(.a(G1138), .O(gate423inter8));
  nand2 gate1480(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate1481(.a(s_133), .b(gate423inter3), .O(gate423inter10));
  nor2  gate1482(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate1483(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate1484(.a(gate423inter12), .b(gate423inter1), .O(G1232));
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );

  xor2  gate1709(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate1710(.a(gate427inter0), .b(s_166), .O(gate427inter1));
  and2  gate1711(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate1712(.a(s_166), .O(gate427inter3));
  inv1  gate1713(.a(s_167), .O(gate427inter4));
  nand2 gate1714(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate1715(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate1716(.a(G5), .O(gate427inter7));
  inv1  gate1717(.a(G1144), .O(gate427inter8));
  nand2 gate1718(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate1719(.a(s_167), .b(gate427inter3), .O(gate427inter10));
  nor2  gate1720(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate1721(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate1722(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate981(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate982(.a(gate430inter0), .b(s_62), .O(gate430inter1));
  and2  gate983(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate984(.a(s_62), .O(gate430inter3));
  inv1  gate985(.a(s_63), .O(gate430inter4));
  nand2 gate986(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate987(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate988(.a(G1051), .O(gate430inter7));
  inv1  gate989(.a(G1147), .O(gate430inter8));
  nand2 gate990(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate991(.a(s_63), .b(gate430inter3), .O(gate430inter10));
  nor2  gate992(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate993(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate994(.a(gate430inter12), .b(gate430inter1), .O(G1239));

  xor2  gate967(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate968(.a(gate431inter0), .b(s_60), .O(gate431inter1));
  and2  gate969(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate970(.a(s_60), .O(gate431inter3));
  inv1  gate971(.a(s_61), .O(gate431inter4));
  nand2 gate972(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate973(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate974(.a(G7), .O(gate431inter7));
  inv1  gate975(.a(G1150), .O(gate431inter8));
  nand2 gate976(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate977(.a(s_61), .b(gate431inter3), .O(gate431inter10));
  nor2  gate978(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate979(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate980(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate1121(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate1122(.a(gate444inter0), .b(s_82), .O(gate444inter1));
  and2  gate1123(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate1124(.a(s_82), .O(gate444inter3));
  inv1  gate1125(.a(s_83), .O(gate444inter4));
  nand2 gate1126(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate1127(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate1128(.a(G1072), .O(gate444inter7));
  inv1  gate1129(.a(G1168), .O(gate444inter8));
  nand2 gate1130(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate1131(.a(s_83), .b(gate444inter3), .O(gate444inter10));
  nor2  gate1132(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate1133(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate1134(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );

  xor2  gate841(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate842(.a(gate450inter0), .b(s_42), .O(gate450inter1));
  and2  gate843(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate844(.a(s_42), .O(gate450inter3));
  inv1  gate845(.a(s_43), .O(gate450inter4));
  nand2 gate846(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate847(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate848(.a(G1081), .O(gate450inter7));
  inv1  gate849(.a(G1177), .O(gate450inter8));
  nand2 gate850(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate851(.a(s_43), .b(gate450inter3), .O(gate450inter10));
  nor2  gate852(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate853(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate854(.a(gate450inter12), .b(gate450inter1), .O(G1259));
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );

  xor2  gate1989(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate1990(.a(gate454inter0), .b(s_206), .O(gate454inter1));
  and2  gate1991(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate1992(.a(s_206), .O(gate454inter3));
  inv1  gate1993(.a(s_207), .O(gate454inter4));
  nand2 gate1994(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate1995(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate1996(.a(G1087), .O(gate454inter7));
  inv1  gate1997(.a(G1183), .O(gate454inter8));
  nand2 gate1998(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate1999(.a(s_207), .b(gate454inter3), .O(gate454inter10));
  nor2  gate2000(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate2001(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate2002(.a(gate454inter12), .b(gate454inter1), .O(G1263));
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate701(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate702(.a(gate463inter0), .b(s_22), .O(gate463inter1));
  and2  gate703(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate704(.a(s_22), .O(gate463inter3));
  inv1  gate705(.a(s_23), .O(gate463inter4));
  nand2 gate706(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate707(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate708(.a(G23), .O(gate463inter7));
  inv1  gate709(.a(G1198), .O(gate463inter8));
  nand2 gate710(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate711(.a(s_23), .b(gate463inter3), .O(gate463inter10));
  nor2  gate712(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate713(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate714(.a(gate463inter12), .b(gate463inter1), .O(G1272));

  xor2  gate729(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate730(.a(gate464inter0), .b(s_26), .O(gate464inter1));
  and2  gate731(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate732(.a(s_26), .O(gate464inter3));
  inv1  gate733(.a(s_27), .O(gate464inter4));
  nand2 gate734(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate735(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate736(.a(G1102), .O(gate464inter7));
  inv1  gate737(.a(G1198), .O(gate464inter8));
  nand2 gate738(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate739(.a(s_27), .b(gate464inter3), .O(gate464inter10));
  nor2  gate740(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate741(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate742(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate1331(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate1332(.a(gate471inter0), .b(s_112), .O(gate471inter1));
  and2  gate1333(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate1334(.a(s_112), .O(gate471inter3));
  inv1  gate1335(.a(s_113), .O(gate471inter4));
  nand2 gate1336(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate1337(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate1338(.a(G27), .O(gate471inter7));
  inv1  gate1339(.a(G1210), .O(gate471inter8));
  nand2 gate1340(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate1341(.a(s_113), .b(gate471inter3), .O(gate471inter10));
  nor2  gate1342(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate1343(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate1344(.a(gate471inter12), .b(gate471inter1), .O(G1280));

  xor2  gate1681(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate1682(.a(gate472inter0), .b(s_162), .O(gate472inter1));
  and2  gate1683(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate1684(.a(s_162), .O(gate472inter3));
  inv1  gate1685(.a(s_163), .O(gate472inter4));
  nand2 gate1686(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate1687(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate1688(.a(G1114), .O(gate472inter7));
  inv1  gate1689(.a(G1210), .O(gate472inter8));
  nand2 gate1690(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate1691(.a(s_163), .b(gate472inter3), .O(gate472inter10));
  nor2  gate1692(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate1693(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate1694(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate1079(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate1080(.a(gate474inter0), .b(s_76), .O(gate474inter1));
  and2  gate1081(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate1082(.a(s_76), .O(gate474inter3));
  inv1  gate1083(.a(s_77), .O(gate474inter4));
  nand2 gate1084(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate1085(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate1086(.a(G1117), .O(gate474inter7));
  inv1  gate1087(.a(G1213), .O(gate474inter8));
  nand2 gate1088(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate1089(.a(s_77), .b(gate474inter3), .O(gate474inter10));
  nor2  gate1090(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate1091(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate1092(.a(gate474inter12), .b(gate474inter1), .O(G1283));

  xor2  gate1135(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate1136(.a(gate475inter0), .b(s_84), .O(gate475inter1));
  and2  gate1137(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate1138(.a(s_84), .O(gate475inter3));
  inv1  gate1139(.a(s_85), .O(gate475inter4));
  nand2 gate1140(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate1141(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate1142(.a(G29), .O(gate475inter7));
  inv1  gate1143(.a(G1216), .O(gate475inter8));
  nand2 gate1144(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate1145(.a(s_85), .b(gate475inter3), .O(gate475inter10));
  nor2  gate1146(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate1147(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate1148(.a(gate475inter12), .b(gate475inter1), .O(G1284));
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );

  xor2  gate1443(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate1444(.a(gate479inter0), .b(s_128), .O(gate479inter1));
  and2  gate1445(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate1446(.a(s_128), .O(gate479inter3));
  inv1  gate1447(.a(s_129), .O(gate479inter4));
  nand2 gate1448(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate1449(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate1450(.a(G31), .O(gate479inter7));
  inv1  gate1451(.a(G1222), .O(gate479inter8));
  nand2 gate1452(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate1453(.a(s_129), .b(gate479inter3), .O(gate479inter10));
  nor2  gate1454(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate1455(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate1456(.a(gate479inter12), .b(gate479inter1), .O(G1288));

  xor2  gate1149(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate1150(.a(gate480inter0), .b(s_86), .O(gate480inter1));
  and2  gate1151(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate1152(.a(s_86), .O(gate480inter3));
  inv1  gate1153(.a(s_87), .O(gate480inter4));
  nand2 gate1154(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate1155(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate1156(.a(G1126), .O(gate480inter7));
  inv1  gate1157(.a(G1222), .O(gate480inter8));
  nand2 gate1158(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate1159(.a(s_87), .b(gate480inter3), .O(gate480inter10));
  nor2  gate1160(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate1161(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate1162(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate1345(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate1346(.a(gate482inter0), .b(s_114), .O(gate482inter1));
  and2  gate1347(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate1348(.a(s_114), .O(gate482inter3));
  inv1  gate1349(.a(s_115), .O(gate482inter4));
  nand2 gate1350(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate1351(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate1352(.a(G1129), .O(gate482inter7));
  inv1  gate1353(.a(G1225), .O(gate482inter8));
  nand2 gate1354(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate1355(.a(s_115), .b(gate482inter3), .O(gate482inter10));
  nor2  gate1356(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate1357(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate1358(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate1051(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate1052(.a(gate485inter0), .b(s_72), .O(gate485inter1));
  and2  gate1053(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate1054(.a(s_72), .O(gate485inter3));
  inv1  gate1055(.a(s_73), .O(gate485inter4));
  nand2 gate1056(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate1057(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate1058(.a(G1232), .O(gate485inter7));
  inv1  gate1059(.a(G1233), .O(gate485inter8));
  nand2 gate1060(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate1061(.a(s_73), .b(gate485inter3), .O(gate485inter10));
  nor2  gate1062(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate1063(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate1064(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );

  xor2  gate1583(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate1584(.a(gate498inter0), .b(s_148), .O(gate498inter1));
  and2  gate1585(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate1586(.a(s_148), .O(gate498inter3));
  inv1  gate1587(.a(s_149), .O(gate498inter4));
  nand2 gate1588(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate1589(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate1590(.a(G1258), .O(gate498inter7));
  inv1  gate1591(.a(G1259), .O(gate498inter8));
  nand2 gate1592(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate1593(.a(s_149), .b(gate498inter3), .O(gate498inter10));
  nor2  gate1594(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate1595(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate1596(.a(gate498inter12), .b(gate498inter1), .O(G1307));

  xor2  gate1667(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate1668(.a(gate499inter0), .b(s_160), .O(gate499inter1));
  and2  gate1669(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate1670(.a(s_160), .O(gate499inter3));
  inv1  gate1671(.a(s_161), .O(gate499inter4));
  nand2 gate1672(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate1673(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate1674(.a(G1260), .O(gate499inter7));
  inv1  gate1675(.a(G1261), .O(gate499inter8));
  nand2 gate1676(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate1677(.a(s_161), .b(gate499inter3), .O(gate499inter10));
  nor2  gate1678(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate1679(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate1680(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate939(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate940(.a(gate501inter0), .b(s_56), .O(gate501inter1));
  and2  gate941(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate942(.a(s_56), .O(gate501inter3));
  inv1  gate943(.a(s_57), .O(gate501inter4));
  nand2 gate944(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate945(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate946(.a(G1264), .O(gate501inter7));
  inv1  gate947(.a(G1265), .O(gate501inter8));
  nand2 gate948(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate949(.a(s_57), .b(gate501inter3), .O(gate501inter10));
  nor2  gate950(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate951(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate952(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );

  xor2  gate1163(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate1164(.a(gate505inter0), .b(s_88), .O(gate505inter1));
  and2  gate1165(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate1166(.a(s_88), .O(gate505inter3));
  inv1  gate1167(.a(s_89), .O(gate505inter4));
  nand2 gate1168(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate1169(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate1170(.a(G1272), .O(gate505inter7));
  inv1  gate1171(.a(G1273), .O(gate505inter8));
  nand2 gate1172(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate1173(.a(s_89), .b(gate505inter3), .O(gate505inter10));
  nor2  gate1174(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate1175(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate1176(.a(gate505inter12), .b(gate505inter1), .O(G1314));
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate771(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate772(.a(gate509inter0), .b(s_32), .O(gate509inter1));
  and2  gate773(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate774(.a(s_32), .O(gate509inter3));
  inv1  gate775(.a(s_33), .O(gate509inter4));
  nand2 gate776(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate777(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate778(.a(G1280), .O(gate509inter7));
  inv1  gate779(.a(G1281), .O(gate509inter8));
  nand2 gate780(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate781(.a(s_33), .b(gate509inter3), .O(gate509inter10));
  nor2  gate782(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate783(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate784(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule