module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate981(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate982(.a(gate17inter0), .b(s_62), .O(gate17inter1));
  and2  gate983(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate984(.a(s_62), .O(gate17inter3));
  inv1  gate985(.a(s_63), .O(gate17inter4));
  nand2 gate986(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate987(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate988(.a(G17), .O(gate17inter7));
  inv1  gate989(.a(G18), .O(gate17inter8));
  nand2 gate990(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate991(.a(s_63), .b(gate17inter3), .O(gate17inter10));
  nor2  gate992(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate993(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate994(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate617(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate618(.a(gate24inter0), .b(s_10), .O(gate24inter1));
  and2  gate619(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate620(.a(s_10), .O(gate24inter3));
  inv1  gate621(.a(s_11), .O(gate24inter4));
  nand2 gate622(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate623(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate624(.a(G31), .O(gate24inter7));
  inv1  gate625(.a(G32), .O(gate24inter8));
  nand2 gate626(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate627(.a(s_11), .b(gate24inter3), .O(gate24inter10));
  nor2  gate628(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate629(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate630(.a(gate24inter12), .b(gate24inter1), .O(G311));

  xor2  gate1149(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate1150(.a(gate25inter0), .b(s_86), .O(gate25inter1));
  and2  gate1151(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate1152(.a(s_86), .O(gate25inter3));
  inv1  gate1153(.a(s_87), .O(gate25inter4));
  nand2 gate1154(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate1155(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate1156(.a(G1), .O(gate25inter7));
  inv1  gate1157(.a(G5), .O(gate25inter8));
  nand2 gate1158(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate1159(.a(s_87), .b(gate25inter3), .O(gate25inter10));
  nor2  gate1160(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate1161(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate1162(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate1023(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate1024(.a(gate37inter0), .b(s_68), .O(gate37inter1));
  and2  gate1025(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate1026(.a(s_68), .O(gate37inter3));
  inv1  gate1027(.a(s_69), .O(gate37inter4));
  nand2 gate1028(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate1029(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate1030(.a(G19), .O(gate37inter7));
  inv1  gate1031(.a(G23), .O(gate37inter8));
  nand2 gate1032(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate1033(.a(s_69), .b(gate37inter3), .O(gate37inter10));
  nor2  gate1034(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate1035(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate1036(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate953(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate954(.a(gate41inter0), .b(s_58), .O(gate41inter1));
  and2  gate955(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate956(.a(s_58), .O(gate41inter3));
  inv1  gate957(.a(s_59), .O(gate41inter4));
  nand2 gate958(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate959(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate960(.a(G1), .O(gate41inter7));
  inv1  gate961(.a(G266), .O(gate41inter8));
  nand2 gate962(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate963(.a(s_59), .b(gate41inter3), .O(gate41inter10));
  nor2  gate964(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate965(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate966(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate659(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate660(.a(gate62inter0), .b(s_16), .O(gate62inter1));
  and2  gate661(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate662(.a(s_16), .O(gate62inter3));
  inv1  gate663(.a(s_17), .O(gate62inter4));
  nand2 gate664(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate665(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate666(.a(G22), .O(gate62inter7));
  inv1  gate667(.a(G296), .O(gate62inter8));
  nand2 gate668(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate669(.a(s_17), .b(gate62inter3), .O(gate62inter10));
  nor2  gate670(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate671(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate672(.a(gate62inter12), .b(gate62inter1), .O(G383));

  xor2  gate883(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate884(.a(gate63inter0), .b(s_48), .O(gate63inter1));
  and2  gate885(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate886(.a(s_48), .O(gate63inter3));
  inv1  gate887(.a(s_49), .O(gate63inter4));
  nand2 gate888(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate889(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate890(.a(G23), .O(gate63inter7));
  inv1  gate891(.a(G299), .O(gate63inter8));
  nand2 gate892(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate893(.a(s_49), .b(gate63inter3), .O(gate63inter10));
  nor2  gate894(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate895(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate896(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate687(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate688(.a(gate69inter0), .b(s_20), .O(gate69inter1));
  and2  gate689(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate690(.a(s_20), .O(gate69inter3));
  inv1  gate691(.a(s_21), .O(gate69inter4));
  nand2 gate692(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate693(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate694(.a(G29), .O(gate69inter7));
  inv1  gate695(.a(G308), .O(gate69inter8));
  nand2 gate696(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate697(.a(s_21), .b(gate69inter3), .O(gate69inter10));
  nor2  gate698(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate699(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate700(.a(gate69inter12), .b(gate69inter1), .O(G390));

  xor2  gate1079(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate1080(.a(gate70inter0), .b(s_76), .O(gate70inter1));
  and2  gate1081(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate1082(.a(s_76), .O(gate70inter3));
  inv1  gate1083(.a(s_77), .O(gate70inter4));
  nand2 gate1084(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate1085(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate1086(.a(G30), .O(gate70inter7));
  inv1  gate1087(.a(G308), .O(gate70inter8));
  nand2 gate1088(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate1089(.a(s_77), .b(gate70inter3), .O(gate70inter10));
  nor2  gate1090(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate1091(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate1092(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );

  xor2  gate1107(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate1108(.a(gate72inter0), .b(s_80), .O(gate72inter1));
  and2  gate1109(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate1110(.a(s_80), .O(gate72inter3));
  inv1  gate1111(.a(s_81), .O(gate72inter4));
  nand2 gate1112(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate1113(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate1114(.a(G32), .O(gate72inter7));
  inv1  gate1115(.a(G311), .O(gate72inter8));
  nand2 gate1116(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate1117(.a(s_81), .b(gate72inter3), .O(gate72inter10));
  nor2  gate1118(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate1119(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate1120(.a(gate72inter12), .b(gate72inter1), .O(G393));
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );

  xor2  gate1331(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate1332(.a(gate76inter0), .b(s_112), .O(gate76inter1));
  and2  gate1333(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate1334(.a(s_112), .O(gate76inter3));
  inv1  gate1335(.a(s_113), .O(gate76inter4));
  nand2 gate1336(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate1337(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate1338(.a(G13), .O(gate76inter7));
  inv1  gate1339(.a(G317), .O(gate76inter8));
  nand2 gate1340(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate1341(.a(s_113), .b(gate76inter3), .O(gate76inter10));
  nor2  gate1342(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate1343(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate1344(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate1065(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate1066(.a(gate81inter0), .b(s_74), .O(gate81inter1));
  and2  gate1067(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate1068(.a(s_74), .O(gate81inter3));
  inv1  gate1069(.a(s_75), .O(gate81inter4));
  nand2 gate1070(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate1071(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate1072(.a(G3), .O(gate81inter7));
  inv1  gate1073(.a(G326), .O(gate81inter8));
  nand2 gate1074(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate1075(.a(s_75), .b(gate81inter3), .O(gate81inter10));
  nor2  gate1076(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate1077(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate1078(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );

  xor2  gate925(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate926(.a(gate83inter0), .b(s_54), .O(gate83inter1));
  and2  gate927(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate928(.a(s_54), .O(gate83inter3));
  inv1  gate929(.a(s_55), .O(gate83inter4));
  nand2 gate930(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate931(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate932(.a(G11), .O(gate83inter7));
  inv1  gate933(.a(G329), .O(gate83inter8));
  nand2 gate934(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate935(.a(s_55), .b(gate83inter3), .O(gate83inter10));
  nor2  gate936(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate937(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate938(.a(gate83inter12), .b(gate83inter1), .O(G404));

  xor2  gate855(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate856(.a(gate84inter0), .b(s_44), .O(gate84inter1));
  and2  gate857(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate858(.a(s_44), .O(gate84inter3));
  inv1  gate859(.a(s_45), .O(gate84inter4));
  nand2 gate860(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate861(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate862(.a(G15), .O(gate84inter7));
  inv1  gate863(.a(G329), .O(gate84inter8));
  nand2 gate864(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate865(.a(s_45), .b(gate84inter3), .O(gate84inter10));
  nor2  gate866(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate867(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate868(.a(gate84inter12), .b(gate84inter1), .O(G405));
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate603(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate604(.a(gate86inter0), .b(s_8), .O(gate86inter1));
  and2  gate605(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate606(.a(s_8), .O(gate86inter3));
  inv1  gate607(.a(s_9), .O(gate86inter4));
  nand2 gate608(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate609(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate610(.a(G8), .O(gate86inter7));
  inv1  gate611(.a(G332), .O(gate86inter8));
  nand2 gate612(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate613(.a(s_9), .b(gate86inter3), .O(gate86inter10));
  nor2  gate614(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate615(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate616(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate785(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate786(.a(gate98inter0), .b(s_34), .O(gate98inter1));
  and2  gate787(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate788(.a(s_34), .O(gate98inter3));
  inv1  gate789(.a(s_35), .O(gate98inter4));
  nand2 gate790(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate791(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate792(.a(G23), .O(gate98inter7));
  inv1  gate793(.a(G350), .O(gate98inter8));
  nand2 gate794(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate795(.a(s_35), .b(gate98inter3), .O(gate98inter10));
  nor2  gate796(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate797(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate798(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );

  xor2  gate589(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate590(.a(gate101inter0), .b(s_6), .O(gate101inter1));
  and2  gate591(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate592(.a(s_6), .O(gate101inter3));
  inv1  gate593(.a(s_7), .O(gate101inter4));
  nand2 gate594(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate595(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate596(.a(G20), .O(gate101inter7));
  inv1  gate597(.a(G356), .O(gate101inter8));
  nand2 gate598(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate599(.a(s_7), .b(gate101inter3), .O(gate101inter10));
  nor2  gate600(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate601(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate602(.a(gate101inter12), .b(gate101inter1), .O(G422));
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate1177(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate1178(.a(gate108inter0), .b(s_90), .O(gate108inter1));
  and2  gate1179(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate1180(.a(s_90), .O(gate108inter3));
  inv1  gate1181(.a(s_91), .O(gate108inter4));
  nand2 gate1182(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate1183(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate1184(.a(G368), .O(gate108inter7));
  inv1  gate1185(.a(G369), .O(gate108inter8));
  nand2 gate1186(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate1187(.a(s_91), .b(gate108inter3), .O(gate108inter10));
  nor2  gate1188(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate1189(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate1190(.a(gate108inter12), .b(gate108inter1), .O(G435));
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate1359(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate1360(.a(gate110inter0), .b(s_116), .O(gate110inter1));
  and2  gate1361(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate1362(.a(s_116), .O(gate110inter3));
  inv1  gate1363(.a(s_117), .O(gate110inter4));
  nand2 gate1364(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1365(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1366(.a(G372), .O(gate110inter7));
  inv1  gate1367(.a(G373), .O(gate110inter8));
  nand2 gate1368(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1369(.a(s_117), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1370(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1371(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1372(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate1205(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate1206(.a(gate116inter0), .b(s_94), .O(gate116inter1));
  and2  gate1207(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate1208(.a(s_94), .O(gate116inter3));
  inv1  gate1209(.a(s_95), .O(gate116inter4));
  nand2 gate1210(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate1211(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate1212(.a(G384), .O(gate116inter7));
  inv1  gate1213(.a(G385), .O(gate116inter8));
  nand2 gate1214(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate1215(.a(s_95), .b(gate116inter3), .O(gate116inter10));
  nor2  gate1216(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate1217(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate1218(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate1051(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate1052(.a(gate123inter0), .b(s_72), .O(gate123inter1));
  and2  gate1053(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate1054(.a(s_72), .O(gate123inter3));
  inv1  gate1055(.a(s_73), .O(gate123inter4));
  nand2 gate1056(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate1057(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate1058(.a(G398), .O(gate123inter7));
  inv1  gate1059(.a(G399), .O(gate123inter8));
  nand2 gate1060(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate1061(.a(s_73), .b(gate123inter3), .O(gate123inter10));
  nor2  gate1062(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate1063(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate1064(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate673(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate674(.a(gate125inter0), .b(s_18), .O(gate125inter1));
  and2  gate675(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate676(.a(s_18), .O(gate125inter3));
  inv1  gate677(.a(s_19), .O(gate125inter4));
  nand2 gate678(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate679(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate680(.a(G402), .O(gate125inter7));
  inv1  gate681(.a(G403), .O(gate125inter8));
  nand2 gate682(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate683(.a(s_19), .b(gate125inter3), .O(gate125inter10));
  nor2  gate684(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate685(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate686(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate715(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate716(.a(gate144inter0), .b(s_24), .O(gate144inter1));
  and2  gate717(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate718(.a(s_24), .O(gate144inter3));
  inv1  gate719(.a(s_25), .O(gate144inter4));
  nand2 gate720(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate721(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate722(.a(G468), .O(gate144inter7));
  inv1  gate723(.a(G471), .O(gate144inter8));
  nand2 gate724(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate725(.a(s_25), .b(gate144inter3), .O(gate144inter10));
  nor2  gate726(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate727(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate728(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate1037(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate1038(.a(gate147inter0), .b(s_70), .O(gate147inter1));
  and2  gate1039(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate1040(.a(s_70), .O(gate147inter3));
  inv1  gate1041(.a(s_71), .O(gate147inter4));
  nand2 gate1042(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate1043(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate1044(.a(G486), .O(gate147inter7));
  inv1  gate1045(.a(G489), .O(gate147inter8));
  nand2 gate1046(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate1047(.a(s_71), .b(gate147inter3), .O(gate147inter10));
  nor2  gate1048(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate1049(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate1050(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate771(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate772(.a(gate159inter0), .b(s_32), .O(gate159inter1));
  and2  gate773(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate774(.a(s_32), .O(gate159inter3));
  inv1  gate775(.a(s_33), .O(gate159inter4));
  nand2 gate776(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate777(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate778(.a(G444), .O(gate159inter7));
  inv1  gate779(.a(G531), .O(gate159inter8));
  nand2 gate780(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate781(.a(s_33), .b(gate159inter3), .O(gate159inter10));
  nor2  gate782(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate783(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate784(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate967(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate968(.a(gate161inter0), .b(s_60), .O(gate161inter1));
  and2  gate969(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate970(.a(s_60), .O(gate161inter3));
  inv1  gate971(.a(s_61), .O(gate161inter4));
  nand2 gate972(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate973(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate974(.a(G450), .O(gate161inter7));
  inv1  gate975(.a(G534), .O(gate161inter8));
  nand2 gate976(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate977(.a(s_61), .b(gate161inter3), .O(gate161inter10));
  nor2  gate978(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate979(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate980(.a(gate161inter12), .b(gate161inter1), .O(G578));

  xor2  gate1121(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate1122(.a(gate162inter0), .b(s_82), .O(gate162inter1));
  and2  gate1123(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate1124(.a(s_82), .O(gate162inter3));
  inv1  gate1125(.a(s_83), .O(gate162inter4));
  nand2 gate1126(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate1127(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate1128(.a(G453), .O(gate162inter7));
  inv1  gate1129(.a(G534), .O(gate162inter8));
  nand2 gate1130(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate1131(.a(s_83), .b(gate162inter3), .O(gate162inter10));
  nor2  gate1132(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate1133(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate1134(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate575(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate576(.a(gate164inter0), .b(s_4), .O(gate164inter1));
  and2  gate577(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate578(.a(s_4), .O(gate164inter3));
  inv1  gate579(.a(s_5), .O(gate164inter4));
  nand2 gate580(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate581(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate582(.a(G459), .O(gate164inter7));
  inv1  gate583(.a(G537), .O(gate164inter8));
  nand2 gate584(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate585(.a(s_5), .b(gate164inter3), .O(gate164inter10));
  nor2  gate586(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate587(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate588(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );

  xor2  gate1275(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate1276(.a(gate167inter0), .b(s_104), .O(gate167inter1));
  and2  gate1277(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate1278(.a(s_104), .O(gate167inter3));
  inv1  gate1279(.a(s_105), .O(gate167inter4));
  nand2 gate1280(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate1281(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate1282(.a(G468), .O(gate167inter7));
  inv1  gate1283(.a(G543), .O(gate167inter8));
  nand2 gate1284(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate1285(.a(s_105), .b(gate167inter3), .O(gate167inter10));
  nor2  gate1286(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate1287(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate1288(.a(gate167inter12), .b(gate167inter1), .O(G584));
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate841(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate842(.a(gate198inter0), .b(s_42), .O(gate198inter1));
  and2  gate843(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate844(.a(s_42), .O(gate198inter3));
  inv1  gate845(.a(s_43), .O(gate198inter4));
  nand2 gate846(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate847(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate848(.a(G596), .O(gate198inter7));
  inv1  gate849(.a(G597), .O(gate198inter8));
  nand2 gate850(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate851(.a(s_43), .b(gate198inter3), .O(gate198inter10));
  nor2  gate852(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate853(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate854(.a(gate198inter12), .b(gate198inter1), .O(G657));
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );

  xor2  gate1387(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate1388(.a(gate209inter0), .b(s_120), .O(gate209inter1));
  and2  gate1389(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate1390(.a(s_120), .O(gate209inter3));
  inv1  gate1391(.a(s_121), .O(gate209inter4));
  nand2 gate1392(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate1393(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate1394(.a(G602), .O(gate209inter7));
  inv1  gate1395(.a(G666), .O(gate209inter8));
  nand2 gate1396(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate1397(.a(s_121), .b(gate209inter3), .O(gate209inter10));
  nor2  gate1398(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate1399(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate1400(.a(gate209inter12), .b(gate209inter1), .O(G690));
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate911(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate912(.a(gate224inter0), .b(s_52), .O(gate224inter1));
  and2  gate913(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate914(.a(s_52), .O(gate224inter3));
  inv1  gate915(.a(s_53), .O(gate224inter4));
  nand2 gate916(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate917(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate918(.a(G637), .O(gate224inter7));
  inv1  gate919(.a(G687), .O(gate224inter8));
  nand2 gate920(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate921(.a(s_53), .b(gate224inter3), .O(gate224inter10));
  nor2  gate922(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate923(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate924(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );

  xor2  gate561(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate562(.a(gate239inter0), .b(s_2), .O(gate239inter1));
  and2  gate563(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate564(.a(s_2), .O(gate239inter3));
  inv1  gate565(.a(s_3), .O(gate239inter4));
  nand2 gate566(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate567(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate568(.a(G260), .O(gate239inter7));
  inv1  gate569(.a(G712), .O(gate239inter8));
  nand2 gate570(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate571(.a(s_3), .b(gate239inter3), .O(gate239inter10));
  nor2  gate572(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate573(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate574(.a(gate239inter12), .b(gate239inter1), .O(G748));

  xor2  gate757(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate758(.a(gate240inter0), .b(s_30), .O(gate240inter1));
  and2  gate759(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate760(.a(s_30), .O(gate240inter3));
  inv1  gate761(.a(s_31), .O(gate240inter4));
  nand2 gate762(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate763(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate764(.a(G263), .O(gate240inter7));
  inv1  gate765(.a(G715), .O(gate240inter8));
  nand2 gate766(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate767(.a(s_31), .b(gate240inter3), .O(gate240inter10));
  nor2  gate768(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate769(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate770(.a(gate240inter12), .b(gate240inter1), .O(G751));

  xor2  gate1009(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate1010(.a(gate241inter0), .b(s_66), .O(gate241inter1));
  and2  gate1011(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate1012(.a(s_66), .O(gate241inter3));
  inv1  gate1013(.a(s_67), .O(gate241inter4));
  nand2 gate1014(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate1015(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate1016(.a(G242), .O(gate241inter7));
  inv1  gate1017(.a(G730), .O(gate241inter8));
  nand2 gate1018(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate1019(.a(s_67), .b(gate241inter3), .O(gate241inter10));
  nor2  gate1020(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate1021(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate1022(.a(gate241inter12), .b(gate241inter1), .O(G754));

  xor2  gate1289(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate1290(.a(gate242inter0), .b(s_106), .O(gate242inter1));
  and2  gate1291(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate1292(.a(s_106), .O(gate242inter3));
  inv1  gate1293(.a(s_107), .O(gate242inter4));
  nand2 gate1294(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate1295(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate1296(.a(G718), .O(gate242inter7));
  inv1  gate1297(.a(G730), .O(gate242inter8));
  nand2 gate1298(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate1299(.a(s_107), .b(gate242inter3), .O(gate242inter10));
  nor2  gate1300(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate1301(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate1302(.a(gate242inter12), .b(gate242inter1), .O(G755));
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate827(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate828(.a(gate250inter0), .b(s_40), .O(gate250inter1));
  and2  gate829(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate830(.a(s_40), .O(gate250inter3));
  inv1  gate831(.a(s_41), .O(gate250inter4));
  nand2 gate832(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate833(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate834(.a(G706), .O(gate250inter7));
  inv1  gate835(.a(G742), .O(gate250inter8));
  nand2 gate836(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate837(.a(s_41), .b(gate250inter3), .O(gate250inter10));
  nor2  gate838(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate839(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate840(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate1373(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate1374(.a(gate258inter0), .b(s_118), .O(gate258inter1));
  and2  gate1375(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate1376(.a(s_118), .O(gate258inter3));
  inv1  gate1377(.a(s_119), .O(gate258inter4));
  nand2 gate1378(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate1379(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate1380(.a(G756), .O(gate258inter7));
  inv1  gate1381(.a(G757), .O(gate258inter8));
  nand2 gate1382(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate1383(.a(s_119), .b(gate258inter3), .O(gate258inter10));
  nor2  gate1384(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate1385(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate1386(.a(gate258inter12), .b(gate258inter1), .O(G773));

  xor2  gate743(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate744(.a(gate259inter0), .b(s_28), .O(gate259inter1));
  and2  gate745(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate746(.a(s_28), .O(gate259inter3));
  inv1  gate747(.a(s_29), .O(gate259inter4));
  nand2 gate748(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate749(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate750(.a(G758), .O(gate259inter7));
  inv1  gate751(.a(G759), .O(gate259inter8));
  nand2 gate752(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate753(.a(s_29), .b(gate259inter3), .O(gate259inter10));
  nor2  gate754(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate755(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate756(.a(gate259inter12), .b(gate259inter1), .O(G776));
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate1303(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate1304(.a(gate271inter0), .b(s_108), .O(gate271inter1));
  and2  gate1305(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate1306(.a(s_108), .O(gate271inter3));
  inv1  gate1307(.a(s_109), .O(gate271inter4));
  nand2 gate1308(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate1309(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate1310(.a(G660), .O(gate271inter7));
  inv1  gate1311(.a(G788), .O(gate271inter8));
  nand2 gate1312(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate1313(.a(s_109), .b(gate271inter3), .O(gate271inter10));
  nor2  gate1314(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate1315(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate1316(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate869(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate870(.a(gate285inter0), .b(s_46), .O(gate285inter1));
  and2  gate871(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate872(.a(s_46), .O(gate285inter3));
  inv1  gate873(.a(s_47), .O(gate285inter4));
  nand2 gate874(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate875(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate876(.a(G660), .O(gate285inter7));
  inv1  gate877(.a(G812), .O(gate285inter8));
  nand2 gate878(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate879(.a(s_47), .b(gate285inter3), .O(gate285inter10));
  nor2  gate880(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate881(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate882(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate701(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate702(.a(gate292inter0), .b(s_22), .O(gate292inter1));
  and2  gate703(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate704(.a(s_22), .O(gate292inter3));
  inv1  gate705(.a(s_23), .O(gate292inter4));
  nand2 gate706(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate707(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate708(.a(G824), .O(gate292inter7));
  inv1  gate709(.a(G825), .O(gate292inter8));
  nand2 gate710(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate711(.a(s_23), .b(gate292inter3), .O(gate292inter10));
  nor2  gate712(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate713(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate714(.a(gate292inter12), .b(gate292inter1), .O(G873));

  xor2  gate813(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate814(.a(gate293inter0), .b(s_38), .O(gate293inter1));
  and2  gate815(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate816(.a(s_38), .O(gate293inter3));
  inv1  gate817(.a(s_39), .O(gate293inter4));
  nand2 gate818(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate819(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate820(.a(G828), .O(gate293inter7));
  inv1  gate821(.a(G829), .O(gate293inter8));
  nand2 gate822(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate823(.a(s_39), .b(gate293inter3), .O(gate293inter10));
  nor2  gate824(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate825(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate826(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate1093(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate1094(.a(gate296inter0), .b(s_78), .O(gate296inter1));
  and2  gate1095(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate1096(.a(s_78), .O(gate296inter3));
  inv1  gate1097(.a(s_79), .O(gate296inter4));
  nand2 gate1098(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate1099(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate1100(.a(G826), .O(gate296inter7));
  inv1  gate1101(.a(G827), .O(gate296inter8));
  nand2 gate1102(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate1103(.a(s_79), .b(gate296inter3), .O(gate296inter10));
  nor2  gate1104(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate1105(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate1106(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate729(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate730(.a(gate391inter0), .b(s_26), .O(gate391inter1));
  and2  gate731(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate732(.a(s_26), .O(gate391inter3));
  inv1  gate733(.a(s_27), .O(gate391inter4));
  nand2 gate734(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate735(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate736(.a(G5), .O(gate391inter7));
  inv1  gate737(.a(G1048), .O(gate391inter8));
  nand2 gate738(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate739(.a(s_27), .b(gate391inter3), .O(gate391inter10));
  nor2  gate740(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate741(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate742(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate1135(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate1136(.a(gate394inter0), .b(s_84), .O(gate394inter1));
  and2  gate1137(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate1138(.a(s_84), .O(gate394inter3));
  inv1  gate1139(.a(s_85), .O(gate394inter4));
  nand2 gate1140(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate1141(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate1142(.a(G8), .O(gate394inter7));
  inv1  gate1143(.a(G1057), .O(gate394inter8));
  nand2 gate1144(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate1145(.a(s_85), .b(gate394inter3), .O(gate394inter10));
  nor2  gate1146(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate1147(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate1148(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );

  xor2  gate897(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate898(.a(gate396inter0), .b(s_50), .O(gate396inter1));
  and2  gate899(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate900(.a(s_50), .O(gate396inter3));
  inv1  gate901(.a(s_51), .O(gate396inter4));
  nand2 gate902(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate903(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate904(.a(G10), .O(gate396inter7));
  inv1  gate905(.a(G1063), .O(gate396inter8));
  nand2 gate906(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate907(.a(s_51), .b(gate396inter3), .O(gate396inter10));
  nor2  gate908(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate909(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate910(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate1191(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate1192(.a(gate398inter0), .b(s_92), .O(gate398inter1));
  and2  gate1193(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate1194(.a(s_92), .O(gate398inter3));
  inv1  gate1195(.a(s_93), .O(gate398inter4));
  nand2 gate1196(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate1197(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate1198(.a(G12), .O(gate398inter7));
  inv1  gate1199(.a(G1069), .O(gate398inter8));
  nand2 gate1200(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate1201(.a(s_93), .b(gate398inter3), .O(gate398inter10));
  nor2  gate1202(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate1203(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate1204(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate1247(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate1248(.a(gate415inter0), .b(s_100), .O(gate415inter1));
  and2  gate1249(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate1250(.a(s_100), .O(gate415inter3));
  inv1  gate1251(.a(s_101), .O(gate415inter4));
  nand2 gate1252(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate1253(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate1254(.a(G29), .O(gate415inter7));
  inv1  gate1255(.a(G1120), .O(gate415inter8));
  nand2 gate1256(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate1257(.a(s_101), .b(gate415inter3), .O(gate415inter10));
  nor2  gate1258(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate1259(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate1260(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate799(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate800(.a(gate431inter0), .b(s_36), .O(gate431inter1));
  and2  gate801(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate802(.a(s_36), .O(gate431inter3));
  inv1  gate803(.a(s_37), .O(gate431inter4));
  nand2 gate804(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate805(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate806(.a(G7), .O(gate431inter7));
  inv1  gate807(.a(G1150), .O(gate431inter8));
  nand2 gate808(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate809(.a(s_37), .b(gate431inter3), .O(gate431inter10));
  nor2  gate810(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate811(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate812(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate1317(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate1318(.a(gate433inter0), .b(s_110), .O(gate433inter1));
  and2  gate1319(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate1320(.a(s_110), .O(gate433inter3));
  inv1  gate1321(.a(s_111), .O(gate433inter4));
  nand2 gate1322(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate1323(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate1324(.a(G8), .O(gate433inter7));
  inv1  gate1325(.a(G1153), .O(gate433inter8));
  nand2 gate1326(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate1327(.a(s_111), .b(gate433inter3), .O(gate433inter10));
  nor2  gate1328(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate1329(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate1330(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );

  xor2  gate1345(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate1346(.a(gate440inter0), .b(s_114), .O(gate440inter1));
  and2  gate1347(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate1348(.a(s_114), .O(gate440inter3));
  inv1  gate1349(.a(s_115), .O(gate440inter4));
  nand2 gate1350(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate1351(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate1352(.a(G1066), .O(gate440inter7));
  inv1  gate1353(.a(G1162), .O(gate440inter8));
  nand2 gate1354(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate1355(.a(s_115), .b(gate440inter3), .O(gate440inter10));
  nor2  gate1356(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate1357(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate1358(.a(gate440inter12), .b(gate440inter1), .O(G1249));
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );

  xor2  gate1219(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate1220(.a(gate449inter0), .b(s_96), .O(gate449inter1));
  and2  gate1221(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate1222(.a(s_96), .O(gate449inter3));
  inv1  gate1223(.a(s_97), .O(gate449inter4));
  nand2 gate1224(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate1225(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate1226(.a(G16), .O(gate449inter7));
  inv1  gate1227(.a(G1177), .O(gate449inter8));
  nand2 gate1228(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate1229(.a(s_97), .b(gate449inter3), .O(gate449inter10));
  nor2  gate1230(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate1231(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate1232(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );

  xor2  gate631(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate632(.a(gate469inter0), .b(s_12), .O(gate469inter1));
  and2  gate633(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate634(.a(s_12), .O(gate469inter3));
  inv1  gate635(.a(s_13), .O(gate469inter4));
  nand2 gate636(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate637(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate638(.a(G26), .O(gate469inter7));
  inv1  gate639(.a(G1207), .O(gate469inter8));
  nand2 gate640(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate641(.a(s_13), .b(gate469inter3), .O(gate469inter10));
  nor2  gate642(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate643(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate644(.a(gate469inter12), .b(gate469inter1), .O(G1278));
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );

  xor2  gate645(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate646(.a(gate489inter0), .b(s_14), .O(gate489inter1));
  and2  gate647(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate648(.a(s_14), .O(gate489inter3));
  inv1  gate649(.a(s_15), .O(gate489inter4));
  nand2 gate650(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate651(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate652(.a(G1240), .O(gate489inter7));
  inv1  gate653(.a(G1241), .O(gate489inter8));
  nand2 gate654(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate655(.a(s_15), .b(gate489inter3), .O(gate489inter10));
  nor2  gate656(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate657(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate658(.a(gate489inter12), .b(gate489inter1), .O(G1298));

  xor2  gate547(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate548(.a(gate490inter0), .b(s_0), .O(gate490inter1));
  and2  gate549(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate550(.a(s_0), .O(gate490inter3));
  inv1  gate551(.a(s_1), .O(gate490inter4));
  nand2 gate552(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate553(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate554(.a(G1242), .O(gate490inter7));
  inv1  gate555(.a(G1243), .O(gate490inter8));
  nand2 gate556(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate557(.a(s_1), .b(gate490inter3), .O(gate490inter10));
  nor2  gate558(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate559(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate560(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate1261(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate1262(.a(gate497inter0), .b(s_102), .O(gate497inter1));
  and2  gate1263(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate1264(.a(s_102), .O(gate497inter3));
  inv1  gate1265(.a(s_103), .O(gate497inter4));
  nand2 gate1266(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate1267(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate1268(.a(G1256), .O(gate497inter7));
  inv1  gate1269(.a(G1257), .O(gate497inter8));
  nand2 gate1270(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate1271(.a(s_103), .b(gate497inter3), .O(gate497inter10));
  nor2  gate1272(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate1273(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate1274(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate995(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate996(.a(gate501inter0), .b(s_64), .O(gate501inter1));
  and2  gate997(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate998(.a(s_64), .O(gate501inter3));
  inv1  gate999(.a(s_65), .O(gate501inter4));
  nand2 gate1000(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1001(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1002(.a(G1264), .O(gate501inter7));
  inv1  gate1003(.a(G1265), .O(gate501inter8));
  nand2 gate1004(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1005(.a(s_65), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1006(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1007(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1008(.a(gate501inter12), .b(gate501inter1), .O(G1310));

  xor2  gate1163(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate1164(.a(gate502inter0), .b(s_88), .O(gate502inter1));
  and2  gate1165(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate1166(.a(s_88), .O(gate502inter3));
  inv1  gate1167(.a(s_89), .O(gate502inter4));
  nand2 gate1168(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate1169(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate1170(.a(G1266), .O(gate502inter7));
  inv1  gate1171(.a(G1267), .O(gate502inter8));
  nand2 gate1172(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate1173(.a(s_89), .b(gate502inter3), .O(gate502inter10));
  nor2  gate1174(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate1175(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate1176(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );

  xor2  gate1233(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate1234(.a(gate507inter0), .b(s_98), .O(gate507inter1));
  and2  gate1235(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate1236(.a(s_98), .O(gate507inter3));
  inv1  gate1237(.a(s_99), .O(gate507inter4));
  nand2 gate1238(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate1239(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate1240(.a(G1276), .O(gate507inter7));
  inv1  gate1241(.a(G1277), .O(gate507inter8));
  nand2 gate1242(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate1243(.a(s_99), .b(gate507inter3), .O(gate507inter10));
  nor2  gate1244(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate1245(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate1246(.a(gate507inter12), .b(gate507inter1), .O(G1316));
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );

  xor2  gate939(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate940(.a(gate512inter0), .b(s_56), .O(gate512inter1));
  and2  gate941(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate942(.a(s_56), .O(gate512inter3));
  inv1  gate943(.a(s_57), .O(gate512inter4));
  nand2 gate944(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate945(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate946(.a(G1286), .O(gate512inter7));
  inv1  gate947(.a(G1287), .O(gate512inter8));
  nand2 gate948(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate949(.a(s_57), .b(gate512inter3), .O(gate512inter10));
  nor2  gate950(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate951(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate952(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule