module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate429inter0, gate429inter1, gate429inter2, gate429inter3, gate429inter4, gate429inter5, gate429inter6, gate429inter7, gate429inter8, gate429inter9, gate429inter10, gate429inter11, gate429inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );

  xor2  gate1541(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate1542(.a(gate14inter0), .b(s_142), .O(gate14inter1));
  and2  gate1543(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate1544(.a(s_142), .O(gate14inter3));
  inv1  gate1545(.a(s_143), .O(gate14inter4));
  nand2 gate1546(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate1547(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate1548(.a(G11), .O(gate14inter7));
  inv1  gate1549(.a(G12), .O(gate14inter8));
  nand2 gate1550(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate1551(.a(s_143), .b(gate14inter3), .O(gate14inter10));
  nor2  gate1552(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate1553(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate1554(.a(gate14inter12), .b(gate14inter1), .O(G281));

  xor2  gate561(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate562(.a(gate15inter0), .b(s_2), .O(gate15inter1));
  and2  gate563(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate564(.a(s_2), .O(gate15inter3));
  inv1  gate565(.a(s_3), .O(gate15inter4));
  nand2 gate566(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate567(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate568(.a(G13), .O(gate15inter7));
  inv1  gate569(.a(G14), .O(gate15inter8));
  nand2 gate570(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate571(.a(s_3), .b(gate15inter3), .O(gate15inter10));
  nor2  gate572(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate573(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate574(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate1821(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate1822(.a(gate19inter0), .b(s_182), .O(gate19inter1));
  and2  gate1823(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate1824(.a(s_182), .O(gate19inter3));
  inv1  gate1825(.a(s_183), .O(gate19inter4));
  nand2 gate1826(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate1827(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate1828(.a(G21), .O(gate19inter7));
  inv1  gate1829(.a(G22), .O(gate19inter8));
  nand2 gate1830(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate1831(.a(s_183), .b(gate19inter3), .O(gate19inter10));
  nor2  gate1832(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate1833(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate1834(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate1765(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate1766(.a(gate21inter0), .b(s_174), .O(gate21inter1));
  and2  gate1767(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate1768(.a(s_174), .O(gate21inter3));
  inv1  gate1769(.a(s_175), .O(gate21inter4));
  nand2 gate1770(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate1771(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate1772(.a(G25), .O(gate21inter7));
  inv1  gate1773(.a(G26), .O(gate21inter8));
  nand2 gate1774(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate1775(.a(s_175), .b(gate21inter3), .O(gate21inter10));
  nor2  gate1776(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate1777(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate1778(.a(gate21inter12), .b(gate21inter1), .O(G302));
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate743(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate744(.a(gate26inter0), .b(s_28), .O(gate26inter1));
  and2  gate745(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate746(.a(s_28), .O(gate26inter3));
  inv1  gate747(.a(s_29), .O(gate26inter4));
  nand2 gate748(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate749(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate750(.a(G9), .O(gate26inter7));
  inv1  gate751(.a(G13), .O(gate26inter8));
  nand2 gate752(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate753(.a(s_29), .b(gate26inter3), .O(gate26inter10));
  nor2  gate754(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate755(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate756(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate2059(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate2060(.a(gate36inter0), .b(s_216), .O(gate36inter1));
  and2  gate2061(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate2062(.a(s_216), .O(gate36inter3));
  inv1  gate2063(.a(s_217), .O(gate36inter4));
  nand2 gate2064(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate2065(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate2066(.a(G26), .O(gate36inter7));
  inv1  gate2067(.a(G30), .O(gate36inter8));
  nand2 gate2068(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate2069(.a(s_217), .b(gate36inter3), .O(gate36inter10));
  nor2  gate2070(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate2071(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate2072(.a(gate36inter12), .b(gate36inter1), .O(G347));

  xor2  gate981(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate982(.a(gate37inter0), .b(s_62), .O(gate37inter1));
  and2  gate983(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate984(.a(s_62), .O(gate37inter3));
  inv1  gate985(.a(s_63), .O(gate37inter4));
  nand2 gate986(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate987(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate988(.a(G19), .O(gate37inter7));
  inv1  gate989(.a(G23), .O(gate37inter8));
  nand2 gate990(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate991(.a(s_63), .b(gate37inter3), .O(gate37inter10));
  nor2  gate992(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate993(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate994(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate631(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate632(.a(gate44inter0), .b(s_12), .O(gate44inter1));
  and2  gate633(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate634(.a(s_12), .O(gate44inter3));
  inv1  gate635(.a(s_13), .O(gate44inter4));
  nand2 gate636(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate637(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate638(.a(G4), .O(gate44inter7));
  inv1  gate639(.a(G269), .O(gate44inter8));
  nand2 gate640(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate641(.a(s_13), .b(gate44inter3), .O(gate44inter10));
  nor2  gate642(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate643(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate644(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );

  xor2  gate1135(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate1136(.a(gate47inter0), .b(s_84), .O(gate47inter1));
  and2  gate1137(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate1138(.a(s_84), .O(gate47inter3));
  inv1  gate1139(.a(s_85), .O(gate47inter4));
  nand2 gate1140(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate1141(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate1142(.a(G7), .O(gate47inter7));
  inv1  gate1143(.a(G275), .O(gate47inter8));
  nand2 gate1144(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate1145(.a(s_85), .b(gate47inter3), .O(gate47inter10));
  nor2  gate1146(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate1147(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate1148(.a(gate47inter12), .b(gate47inter1), .O(G368));
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate2017(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate2018(.a(gate51inter0), .b(s_210), .O(gate51inter1));
  and2  gate2019(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate2020(.a(s_210), .O(gate51inter3));
  inv1  gate2021(.a(s_211), .O(gate51inter4));
  nand2 gate2022(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate2023(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate2024(.a(G11), .O(gate51inter7));
  inv1  gate2025(.a(G281), .O(gate51inter8));
  nand2 gate2026(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate2027(.a(s_211), .b(gate51inter3), .O(gate51inter10));
  nor2  gate2028(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate2029(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate2030(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate1877(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate1878(.a(gate54inter0), .b(s_190), .O(gate54inter1));
  and2  gate1879(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate1880(.a(s_190), .O(gate54inter3));
  inv1  gate1881(.a(s_191), .O(gate54inter4));
  nand2 gate1882(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate1883(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate1884(.a(G14), .O(gate54inter7));
  inv1  gate1885(.a(G284), .O(gate54inter8));
  nand2 gate1886(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate1887(.a(s_191), .b(gate54inter3), .O(gate54inter10));
  nor2  gate1888(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate1889(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate1890(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );

  xor2  gate1373(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate1374(.a(gate56inter0), .b(s_118), .O(gate56inter1));
  and2  gate1375(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate1376(.a(s_118), .O(gate56inter3));
  inv1  gate1377(.a(s_119), .O(gate56inter4));
  nand2 gate1378(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate1379(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate1380(.a(G16), .O(gate56inter7));
  inv1  gate1381(.a(G287), .O(gate56inter8));
  nand2 gate1382(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate1383(.a(s_119), .b(gate56inter3), .O(gate56inter10));
  nor2  gate1384(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate1385(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate1386(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );

  xor2  gate1387(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate1388(.a(gate61inter0), .b(s_120), .O(gate61inter1));
  and2  gate1389(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate1390(.a(s_120), .O(gate61inter3));
  inv1  gate1391(.a(s_121), .O(gate61inter4));
  nand2 gate1392(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate1393(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate1394(.a(G21), .O(gate61inter7));
  inv1  gate1395(.a(G296), .O(gate61inter8));
  nand2 gate1396(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate1397(.a(s_121), .b(gate61inter3), .O(gate61inter10));
  nor2  gate1398(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate1399(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate1400(.a(gate61inter12), .b(gate61inter1), .O(G382));
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );

  xor2  gate1177(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate1178(.a(gate64inter0), .b(s_90), .O(gate64inter1));
  and2  gate1179(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate1180(.a(s_90), .O(gate64inter3));
  inv1  gate1181(.a(s_91), .O(gate64inter4));
  nand2 gate1182(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate1183(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate1184(.a(G24), .O(gate64inter7));
  inv1  gate1185(.a(G299), .O(gate64inter8));
  nand2 gate1186(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate1187(.a(s_91), .b(gate64inter3), .O(gate64inter10));
  nor2  gate1188(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate1189(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate1190(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );

  xor2  gate1667(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate1668(.a(gate72inter0), .b(s_160), .O(gate72inter1));
  and2  gate1669(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate1670(.a(s_160), .O(gate72inter3));
  inv1  gate1671(.a(s_161), .O(gate72inter4));
  nand2 gate1672(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate1673(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate1674(.a(G32), .O(gate72inter7));
  inv1  gate1675(.a(G311), .O(gate72inter8));
  nand2 gate1676(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate1677(.a(s_161), .b(gate72inter3), .O(gate72inter10));
  nor2  gate1678(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate1679(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate1680(.a(gate72inter12), .b(gate72inter1), .O(G393));
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );

  xor2  gate1933(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate1934(.a(gate76inter0), .b(s_198), .O(gate76inter1));
  and2  gate1935(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate1936(.a(s_198), .O(gate76inter3));
  inv1  gate1937(.a(s_199), .O(gate76inter4));
  nand2 gate1938(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate1939(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate1940(.a(G13), .O(gate76inter7));
  inv1  gate1941(.a(G317), .O(gate76inter8));
  nand2 gate1942(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate1943(.a(s_199), .b(gate76inter3), .O(gate76inter10));
  nor2  gate1944(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate1945(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate1946(.a(gate76inter12), .b(gate76inter1), .O(G397));

  xor2  gate1905(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate1906(.a(gate77inter0), .b(s_194), .O(gate77inter1));
  and2  gate1907(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate1908(.a(s_194), .O(gate77inter3));
  inv1  gate1909(.a(s_195), .O(gate77inter4));
  nand2 gate1910(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate1911(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate1912(.a(G2), .O(gate77inter7));
  inv1  gate1913(.a(G320), .O(gate77inter8));
  nand2 gate1914(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate1915(.a(s_195), .b(gate77inter3), .O(gate77inter10));
  nor2  gate1916(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate1917(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate1918(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate2227(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate2228(.a(gate80inter0), .b(s_240), .O(gate80inter1));
  and2  gate2229(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate2230(.a(s_240), .O(gate80inter3));
  inv1  gate2231(.a(s_241), .O(gate80inter4));
  nand2 gate2232(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate2233(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate2234(.a(G14), .O(gate80inter7));
  inv1  gate2235(.a(G323), .O(gate80inter8));
  nand2 gate2236(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate2237(.a(s_241), .b(gate80inter3), .O(gate80inter10));
  nor2  gate2238(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate2239(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate2240(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate1261(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate1262(.a(gate82inter0), .b(s_102), .O(gate82inter1));
  and2  gate1263(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate1264(.a(s_102), .O(gate82inter3));
  inv1  gate1265(.a(s_103), .O(gate82inter4));
  nand2 gate1266(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate1267(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate1268(.a(G7), .O(gate82inter7));
  inv1  gate1269(.a(G326), .O(gate82inter8));
  nand2 gate1270(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate1271(.a(s_103), .b(gate82inter3), .O(gate82inter10));
  nor2  gate1272(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate1273(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate1274(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );

  xor2  gate2143(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate2144(.a(gate84inter0), .b(s_228), .O(gate84inter1));
  and2  gate2145(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate2146(.a(s_228), .O(gate84inter3));
  inv1  gate2147(.a(s_229), .O(gate84inter4));
  nand2 gate2148(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate2149(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate2150(.a(G15), .O(gate84inter7));
  inv1  gate2151(.a(G329), .O(gate84inter8));
  nand2 gate2152(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate2153(.a(s_229), .b(gate84inter3), .O(gate84inter10));
  nor2  gate2154(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate2155(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate2156(.a(gate84inter12), .b(gate84inter1), .O(G405));

  xor2  gate1695(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate1696(.a(gate85inter0), .b(s_164), .O(gate85inter1));
  and2  gate1697(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate1698(.a(s_164), .O(gate85inter3));
  inv1  gate1699(.a(s_165), .O(gate85inter4));
  nand2 gate1700(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate1701(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate1702(.a(G4), .O(gate85inter7));
  inv1  gate1703(.a(G332), .O(gate85inter8));
  nand2 gate1704(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate1705(.a(s_165), .b(gate85inter3), .O(gate85inter10));
  nor2  gate1706(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate1707(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate1708(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );

  xor2  gate1009(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate1010(.a(gate87inter0), .b(s_66), .O(gate87inter1));
  and2  gate1011(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate1012(.a(s_66), .O(gate87inter3));
  inv1  gate1013(.a(s_67), .O(gate87inter4));
  nand2 gate1014(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate1015(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate1016(.a(G12), .O(gate87inter7));
  inv1  gate1017(.a(G335), .O(gate87inter8));
  nand2 gate1018(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate1019(.a(s_67), .b(gate87inter3), .O(gate87inter10));
  nor2  gate1020(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate1021(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate1022(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate757(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate758(.a(gate90inter0), .b(s_30), .O(gate90inter1));
  and2  gate759(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate760(.a(s_30), .O(gate90inter3));
  inv1  gate761(.a(s_31), .O(gate90inter4));
  nand2 gate762(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate763(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate764(.a(G21), .O(gate90inter7));
  inv1  gate765(.a(G338), .O(gate90inter8));
  nand2 gate766(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate767(.a(s_31), .b(gate90inter3), .O(gate90inter10));
  nor2  gate768(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate769(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate770(.a(gate90inter12), .b(gate90inter1), .O(G411));

  xor2  gate547(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate548(.a(gate91inter0), .b(s_0), .O(gate91inter1));
  and2  gate549(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate550(.a(s_0), .O(gate91inter3));
  inv1  gate551(.a(s_1), .O(gate91inter4));
  nand2 gate552(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate553(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate554(.a(G25), .O(gate91inter7));
  inv1  gate555(.a(G341), .O(gate91inter8));
  nand2 gate556(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate557(.a(s_1), .b(gate91inter3), .O(gate91inter10));
  nor2  gate558(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate559(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate560(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate2199(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate2200(.a(gate94inter0), .b(s_236), .O(gate94inter1));
  and2  gate2201(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate2202(.a(s_236), .O(gate94inter3));
  inv1  gate2203(.a(s_237), .O(gate94inter4));
  nand2 gate2204(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate2205(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate2206(.a(G22), .O(gate94inter7));
  inv1  gate2207(.a(G344), .O(gate94inter8));
  nand2 gate2208(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate2209(.a(s_237), .b(gate94inter3), .O(gate94inter10));
  nor2  gate2210(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate2211(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate2212(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate2241(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate2242(.a(gate96inter0), .b(s_242), .O(gate96inter1));
  and2  gate2243(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate2244(.a(s_242), .O(gate96inter3));
  inv1  gate2245(.a(s_243), .O(gate96inter4));
  nand2 gate2246(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate2247(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate2248(.a(G30), .O(gate96inter7));
  inv1  gate2249(.a(G347), .O(gate96inter8));
  nand2 gate2250(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate2251(.a(s_243), .b(gate96inter3), .O(gate96inter10));
  nor2  gate2252(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate2253(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate2254(.a(gate96inter12), .b(gate96inter1), .O(G417));

  xor2  gate1345(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate1346(.a(gate97inter0), .b(s_114), .O(gate97inter1));
  and2  gate1347(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate1348(.a(s_114), .O(gate97inter3));
  inv1  gate1349(.a(s_115), .O(gate97inter4));
  nand2 gate1350(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate1351(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate1352(.a(G19), .O(gate97inter7));
  inv1  gate1353(.a(G350), .O(gate97inter8));
  nand2 gate1354(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate1355(.a(s_115), .b(gate97inter3), .O(gate97inter10));
  nor2  gate1356(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate1357(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate1358(.a(gate97inter12), .b(gate97inter1), .O(G418));

  xor2  gate1751(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate1752(.a(gate98inter0), .b(s_172), .O(gate98inter1));
  and2  gate1753(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate1754(.a(s_172), .O(gate98inter3));
  inv1  gate1755(.a(s_173), .O(gate98inter4));
  nand2 gate1756(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1757(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1758(.a(G23), .O(gate98inter7));
  inv1  gate1759(.a(G350), .O(gate98inter8));
  nand2 gate1760(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1761(.a(s_173), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1762(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1763(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1764(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );

  xor2  gate1471(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate1472(.a(gate101inter0), .b(s_132), .O(gate101inter1));
  and2  gate1473(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate1474(.a(s_132), .O(gate101inter3));
  inv1  gate1475(.a(s_133), .O(gate101inter4));
  nand2 gate1476(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate1477(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate1478(.a(G20), .O(gate101inter7));
  inv1  gate1479(.a(G356), .O(gate101inter8));
  nand2 gate1480(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate1481(.a(s_133), .b(gate101inter3), .O(gate101inter10));
  nor2  gate1482(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate1483(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate1484(.a(gate101inter12), .b(gate101inter1), .O(G422));

  xor2  gate1219(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate1220(.a(gate102inter0), .b(s_96), .O(gate102inter1));
  and2  gate1221(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate1222(.a(s_96), .O(gate102inter3));
  inv1  gate1223(.a(s_97), .O(gate102inter4));
  nand2 gate1224(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate1225(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate1226(.a(G24), .O(gate102inter7));
  inv1  gate1227(.a(G356), .O(gate102inter8));
  nand2 gate1228(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate1229(.a(s_97), .b(gate102inter3), .O(gate102inter10));
  nor2  gate1230(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate1231(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate1232(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate1611(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate1612(.a(gate108inter0), .b(s_152), .O(gate108inter1));
  and2  gate1613(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate1614(.a(s_152), .O(gate108inter3));
  inv1  gate1615(.a(s_153), .O(gate108inter4));
  nand2 gate1616(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate1617(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate1618(.a(G368), .O(gate108inter7));
  inv1  gate1619(.a(G369), .O(gate108inter8));
  nand2 gate1620(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate1621(.a(s_153), .b(gate108inter3), .O(gate108inter10));
  nor2  gate1622(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate1623(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate1624(.a(gate108inter12), .b(gate108inter1), .O(G435));

  xor2  gate1303(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate1304(.a(gate109inter0), .b(s_108), .O(gate109inter1));
  and2  gate1305(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate1306(.a(s_108), .O(gate109inter3));
  inv1  gate1307(.a(s_109), .O(gate109inter4));
  nand2 gate1308(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate1309(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate1310(.a(G370), .O(gate109inter7));
  inv1  gate1311(.a(G371), .O(gate109inter8));
  nand2 gate1312(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate1313(.a(s_109), .b(gate109inter3), .O(gate109inter10));
  nor2  gate1314(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate1315(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate1316(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate1919(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate1920(.a(gate117inter0), .b(s_196), .O(gate117inter1));
  and2  gate1921(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate1922(.a(s_196), .O(gate117inter3));
  inv1  gate1923(.a(s_197), .O(gate117inter4));
  nand2 gate1924(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate1925(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate1926(.a(G386), .O(gate117inter7));
  inv1  gate1927(.a(G387), .O(gate117inter8));
  nand2 gate1928(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate1929(.a(s_197), .b(gate117inter3), .O(gate117inter10));
  nor2  gate1930(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate1931(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate1932(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate1737(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate1738(.a(gate121inter0), .b(s_170), .O(gate121inter1));
  and2  gate1739(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate1740(.a(s_170), .O(gate121inter3));
  inv1  gate1741(.a(s_171), .O(gate121inter4));
  nand2 gate1742(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate1743(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate1744(.a(G394), .O(gate121inter7));
  inv1  gate1745(.a(G395), .O(gate121inter8));
  nand2 gate1746(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate1747(.a(s_171), .b(gate121inter3), .O(gate121inter10));
  nor2  gate1748(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate1749(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate1750(.a(gate121inter12), .b(gate121inter1), .O(G474));

  xor2  gate785(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate786(.a(gate122inter0), .b(s_34), .O(gate122inter1));
  and2  gate787(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate788(.a(s_34), .O(gate122inter3));
  inv1  gate789(.a(s_35), .O(gate122inter4));
  nand2 gate790(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate791(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate792(.a(G396), .O(gate122inter7));
  inv1  gate793(.a(G397), .O(gate122inter8));
  nand2 gate794(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate795(.a(s_35), .b(gate122inter3), .O(gate122inter10));
  nor2  gate796(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate797(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate798(.a(gate122inter12), .b(gate122inter1), .O(G477));

  xor2  gate1513(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate1514(.a(gate123inter0), .b(s_138), .O(gate123inter1));
  and2  gate1515(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate1516(.a(s_138), .O(gate123inter3));
  inv1  gate1517(.a(s_139), .O(gate123inter4));
  nand2 gate1518(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate1519(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate1520(.a(G398), .O(gate123inter7));
  inv1  gate1521(.a(G399), .O(gate123inter8));
  nand2 gate1522(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate1523(.a(s_139), .b(gate123inter3), .O(gate123inter10));
  nor2  gate1524(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate1525(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate1526(.a(gate123inter12), .b(gate123inter1), .O(G480));

  xor2  gate1863(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate1864(.a(gate124inter0), .b(s_188), .O(gate124inter1));
  and2  gate1865(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate1866(.a(s_188), .O(gate124inter3));
  inv1  gate1867(.a(s_189), .O(gate124inter4));
  nand2 gate1868(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate1869(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate1870(.a(G400), .O(gate124inter7));
  inv1  gate1871(.a(G401), .O(gate124inter8));
  nand2 gate1872(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate1873(.a(s_189), .b(gate124inter3), .O(gate124inter10));
  nor2  gate1874(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate1875(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate1876(.a(gate124inter12), .b(gate124inter1), .O(G483));

  xor2  gate1093(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate1094(.a(gate125inter0), .b(s_78), .O(gate125inter1));
  and2  gate1095(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate1096(.a(s_78), .O(gate125inter3));
  inv1  gate1097(.a(s_79), .O(gate125inter4));
  nand2 gate1098(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate1099(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate1100(.a(G402), .O(gate125inter7));
  inv1  gate1101(.a(G403), .O(gate125inter8));
  nand2 gate1102(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate1103(.a(s_79), .b(gate125inter3), .O(gate125inter10));
  nor2  gate1104(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate1105(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate1106(.a(gate125inter12), .b(gate125inter1), .O(G486));

  xor2  gate1849(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate1850(.a(gate126inter0), .b(s_186), .O(gate126inter1));
  and2  gate1851(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate1852(.a(s_186), .O(gate126inter3));
  inv1  gate1853(.a(s_187), .O(gate126inter4));
  nand2 gate1854(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate1855(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate1856(.a(G404), .O(gate126inter7));
  inv1  gate1857(.a(G405), .O(gate126inter8));
  nand2 gate1858(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate1859(.a(s_187), .b(gate126inter3), .O(gate126inter10));
  nor2  gate1860(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate1861(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate1862(.a(gate126inter12), .b(gate126inter1), .O(G489));

  xor2  gate1947(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate1948(.a(gate127inter0), .b(s_200), .O(gate127inter1));
  and2  gate1949(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate1950(.a(s_200), .O(gate127inter3));
  inv1  gate1951(.a(s_201), .O(gate127inter4));
  nand2 gate1952(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate1953(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate1954(.a(G406), .O(gate127inter7));
  inv1  gate1955(.a(G407), .O(gate127inter8));
  nand2 gate1956(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate1957(.a(s_201), .b(gate127inter3), .O(gate127inter10));
  nor2  gate1958(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate1959(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate1960(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate2185(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate2186(.a(gate130inter0), .b(s_234), .O(gate130inter1));
  and2  gate2187(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate2188(.a(s_234), .O(gate130inter3));
  inv1  gate2189(.a(s_235), .O(gate130inter4));
  nand2 gate2190(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate2191(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate2192(.a(G412), .O(gate130inter7));
  inv1  gate2193(.a(G413), .O(gate130inter8));
  nand2 gate2194(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate2195(.a(s_235), .b(gate130inter3), .O(gate130inter10));
  nor2  gate2196(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate2197(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate2198(.a(gate130inter12), .b(gate130inter1), .O(G501));
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );

  xor2  gate2157(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate2158(.a(gate133inter0), .b(s_230), .O(gate133inter1));
  and2  gate2159(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate2160(.a(s_230), .O(gate133inter3));
  inv1  gate2161(.a(s_231), .O(gate133inter4));
  nand2 gate2162(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate2163(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate2164(.a(G418), .O(gate133inter7));
  inv1  gate2165(.a(G419), .O(gate133inter8));
  nand2 gate2166(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate2167(.a(s_231), .b(gate133inter3), .O(gate133inter10));
  nor2  gate2168(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate2169(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate2170(.a(gate133inter12), .b(gate133inter1), .O(G510));

  xor2  gate1625(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate1626(.a(gate134inter0), .b(s_154), .O(gate134inter1));
  and2  gate1627(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate1628(.a(s_154), .O(gate134inter3));
  inv1  gate1629(.a(s_155), .O(gate134inter4));
  nand2 gate1630(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate1631(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate1632(.a(G420), .O(gate134inter7));
  inv1  gate1633(.a(G421), .O(gate134inter8));
  nand2 gate1634(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate1635(.a(s_155), .b(gate134inter3), .O(gate134inter10));
  nor2  gate1636(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate1637(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate1638(.a(gate134inter12), .b(gate134inter1), .O(G513));
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate855(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate856(.a(gate136inter0), .b(s_44), .O(gate136inter1));
  and2  gate857(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate858(.a(s_44), .O(gate136inter3));
  inv1  gate859(.a(s_45), .O(gate136inter4));
  nand2 gate860(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate861(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate862(.a(G424), .O(gate136inter7));
  inv1  gate863(.a(G425), .O(gate136inter8));
  nand2 gate864(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate865(.a(s_45), .b(gate136inter3), .O(gate136inter10));
  nor2  gate866(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate867(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate868(.a(gate136inter12), .b(gate136inter1), .O(G519));

  xor2  gate2269(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate2270(.a(gate137inter0), .b(s_246), .O(gate137inter1));
  and2  gate2271(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate2272(.a(s_246), .O(gate137inter3));
  inv1  gate2273(.a(s_247), .O(gate137inter4));
  nand2 gate2274(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate2275(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate2276(.a(G426), .O(gate137inter7));
  inv1  gate2277(.a(G429), .O(gate137inter8));
  nand2 gate2278(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate2279(.a(s_247), .b(gate137inter3), .O(gate137inter10));
  nor2  gate2280(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate2281(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate2282(.a(gate137inter12), .b(gate137inter1), .O(G522));

  xor2  gate813(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate814(.a(gate138inter0), .b(s_38), .O(gate138inter1));
  and2  gate815(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate816(.a(s_38), .O(gate138inter3));
  inv1  gate817(.a(s_39), .O(gate138inter4));
  nand2 gate818(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate819(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate820(.a(G432), .O(gate138inter7));
  inv1  gate821(.a(G435), .O(gate138inter8));
  nand2 gate822(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate823(.a(s_39), .b(gate138inter3), .O(gate138inter10));
  nor2  gate824(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate825(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate826(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate897(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate898(.a(gate142inter0), .b(s_50), .O(gate142inter1));
  and2  gate899(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate900(.a(s_50), .O(gate142inter3));
  inv1  gate901(.a(s_51), .O(gate142inter4));
  nand2 gate902(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate903(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate904(.a(G456), .O(gate142inter7));
  inv1  gate905(.a(G459), .O(gate142inter8));
  nand2 gate906(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate907(.a(s_51), .b(gate142inter3), .O(gate142inter10));
  nor2  gate908(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate909(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate910(.a(gate142inter12), .b(gate142inter1), .O(G537));
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );

  xor2  gate1779(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate1780(.a(gate145inter0), .b(s_176), .O(gate145inter1));
  and2  gate1781(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate1782(.a(s_176), .O(gate145inter3));
  inv1  gate1783(.a(s_177), .O(gate145inter4));
  nand2 gate1784(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate1785(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate1786(.a(G474), .O(gate145inter7));
  inv1  gate1787(.a(G477), .O(gate145inter8));
  nand2 gate1788(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate1789(.a(s_177), .b(gate145inter3), .O(gate145inter10));
  nor2  gate1790(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate1791(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate1792(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate995(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate996(.a(gate151inter0), .b(s_64), .O(gate151inter1));
  and2  gate997(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate998(.a(s_64), .O(gate151inter3));
  inv1  gate999(.a(s_65), .O(gate151inter4));
  nand2 gate1000(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate1001(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate1002(.a(G510), .O(gate151inter7));
  inv1  gate1003(.a(G513), .O(gate151inter8));
  nand2 gate1004(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate1005(.a(s_65), .b(gate151inter3), .O(gate151inter10));
  nor2  gate1006(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate1007(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate1008(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate2031(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate2032(.a(gate153inter0), .b(s_212), .O(gate153inter1));
  and2  gate2033(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate2034(.a(s_212), .O(gate153inter3));
  inv1  gate2035(.a(s_213), .O(gate153inter4));
  nand2 gate2036(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate2037(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate2038(.a(G426), .O(gate153inter7));
  inv1  gate2039(.a(G522), .O(gate153inter8));
  nand2 gate2040(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate2041(.a(s_213), .b(gate153inter3), .O(gate153inter10));
  nor2  gate2042(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate2043(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate2044(.a(gate153inter12), .b(gate153inter1), .O(G570));

  xor2  gate1247(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate1248(.a(gate154inter0), .b(s_100), .O(gate154inter1));
  and2  gate1249(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate1250(.a(s_100), .O(gate154inter3));
  inv1  gate1251(.a(s_101), .O(gate154inter4));
  nand2 gate1252(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate1253(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate1254(.a(G429), .O(gate154inter7));
  inv1  gate1255(.a(G522), .O(gate154inter8));
  nand2 gate1256(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate1257(.a(s_101), .b(gate154inter3), .O(gate154inter10));
  nor2  gate1258(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate1259(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate1260(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate1289(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate1290(.a(gate161inter0), .b(s_106), .O(gate161inter1));
  and2  gate1291(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate1292(.a(s_106), .O(gate161inter3));
  inv1  gate1293(.a(s_107), .O(gate161inter4));
  nand2 gate1294(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate1295(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate1296(.a(G450), .O(gate161inter7));
  inv1  gate1297(.a(G534), .O(gate161inter8));
  nand2 gate1298(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate1299(.a(s_107), .b(gate161inter3), .O(gate161inter10));
  nor2  gate1300(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate1301(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate1302(.a(gate161inter12), .b(gate161inter1), .O(G578));

  xor2  gate1457(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate1458(.a(gate162inter0), .b(s_130), .O(gate162inter1));
  and2  gate1459(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate1460(.a(s_130), .O(gate162inter3));
  inv1  gate1461(.a(s_131), .O(gate162inter4));
  nand2 gate1462(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate1463(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate1464(.a(G453), .O(gate162inter7));
  inv1  gate1465(.a(G534), .O(gate162inter8));
  nand2 gate1466(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate1467(.a(s_131), .b(gate162inter3), .O(gate162inter10));
  nor2  gate1468(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate1469(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate1470(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );

  xor2  gate589(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate590(.a(gate166inter0), .b(s_6), .O(gate166inter1));
  and2  gate591(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate592(.a(s_6), .O(gate166inter3));
  inv1  gate593(.a(s_7), .O(gate166inter4));
  nand2 gate594(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate595(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate596(.a(G465), .O(gate166inter7));
  inv1  gate597(.a(G540), .O(gate166inter8));
  nand2 gate598(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate599(.a(s_7), .b(gate166inter3), .O(gate166inter10));
  nor2  gate600(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate601(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate602(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate1037(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate1038(.a(gate174inter0), .b(s_70), .O(gate174inter1));
  and2  gate1039(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate1040(.a(s_70), .O(gate174inter3));
  inv1  gate1041(.a(s_71), .O(gate174inter4));
  nand2 gate1042(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate1043(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate1044(.a(G489), .O(gate174inter7));
  inv1  gate1045(.a(G552), .O(gate174inter8));
  nand2 gate1046(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate1047(.a(s_71), .b(gate174inter3), .O(gate174inter10));
  nor2  gate1048(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate1049(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate1050(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );

  xor2  gate939(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate940(.a(gate176inter0), .b(s_56), .O(gate176inter1));
  and2  gate941(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate942(.a(s_56), .O(gate176inter3));
  inv1  gate943(.a(s_57), .O(gate176inter4));
  nand2 gate944(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate945(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate946(.a(G495), .O(gate176inter7));
  inv1  gate947(.a(G555), .O(gate176inter8));
  nand2 gate948(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate949(.a(s_57), .b(gate176inter3), .O(gate176inter10));
  nor2  gate950(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate951(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate952(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate2283(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate2284(.a(gate180inter0), .b(s_248), .O(gate180inter1));
  and2  gate2285(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate2286(.a(s_248), .O(gate180inter3));
  inv1  gate2287(.a(s_249), .O(gate180inter4));
  nand2 gate2288(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate2289(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate2290(.a(G507), .O(gate180inter7));
  inv1  gate2291(.a(G561), .O(gate180inter8));
  nand2 gate2292(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate2293(.a(s_249), .b(gate180inter3), .O(gate180inter10));
  nor2  gate2294(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate2295(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate2296(.a(gate180inter12), .b(gate180inter1), .O(G597));
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate1107(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1108(.a(gate186inter0), .b(s_80), .O(gate186inter1));
  and2  gate1109(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1110(.a(s_80), .O(gate186inter3));
  inv1  gate1111(.a(s_81), .O(gate186inter4));
  nand2 gate1112(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1113(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1114(.a(G572), .O(gate186inter7));
  inv1  gate1115(.a(G573), .O(gate186inter8));
  nand2 gate1116(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1117(.a(s_81), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1118(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1119(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1120(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate1485(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate1486(.a(gate195inter0), .b(s_134), .O(gate195inter1));
  and2  gate1487(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate1488(.a(s_134), .O(gate195inter3));
  inv1  gate1489(.a(s_135), .O(gate195inter4));
  nand2 gate1490(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate1491(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate1492(.a(G590), .O(gate195inter7));
  inv1  gate1493(.a(G591), .O(gate195inter8));
  nand2 gate1494(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate1495(.a(s_135), .b(gate195inter3), .O(gate195inter10));
  nor2  gate1496(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate1497(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate1498(.a(gate195inter12), .b(gate195inter1), .O(G648));

  xor2  gate673(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate674(.a(gate196inter0), .b(s_18), .O(gate196inter1));
  and2  gate675(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate676(.a(s_18), .O(gate196inter3));
  inv1  gate677(.a(s_19), .O(gate196inter4));
  nand2 gate678(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate679(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate680(.a(G592), .O(gate196inter7));
  inv1  gate681(.a(G593), .O(gate196inter8));
  nand2 gate682(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate683(.a(s_19), .b(gate196inter3), .O(gate196inter10));
  nor2  gate684(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate685(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate686(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate1401(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate1402(.a(gate198inter0), .b(s_122), .O(gate198inter1));
  and2  gate1403(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate1404(.a(s_122), .O(gate198inter3));
  inv1  gate1405(.a(s_123), .O(gate198inter4));
  nand2 gate1406(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate1407(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate1408(.a(G596), .O(gate198inter7));
  inv1  gate1409(.a(G597), .O(gate198inter8));
  nand2 gate1410(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate1411(.a(s_123), .b(gate198inter3), .O(gate198inter10));
  nor2  gate1412(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate1413(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate1414(.a(gate198inter12), .b(gate198inter1), .O(G657));

  xor2  gate799(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate800(.a(gate199inter0), .b(s_36), .O(gate199inter1));
  and2  gate801(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate802(.a(s_36), .O(gate199inter3));
  inv1  gate803(.a(s_37), .O(gate199inter4));
  nand2 gate804(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate805(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate806(.a(G598), .O(gate199inter7));
  inv1  gate807(.a(G599), .O(gate199inter8));
  nand2 gate808(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate809(.a(s_37), .b(gate199inter3), .O(gate199inter10));
  nor2  gate810(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate811(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate812(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate869(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate870(.a(gate203inter0), .b(s_46), .O(gate203inter1));
  and2  gate871(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate872(.a(s_46), .O(gate203inter3));
  inv1  gate873(.a(s_47), .O(gate203inter4));
  nand2 gate874(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate875(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate876(.a(G602), .O(gate203inter7));
  inv1  gate877(.a(G612), .O(gate203inter8));
  nand2 gate878(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate879(.a(s_47), .b(gate203inter3), .O(gate203inter10));
  nor2  gate880(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate881(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate882(.a(gate203inter12), .b(gate203inter1), .O(G672));

  xor2  gate2115(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate2116(.a(gate204inter0), .b(s_224), .O(gate204inter1));
  and2  gate2117(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate2118(.a(s_224), .O(gate204inter3));
  inv1  gate2119(.a(s_225), .O(gate204inter4));
  nand2 gate2120(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate2121(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate2122(.a(G607), .O(gate204inter7));
  inv1  gate2123(.a(G617), .O(gate204inter8));
  nand2 gate2124(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate2125(.a(s_225), .b(gate204inter3), .O(gate204inter10));
  nor2  gate2126(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate2127(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate2128(.a(gate204inter12), .b(gate204inter1), .O(G675));
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );

  xor2  gate2129(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate2130(.a(gate207inter0), .b(s_226), .O(gate207inter1));
  and2  gate2131(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate2132(.a(s_226), .O(gate207inter3));
  inv1  gate2133(.a(s_227), .O(gate207inter4));
  nand2 gate2134(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate2135(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate2136(.a(G622), .O(gate207inter7));
  inv1  gate2137(.a(G632), .O(gate207inter8));
  nand2 gate2138(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate2139(.a(s_227), .b(gate207inter3), .O(gate207inter10));
  nor2  gate2140(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate2141(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate2142(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );

  xor2  gate1793(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate1794(.a(gate209inter0), .b(s_178), .O(gate209inter1));
  and2  gate1795(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate1796(.a(s_178), .O(gate209inter3));
  inv1  gate1797(.a(s_179), .O(gate209inter4));
  nand2 gate1798(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate1799(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate1800(.a(G602), .O(gate209inter7));
  inv1  gate1801(.a(G666), .O(gate209inter8));
  nand2 gate1802(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate1803(.a(s_179), .b(gate209inter3), .O(gate209inter10));
  nor2  gate1804(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate1805(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate1806(.a(gate209inter12), .b(gate209inter1), .O(G690));
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );

  xor2  gate953(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate954(.a(gate212inter0), .b(s_58), .O(gate212inter1));
  and2  gate955(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate956(.a(s_58), .O(gate212inter3));
  inv1  gate957(.a(s_59), .O(gate212inter4));
  nand2 gate958(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate959(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate960(.a(G617), .O(gate212inter7));
  inv1  gate961(.a(G669), .O(gate212inter8));
  nand2 gate962(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate963(.a(s_59), .b(gate212inter3), .O(gate212inter10));
  nor2  gate964(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate965(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate966(.a(gate212inter12), .b(gate212inter1), .O(G693));

  xor2  gate2297(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate2298(.a(gate213inter0), .b(s_250), .O(gate213inter1));
  and2  gate2299(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate2300(.a(s_250), .O(gate213inter3));
  inv1  gate2301(.a(s_251), .O(gate213inter4));
  nand2 gate2302(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate2303(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate2304(.a(G602), .O(gate213inter7));
  inv1  gate2305(.a(G672), .O(gate213inter8));
  nand2 gate2306(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate2307(.a(s_251), .b(gate213inter3), .O(gate213inter10));
  nor2  gate2308(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate2309(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate2310(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate2171(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate2172(.a(gate215inter0), .b(s_232), .O(gate215inter1));
  and2  gate2173(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate2174(.a(s_232), .O(gate215inter3));
  inv1  gate2175(.a(s_233), .O(gate215inter4));
  nand2 gate2176(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate2177(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate2178(.a(G607), .O(gate215inter7));
  inv1  gate2179(.a(G675), .O(gate215inter8));
  nand2 gate2180(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate2181(.a(s_233), .b(gate215inter3), .O(gate215inter10));
  nor2  gate2182(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate2183(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate2184(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate1975(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate1976(.a(gate223inter0), .b(s_204), .O(gate223inter1));
  and2  gate1977(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate1978(.a(s_204), .O(gate223inter3));
  inv1  gate1979(.a(s_205), .O(gate223inter4));
  nand2 gate1980(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate1981(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate1982(.a(G627), .O(gate223inter7));
  inv1  gate1983(.a(G687), .O(gate223inter8));
  nand2 gate1984(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate1985(.a(s_205), .b(gate223inter3), .O(gate223inter10));
  nor2  gate1986(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate1987(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate1988(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate841(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate842(.a(gate227inter0), .b(s_42), .O(gate227inter1));
  and2  gate843(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate844(.a(s_42), .O(gate227inter3));
  inv1  gate845(.a(s_43), .O(gate227inter4));
  nand2 gate846(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate847(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate848(.a(G694), .O(gate227inter7));
  inv1  gate849(.a(G695), .O(gate227inter8));
  nand2 gate850(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate851(.a(s_43), .b(gate227inter3), .O(gate227inter10));
  nor2  gate852(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate853(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate854(.a(gate227inter12), .b(gate227inter1), .O(G712));

  xor2  gate1527(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate1528(.a(gate228inter0), .b(s_140), .O(gate228inter1));
  and2  gate1529(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate1530(.a(s_140), .O(gate228inter3));
  inv1  gate1531(.a(s_141), .O(gate228inter4));
  nand2 gate1532(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate1533(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate1534(.a(G696), .O(gate228inter7));
  inv1  gate1535(.a(G697), .O(gate228inter8));
  nand2 gate1536(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate1537(.a(s_141), .b(gate228inter3), .O(gate228inter10));
  nor2  gate1538(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate1539(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate1540(.a(gate228inter12), .b(gate228inter1), .O(G715));

  xor2  gate1681(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate1682(.a(gate229inter0), .b(s_162), .O(gate229inter1));
  and2  gate1683(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate1684(.a(s_162), .O(gate229inter3));
  inv1  gate1685(.a(s_163), .O(gate229inter4));
  nand2 gate1686(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate1687(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate1688(.a(G698), .O(gate229inter7));
  inv1  gate1689(.a(G699), .O(gate229inter8));
  nand2 gate1690(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate1691(.a(s_163), .b(gate229inter3), .O(gate229inter10));
  nor2  gate1692(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate1693(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate1694(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );

  xor2  gate617(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate618(.a(gate232inter0), .b(s_10), .O(gate232inter1));
  and2  gate619(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate620(.a(s_10), .O(gate232inter3));
  inv1  gate621(.a(s_11), .O(gate232inter4));
  nand2 gate622(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate623(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate624(.a(G704), .O(gate232inter7));
  inv1  gate625(.a(G705), .O(gate232inter8));
  nand2 gate626(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate627(.a(s_11), .b(gate232inter3), .O(gate232inter10));
  nor2  gate628(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate629(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate630(.a(gate232inter12), .b(gate232inter1), .O(G727));
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate2101(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate2102(.a(gate234inter0), .b(s_222), .O(gate234inter1));
  and2  gate2103(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate2104(.a(s_222), .O(gate234inter3));
  inv1  gate2105(.a(s_223), .O(gate234inter4));
  nand2 gate2106(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate2107(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate2108(.a(G245), .O(gate234inter7));
  inv1  gate2109(.a(G721), .O(gate234inter8));
  nand2 gate2110(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate2111(.a(s_223), .b(gate234inter3), .O(gate234inter10));
  nor2  gate2112(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate2113(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate2114(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate1569(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate1570(.a(gate236inter0), .b(s_146), .O(gate236inter1));
  and2  gate1571(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate1572(.a(s_146), .O(gate236inter3));
  inv1  gate1573(.a(s_147), .O(gate236inter4));
  nand2 gate1574(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate1575(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate1576(.a(G251), .O(gate236inter7));
  inv1  gate1577(.a(G727), .O(gate236inter8));
  nand2 gate1578(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate1579(.a(s_147), .b(gate236inter3), .O(gate236inter10));
  nor2  gate1580(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate1581(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate1582(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );

  xor2  gate883(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate884(.a(gate239inter0), .b(s_48), .O(gate239inter1));
  and2  gate885(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate886(.a(s_48), .O(gate239inter3));
  inv1  gate887(.a(s_49), .O(gate239inter4));
  nand2 gate888(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate889(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate890(.a(G260), .O(gate239inter7));
  inv1  gate891(.a(G712), .O(gate239inter8));
  nand2 gate892(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate893(.a(s_49), .b(gate239inter3), .O(gate239inter10));
  nor2  gate894(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate895(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate896(.a(gate239inter12), .b(gate239inter1), .O(G748));

  xor2  gate967(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate968(.a(gate240inter0), .b(s_60), .O(gate240inter1));
  and2  gate969(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate970(.a(s_60), .O(gate240inter3));
  inv1  gate971(.a(s_61), .O(gate240inter4));
  nand2 gate972(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate973(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate974(.a(G263), .O(gate240inter7));
  inv1  gate975(.a(G715), .O(gate240inter8));
  nand2 gate976(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate977(.a(s_61), .b(gate240inter3), .O(gate240inter10));
  nor2  gate978(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate979(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate980(.a(gate240inter12), .b(gate240inter1), .O(G751));

  xor2  gate2073(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate2074(.a(gate241inter0), .b(s_218), .O(gate241inter1));
  and2  gate2075(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate2076(.a(s_218), .O(gate241inter3));
  inv1  gate2077(.a(s_219), .O(gate241inter4));
  nand2 gate2078(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate2079(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate2080(.a(G242), .O(gate241inter7));
  inv1  gate2081(.a(G730), .O(gate241inter8));
  nand2 gate2082(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate2083(.a(s_219), .b(gate241inter3), .O(gate241inter10));
  nor2  gate2084(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate2085(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate2086(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate1639(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate1640(.a(gate248inter0), .b(s_156), .O(gate248inter1));
  and2  gate1641(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate1642(.a(s_156), .O(gate248inter3));
  inv1  gate1643(.a(s_157), .O(gate248inter4));
  nand2 gate1644(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate1645(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate1646(.a(G727), .O(gate248inter7));
  inv1  gate1647(.a(G739), .O(gate248inter8));
  nand2 gate1648(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate1649(.a(s_157), .b(gate248inter3), .O(gate248inter10));
  nor2  gate1650(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate1651(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate1652(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );

  xor2  gate1709(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate1710(.a(gate251inter0), .b(s_166), .O(gate251inter1));
  and2  gate1711(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate1712(.a(s_166), .O(gate251inter3));
  inv1  gate1713(.a(s_167), .O(gate251inter4));
  nand2 gate1714(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate1715(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate1716(.a(G257), .O(gate251inter7));
  inv1  gate1717(.a(G745), .O(gate251inter8));
  nand2 gate1718(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate1719(.a(s_167), .b(gate251inter3), .O(gate251inter10));
  nor2  gate1720(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate1721(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate1722(.a(gate251inter12), .b(gate251inter1), .O(G764));
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate2045(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate2046(.a(gate253inter0), .b(s_214), .O(gate253inter1));
  and2  gate2047(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate2048(.a(s_214), .O(gate253inter3));
  inv1  gate2049(.a(s_215), .O(gate253inter4));
  nand2 gate2050(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate2051(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate2052(.a(G260), .O(gate253inter7));
  inv1  gate2053(.a(G748), .O(gate253inter8));
  nand2 gate2054(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate2055(.a(s_215), .b(gate253inter3), .O(gate253inter10));
  nor2  gate2056(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate2057(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate2058(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate1233(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate1234(.a(gate256inter0), .b(s_98), .O(gate256inter1));
  and2  gate1235(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate1236(.a(s_98), .O(gate256inter3));
  inv1  gate1237(.a(s_99), .O(gate256inter4));
  nand2 gate1238(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate1239(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate1240(.a(G715), .O(gate256inter7));
  inv1  gate1241(.a(G751), .O(gate256inter8));
  nand2 gate1242(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate1243(.a(s_99), .b(gate256inter3), .O(gate256inter10));
  nor2  gate1244(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate1245(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate1246(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate1807(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate1808(.a(gate262inter0), .b(s_180), .O(gate262inter1));
  and2  gate1809(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate1810(.a(s_180), .O(gate262inter3));
  inv1  gate1811(.a(s_181), .O(gate262inter4));
  nand2 gate1812(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate1813(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate1814(.a(G764), .O(gate262inter7));
  inv1  gate1815(.a(G765), .O(gate262inter8));
  nand2 gate1816(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate1817(.a(s_181), .b(gate262inter3), .O(gate262inter10));
  nor2  gate1818(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate1819(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate1820(.a(gate262inter12), .b(gate262inter1), .O(G785));

  xor2  gate827(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate828(.a(gate263inter0), .b(s_40), .O(gate263inter1));
  and2  gate829(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate830(.a(s_40), .O(gate263inter3));
  inv1  gate831(.a(s_41), .O(gate263inter4));
  nand2 gate832(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate833(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate834(.a(G766), .O(gate263inter7));
  inv1  gate835(.a(G767), .O(gate263inter8));
  nand2 gate836(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate837(.a(s_41), .b(gate263inter3), .O(gate263inter10));
  nor2  gate838(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate839(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate840(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate1443(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate1444(.a(gate266inter0), .b(s_128), .O(gate266inter1));
  and2  gate1445(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate1446(.a(s_128), .O(gate266inter3));
  inv1  gate1447(.a(s_129), .O(gate266inter4));
  nand2 gate1448(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate1449(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate1450(.a(G645), .O(gate266inter7));
  inv1  gate1451(.a(G773), .O(gate266inter8));
  nand2 gate1452(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate1453(.a(s_129), .b(gate266inter3), .O(gate266inter10));
  nor2  gate1454(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate1455(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate1456(.a(gate266inter12), .b(gate266inter1), .O(G797));

  xor2  gate2213(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate2214(.a(gate267inter0), .b(s_238), .O(gate267inter1));
  and2  gate2215(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate2216(.a(s_238), .O(gate267inter3));
  inv1  gate2217(.a(s_239), .O(gate267inter4));
  nand2 gate2218(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate2219(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate2220(.a(G648), .O(gate267inter7));
  inv1  gate2221(.a(G776), .O(gate267inter8));
  nand2 gate2222(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate2223(.a(s_239), .b(gate267inter3), .O(gate267inter10));
  nor2  gate2224(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate2225(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate2226(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate1989(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate1990(.a(gate279inter0), .b(s_206), .O(gate279inter1));
  and2  gate1991(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate1992(.a(s_206), .O(gate279inter3));
  inv1  gate1993(.a(s_207), .O(gate279inter4));
  nand2 gate1994(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate1995(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate1996(.a(G651), .O(gate279inter7));
  inv1  gate1997(.a(G803), .O(gate279inter8));
  nand2 gate1998(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate1999(.a(s_207), .b(gate279inter3), .O(gate279inter10));
  nor2  gate2000(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate2001(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate2002(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );

  xor2  gate715(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate716(.a(gate284inter0), .b(s_24), .O(gate284inter1));
  and2  gate717(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate718(.a(s_24), .O(gate284inter3));
  inv1  gate719(.a(s_25), .O(gate284inter4));
  nand2 gate720(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate721(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate722(.a(G785), .O(gate284inter7));
  inv1  gate723(.a(G809), .O(gate284inter8));
  nand2 gate724(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate725(.a(s_25), .b(gate284inter3), .O(gate284inter10));
  nor2  gate726(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate727(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate728(.a(gate284inter12), .b(gate284inter1), .O(G829));
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate1835(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate1836(.a(gate286inter0), .b(s_184), .O(gate286inter1));
  and2  gate1837(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate1838(.a(s_184), .O(gate286inter3));
  inv1  gate1839(.a(s_185), .O(gate286inter4));
  nand2 gate1840(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate1841(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate1842(.a(G788), .O(gate286inter7));
  inv1  gate1843(.a(G812), .O(gate286inter8));
  nand2 gate1844(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate1845(.a(s_185), .b(gate286inter3), .O(gate286inter10));
  nor2  gate1846(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate1847(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate1848(.a(gate286inter12), .b(gate286inter1), .O(G831));
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate1317(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate1318(.a(gate292inter0), .b(s_110), .O(gate292inter1));
  and2  gate1319(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate1320(.a(s_110), .O(gate292inter3));
  inv1  gate1321(.a(s_111), .O(gate292inter4));
  nand2 gate1322(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate1323(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate1324(.a(G824), .O(gate292inter7));
  inv1  gate1325(.a(G825), .O(gate292inter8));
  nand2 gate1326(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate1327(.a(s_111), .b(gate292inter3), .O(gate292inter10));
  nor2  gate1328(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate1329(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate1330(.a(gate292inter12), .b(gate292inter1), .O(G873));

  xor2  gate1079(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate1080(.a(gate293inter0), .b(s_76), .O(gate293inter1));
  and2  gate1081(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate1082(.a(s_76), .O(gate293inter3));
  inv1  gate1083(.a(s_77), .O(gate293inter4));
  nand2 gate1084(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate1085(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate1086(.a(G828), .O(gate293inter7));
  inv1  gate1087(.a(G829), .O(gate293inter8));
  nand2 gate1088(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate1089(.a(s_77), .b(gate293inter3), .O(gate293inter10));
  nor2  gate1090(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate1091(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate1092(.a(gate293inter12), .b(gate293inter1), .O(G886));

  xor2  gate1065(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate1066(.a(gate294inter0), .b(s_74), .O(gate294inter1));
  and2  gate1067(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate1068(.a(s_74), .O(gate294inter3));
  inv1  gate1069(.a(s_75), .O(gate294inter4));
  nand2 gate1070(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate1071(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate1072(.a(G832), .O(gate294inter7));
  inv1  gate1073(.a(G833), .O(gate294inter8));
  nand2 gate1074(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate1075(.a(s_75), .b(gate294inter3), .O(gate294inter10));
  nor2  gate1076(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate1077(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate1078(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );

  xor2  gate687(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate688(.a(gate396inter0), .b(s_20), .O(gate396inter1));
  and2  gate689(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate690(.a(s_20), .O(gate396inter3));
  inv1  gate691(.a(s_21), .O(gate396inter4));
  nand2 gate692(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate693(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate694(.a(G10), .O(gate396inter7));
  inv1  gate695(.a(G1063), .O(gate396inter8));
  nand2 gate696(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate697(.a(s_21), .b(gate396inter3), .O(gate396inter10));
  nor2  gate698(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate699(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate700(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate729(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate730(.a(gate399inter0), .b(s_26), .O(gate399inter1));
  and2  gate731(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate732(.a(s_26), .O(gate399inter3));
  inv1  gate733(.a(s_27), .O(gate399inter4));
  nand2 gate734(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate735(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate736(.a(G13), .O(gate399inter7));
  inv1  gate737(.a(G1072), .O(gate399inter8));
  nand2 gate738(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate739(.a(s_27), .b(gate399inter3), .O(gate399inter10));
  nor2  gate740(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate741(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate742(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );

  xor2  gate2255(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate2256(.a(gate402inter0), .b(s_244), .O(gate402inter1));
  and2  gate2257(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate2258(.a(s_244), .O(gate402inter3));
  inv1  gate2259(.a(s_245), .O(gate402inter4));
  nand2 gate2260(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate2261(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate2262(.a(G16), .O(gate402inter7));
  inv1  gate2263(.a(G1081), .O(gate402inter8));
  nand2 gate2264(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate2265(.a(s_245), .b(gate402inter3), .O(gate402inter10));
  nor2  gate2266(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate2267(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate2268(.a(gate402inter12), .b(gate402inter1), .O(G1177));
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate1205(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate1206(.a(gate417inter0), .b(s_94), .O(gate417inter1));
  and2  gate1207(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate1208(.a(s_94), .O(gate417inter3));
  inv1  gate1209(.a(s_95), .O(gate417inter4));
  nand2 gate1210(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate1211(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate1212(.a(G31), .O(gate417inter7));
  inv1  gate1213(.a(G1126), .O(gate417inter8));
  nand2 gate1214(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate1215(.a(s_95), .b(gate417inter3), .O(gate417inter10));
  nor2  gate1216(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate1217(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate1218(.a(gate417inter12), .b(gate417inter1), .O(G1222));

  xor2  gate575(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate576(.a(gate418inter0), .b(s_4), .O(gate418inter1));
  and2  gate577(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate578(.a(s_4), .O(gate418inter3));
  inv1  gate579(.a(s_5), .O(gate418inter4));
  nand2 gate580(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate581(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate582(.a(G32), .O(gate418inter7));
  inv1  gate583(.a(G1129), .O(gate418inter8));
  nand2 gate584(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate585(.a(s_5), .b(gate418inter3), .O(gate418inter10));
  nor2  gate586(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate587(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate588(.a(gate418inter12), .b(gate418inter1), .O(G1225));

  xor2  gate1583(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate1584(.a(gate419inter0), .b(s_148), .O(gate419inter1));
  and2  gate1585(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate1586(.a(s_148), .O(gate419inter3));
  inv1  gate1587(.a(s_149), .O(gate419inter4));
  nand2 gate1588(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate1589(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate1590(.a(G1), .O(gate419inter7));
  inv1  gate1591(.a(G1132), .O(gate419inter8));
  nand2 gate1592(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate1593(.a(s_149), .b(gate419inter3), .O(gate419inter10));
  nor2  gate1594(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate1595(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate1596(.a(gate419inter12), .b(gate419inter1), .O(G1228));

  xor2  gate1597(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1598(.a(gate420inter0), .b(s_150), .O(gate420inter1));
  and2  gate1599(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1600(.a(s_150), .O(gate420inter3));
  inv1  gate1601(.a(s_151), .O(gate420inter4));
  nand2 gate1602(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1603(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1604(.a(G1036), .O(gate420inter7));
  inv1  gate1605(.a(G1132), .O(gate420inter8));
  nand2 gate1606(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1607(.a(s_151), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1608(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1609(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1610(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );

  xor2  gate1891(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate1892(.a(gate423inter0), .b(s_192), .O(gate423inter1));
  and2  gate1893(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate1894(.a(s_192), .O(gate423inter3));
  inv1  gate1895(.a(s_193), .O(gate423inter4));
  nand2 gate1896(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate1897(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate1898(.a(G3), .O(gate423inter7));
  inv1  gate1899(.a(G1138), .O(gate423inter8));
  nand2 gate1900(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate1901(.a(s_193), .b(gate423inter3), .O(gate423inter10));
  nor2  gate1902(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate1903(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate1904(.a(gate423inter12), .b(gate423inter1), .O(G1232));
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );

  xor2  gate645(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate646(.a(gate427inter0), .b(s_14), .O(gate427inter1));
  and2  gate647(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate648(.a(s_14), .O(gate427inter3));
  inv1  gate649(.a(s_15), .O(gate427inter4));
  nand2 gate650(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate651(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate652(.a(G5), .O(gate427inter7));
  inv1  gate653(.a(G1144), .O(gate427inter8));
  nand2 gate654(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate655(.a(s_15), .b(gate427inter3), .O(gate427inter10));
  nor2  gate656(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate657(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate658(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );

  xor2  gate1051(.a(G1147), .b(G6), .O(gate429inter0));
  nand2 gate1052(.a(gate429inter0), .b(s_72), .O(gate429inter1));
  and2  gate1053(.a(G1147), .b(G6), .O(gate429inter2));
  inv1  gate1054(.a(s_72), .O(gate429inter3));
  inv1  gate1055(.a(s_73), .O(gate429inter4));
  nand2 gate1056(.a(gate429inter4), .b(gate429inter3), .O(gate429inter5));
  nor2  gate1057(.a(gate429inter5), .b(gate429inter2), .O(gate429inter6));
  inv1  gate1058(.a(G6), .O(gate429inter7));
  inv1  gate1059(.a(G1147), .O(gate429inter8));
  nand2 gate1060(.a(gate429inter8), .b(gate429inter7), .O(gate429inter9));
  nand2 gate1061(.a(s_73), .b(gate429inter3), .O(gate429inter10));
  nor2  gate1062(.a(gate429inter10), .b(gate429inter9), .O(gate429inter11));
  nor2  gate1063(.a(gate429inter11), .b(gate429inter6), .O(gate429inter12));
  nand2 gate1064(.a(gate429inter12), .b(gate429inter1), .O(G1238));
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate1653(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate1654(.a(gate433inter0), .b(s_158), .O(gate433inter1));
  and2  gate1655(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate1656(.a(s_158), .O(gate433inter3));
  inv1  gate1657(.a(s_159), .O(gate433inter4));
  nand2 gate1658(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate1659(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate1660(.a(G8), .O(gate433inter7));
  inv1  gate1661(.a(G1153), .O(gate433inter8));
  nand2 gate1662(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate1663(.a(s_159), .b(gate433inter3), .O(gate433inter10));
  nor2  gate1664(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate1665(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate1666(.a(gate433inter12), .b(gate433inter1), .O(G1242));

  xor2  gate1149(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate1150(.a(gate434inter0), .b(s_86), .O(gate434inter1));
  and2  gate1151(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate1152(.a(s_86), .O(gate434inter3));
  inv1  gate1153(.a(s_87), .O(gate434inter4));
  nand2 gate1154(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate1155(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate1156(.a(G1057), .O(gate434inter7));
  inv1  gate1157(.a(G1153), .O(gate434inter8));
  nand2 gate1158(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate1159(.a(s_87), .b(gate434inter3), .O(gate434inter10));
  nor2  gate1160(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate1161(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate1162(.a(gate434inter12), .b(gate434inter1), .O(G1243));

  xor2  gate2003(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate2004(.a(gate435inter0), .b(s_208), .O(gate435inter1));
  and2  gate2005(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate2006(.a(s_208), .O(gate435inter3));
  inv1  gate2007(.a(s_209), .O(gate435inter4));
  nand2 gate2008(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate2009(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate2010(.a(G9), .O(gate435inter7));
  inv1  gate2011(.a(G1156), .O(gate435inter8));
  nand2 gate2012(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate2013(.a(s_209), .b(gate435inter3), .O(gate435inter10));
  nor2  gate2014(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate2015(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate2016(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate1359(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate1360(.a(gate438inter0), .b(s_116), .O(gate438inter1));
  and2  gate1361(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate1362(.a(s_116), .O(gate438inter3));
  inv1  gate1363(.a(s_117), .O(gate438inter4));
  nand2 gate1364(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate1365(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate1366(.a(G1063), .O(gate438inter7));
  inv1  gate1367(.a(G1159), .O(gate438inter8));
  nand2 gate1368(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate1369(.a(s_117), .b(gate438inter3), .O(gate438inter10));
  nor2  gate1370(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate1371(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate1372(.a(gate438inter12), .b(gate438inter1), .O(G1247));

  xor2  gate771(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate772(.a(gate439inter0), .b(s_32), .O(gate439inter1));
  and2  gate773(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate774(.a(s_32), .O(gate439inter3));
  inv1  gate775(.a(s_33), .O(gate439inter4));
  nand2 gate776(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate777(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate778(.a(G11), .O(gate439inter7));
  inv1  gate779(.a(G1162), .O(gate439inter8));
  nand2 gate780(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate781(.a(s_33), .b(gate439inter3), .O(gate439inter10));
  nor2  gate782(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate783(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate784(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate2087(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate2088(.a(gate444inter0), .b(s_220), .O(gate444inter1));
  and2  gate2089(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate2090(.a(s_220), .O(gate444inter3));
  inv1  gate2091(.a(s_221), .O(gate444inter4));
  nand2 gate2092(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate2093(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate2094(.a(G1072), .O(gate444inter7));
  inv1  gate2095(.a(G1168), .O(gate444inter8));
  nand2 gate2096(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate2097(.a(s_221), .b(gate444inter3), .O(gate444inter10));
  nor2  gate2098(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate2099(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate2100(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate1121(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate1122(.a(gate456inter0), .b(s_82), .O(gate456inter1));
  and2  gate1123(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate1124(.a(s_82), .O(gate456inter3));
  inv1  gate1125(.a(s_83), .O(gate456inter4));
  nand2 gate1126(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate1127(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate1128(.a(G1090), .O(gate456inter7));
  inv1  gate1129(.a(G1186), .O(gate456inter8));
  nand2 gate1130(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate1131(.a(s_83), .b(gate456inter3), .O(gate456inter10));
  nor2  gate1132(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate1133(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate1134(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );

  xor2  gate911(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate912(.a(gate458inter0), .b(s_52), .O(gate458inter1));
  and2  gate913(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate914(.a(s_52), .O(gate458inter3));
  inv1  gate915(.a(s_53), .O(gate458inter4));
  nand2 gate916(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate917(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate918(.a(G1093), .O(gate458inter7));
  inv1  gate919(.a(G1189), .O(gate458inter8));
  nand2 gate920(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate921(.a(s_53), .b(gate458inter3), .O(gate458inter10));
  nor2  gate922(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate923(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate924(.a(gate458inter12), .b(gate458inter1), .O(G1267));
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate1163(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate1164(.a(gate464inter0), .b(s_88), .O(gate464inter1));
  and2  gate1165(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate1166(.a(s_88), .O(gate464inter3));
  inv1  gate1167(.a(s_89), .O(gate464inter4));
  nand2 gate1168(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate1169(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate1170(.a(G1102), .O(gate464inter7));
  inv1  gate1171(.a(G1198), .O(gate464inter8));
  nand2 gate1172(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate1173(.a(s_89), .b(gate464inter3), .O(gate464inter10));
  nor2  gate1174(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate1175(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate1176(.a(gate464inter12), .b(gate464inter1), .O(G1273));

  xor2  gate701(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate702(.a(gate465inter0), .b(s_22), .O(gate465inter1));
  and2  gate703(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate704(.a(s_22), .O(gate465inter3));
  inv1  gate705(.a(s_23), .O(gate465inter4));
  nand2 gate706(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate707(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate708(.a(G24), .O(gate465inter7));
  inv1  gate709(.a(G1201), .O(gate465inter8));
  nand2 gate710(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate711(.a(s_23), .b(gate465inter3), .O(gate465inter10));
  nor2  gate712(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate713(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate714(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate1331(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate1332(.a(gate475inter0), .b(s_112), .O(gate475inter1));
  and2  gate1333(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate1334(.a(s_112), .O(gate475inter3));
  inv1  gate1335(.a(s_113), .O(gate475inter4));
  nand2 gate1336(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate1337(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate1338(.a(G29), .O(gate475inter7));
  inv1  gate1339(.a(G1216), .O(gate475inter8));
  nand2 gate1340(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate1341(.a(s_113), .b(gate475inter3), .O(gate475inter10));
  nor2  gate1342(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate1343(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate1344(.a(gate475inter12), .b(gate475inter1), .O(G1284));
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );

  xor2  gate603(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate604(.a(gate479inter0), .b(s_8), .O(gate479inter1));
  and2  gate605(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate606(.a(s_8), .O(gate479inter3));
  inv1  gate607(.a(s_9), .O(gate479inter4));
  nand2 gate608(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate609(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate610(.a(G31), .O(gate479inter7));
  inv1  gate611(.a(G1222), .O(gate479inter8));
  nand2 gate612(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate613(.a(s_9), .b(gate479inter3), .O(gate479inter10));
  nor2  gate614(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate615(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate616(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );

  xor2  gate925(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate926(.a(gate483inter0), .b(s_54), .O(gate483inter1));
  and2  gate927(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate928(.a(s_54), .O(gate483inter3));
  inv1  gate929(.a(s_55), .O(gate483inter4));
  nand2 gate930(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate931(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate932(.a(G1228), .O(gate483inter7));
  inv1  gate933(.a(G1229), .O(gate483inter8));
  nand2 gate934(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate935(.a(s_55), .b(gate483inter3), .O(gate483inter10));
  nor2  gate936(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate937(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate938(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate1555(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate1556(.a(gate486inter0), .b(s_144), .O(gate486inter1));
  and2  gate1557(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate1558(.a(s_144), .O(gate486inter3));
  inv1  gate1559(.a(s_145), .O(gate486inter4));
  nand2 gate1560(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate1561(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate1562(.a(G1234), .O(gate486inter7));
  inv1  gate1563(.a(G1235), .O(gate486inter8));
  nand2 gate1564(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate1565(.a(s_145), .b(gate486inter3), .O(gate486inter10));
  nor2  gate1566(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate1567(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate1568(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate1023(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate1024(.a(gate488inter0), .b(s_68), .O(gate488inter1));
  and2  gate1025(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate1026(.a(s_68), .O(gate488inter3));
  inv1  gate1027(.a(s_69), .O(gate488inter4));
  nand2 gate1028(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate1029(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate1030(.a(G1238), .O(gate488inter7));
  inv1  gate1031(.a(G1239), .O(gate488inter8));
  nand2 gate1032(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate1033(.a(s_69), .b(gate488inter3), .O(gate488inter10));
  nor2  gate1034(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate1035(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate1036(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate1191(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate1192(.a(gate490inter0), .b(s_92), .O(gate490inter1));
  and2  gate1193(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate1194(.a(s_92), .O(gate490inter3));
  inv1  gate1195(.a(s_93), .O(gate490inter4));
  nand2 gate1196(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate1197(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate1198(.a(G1242), .O(gate490inter7));
  inv1  gate1199(.a(G1243), .O(gate490inter8));
  nand2 gate1200(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate1201(.a(s_93), .b(gate490inter3), .O(gate490inter10));
  nor2  gate1202(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate1203(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate1204(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate659(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate660(.a(gate492inter0), .b(s_16), .O(gate492inter1));
  and2  gate661(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate662(.a(s_16), .O(gate492inter3));
  inv1  gate663(.a(s_17), .O(gate492inter4));
  nand2 gate664(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate665(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate666(.a(G1246), .O(gate492inter7));
  inv1  gate667(.a(G1247), .O(gate492inter8));
  nand2 gate668(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate669(.a(s_17), .b(gate492inter3), .O(gate492inter10));
  nor2  gate670(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate671(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate672(.a(gate492inter12), .b(gate492inter1), .O(G1301));

  xor2  gate1429(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate1430(.a(gate493inter0), .b(s_126), .O(gate493inter1));
  and2  gate1431(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate1432(.a(s_126), .O(gate493inter3));
  inv1  gate1433(.a(s_127), .O(gate493inter4));
  nand2 gate1434(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate1435(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate1436(.a(G1248), .O(gate493inter7));
  inv1  gate1437(.a(G1249), .O(gate493inter8));
  nand2 gate1438(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate1439(.a(s_127), .b(gate493inter3), .O(gate493inter10));
  nor2  gate1440(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate1441(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate1442(.a(gate493inter12), .b(gate493inter1), .O(G1302));
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );

  xor2  gate1275(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate1276(.a(gate495inter0), .b(s_104), .O(gate495inter1));
  and2  gate1277(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate1278(.a(s_104), .O(gate495inter3));
  inv1  gate1279(.a(s_105), .O(gate495inter4));
  nand2 gate1280(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate1281(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate1282(.a(G1252), .O(gate495inter7));
  inv1  gate1283(.a(G1253), .O(gate495inter8));
  nand2 gate1284(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate1285(.a(s_105), .b(gate495inter3), .O(gate495inter10));
  nor2  gate1286(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate1287(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate1288(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate1961(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate1962(.a(gate500inter0), .b(s_202), .O(gate500inter1));
  and2  gate1963(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate1964(.a(s_202), .O(gate500inter3));
  inv1  gate1965(.a(s_203), .O(gate500inter4));
  nand2 gate1966(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate1967(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate1968(.a(G1262), .O(gate500inter7));
  inv1  gate1969(.a(G1263), .O(gate500inter8));
  nand2 gate1970(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate1971(.a(s_203), .b(gate500inter3), .O(gate500inter10));
  nor2  gate1972(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate1973(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate1974(.a(gate500inter12), .b(gate500inter1), .O(G1309));
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );

  xor2  gate1723(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate1724(.a(gate507inter0), .b(s_168), .O(gate507inter1));
  and2  gate1725(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate1726(.a(s_168), .O(gate507inter3));
  inv1  gate1727(.a(s_169), .O(gate507inter4));
  nand2 gate1728(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate1729(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate1730(.a(G1276), .O(gate507inter7));
  inv1  gate1731(.a(G1277), .O(gate507inter8));
  nand2 gate1732(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate1733(.a(s_169), .b(gate507inter3), .O(gate507inter10));
  nor2  gate1734(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate1735(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate1736(.a(gate507inter12), .b(gate507inter1), .O(G1316));

  xor2  gate1415(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate1416(.a(gate508inter0), .b(s_124), .O(gate508inter1));
  and2  gate1417(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate1418(.a(s_124), .O(gate508inter3));
  inv1  gate1419(.a(s_125), .O(gate508inter4));
  nand2 gate1420(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate1421(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate1422(.a(G1278), .O(gate508inter7));
  inv1  gate1423(.a(G1279), .O(gate508inter8));
  nand2 gate1424(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate1425(.a(s_125), .b(gate508inter3), .O(gate508inter10));
  nor2  gate1426(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate1427(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate1428(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate1499(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate1500(.a(gate511inter0), .b(s_136), .O(gate511inter1));
  and2  gate1501(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate1502(.a(s_136), .O(gate511inter3));
  inv1  gate1503(.a(s_137), .O(gate511inter4));
  nand2 gate1504(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate1505(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate1506(.a(G1284), .O(gate511inter7));
  inv1  gate1507(.a(G1285), .O(gate511inter8));
  nand2 gate1508(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate1509(.a(s_137), .b(gate511inter3), .O(gate511inter10));
  nor2  gate1510(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate1511(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate1512(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule