module c499 (N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
             N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
             N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
             N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
             N137,N724,N725,N726,N727,N728,N729,N730,N731,N732,
             N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,
             N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,
             N753,N754,N755);
input N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
      N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
      N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
      N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
      N137;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51;
output N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,
       N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
       N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
       N754,N755;
wire N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
     N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
     N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,
     N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,
     N290,N293,N296,N299,N302,N305,N308,N311,N314,N315,
     N316,N317,N318,N319,N320,N321,N338,N339,N340,N341,
     N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,
     N352,N353,N354,N367,N380,N393,N406,N419,N432,N445,
     N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
     N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,
     N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,
     N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,
     N594,N595,N596,N597,N598,N599,N600,N601,N602,N607,
     N620,N625,N630,N635,N640,N645,N650,N655,N692,N693,
     N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,
     N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,
     N714,N715,N716,N717,N718,N719,N720,N721,N722,N723, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate3inter0, gate3inter1, gate3inter2, gate3inter3, gate3inter4, gate3inter5, gate3inter6, gate3inter7, gate3inter8, gate3inter9, gate3inter10, gate3inter11, gate3inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12;


xor2 gate1( .a(N1), .b(N5), .O(N250) );
xor2 gate2( .a(N9), .b(N13), .O(N251) );

  xor2  gate259(.a(N21), .b(N17), .O(gate3inter0));
  nand2 gate260(.a(gate3inter0), .b(s_8), .O(gate3inter1));
  and2  gate261(.a(N21), .b(N17), .O(gate3inter2));
  inv1  gate262(.a(s_8), .O(gate3inter3));
  inv1  gate263(.a(s_9), .O(gate3inter4));
  nand2 gate264(.a(gate3inter4), .b(gate3inter3), .O(gate3inter5));
  nor2  gate265(.a(gate3inter5), .b(gate3inter2), .O(gate3inter6));
  inv1  gate266(.a(N17), .O(gate3inter7));
  inv1  gate267(.a(N21), .O(gate3inter8));
  nand2 gate268(.a(gate3inter8), .b(gate3inter7), .O(gate3inter9));
  nand2 gate269(.a(s_9), .b(gate3inter3), .O(gate3inter10));
  nor2  gate270(.a(gate3inter10), .b(gate3inter9), .O(gate3inter11));
  nor2  gate271(.a(gate3inter11), .b(gate3inter6), .O(gate3inter12));
  nand2 gate272(.a(gate3inter12), .b(gate3inter1), .O(N252));
xor2 gate4( .a(N25), .b(N29), .O(N253) );
xor2 gate5( .a(N33), .b(N37), .O(N254) );
xor2 gate6( .a(N41), .b(N45), .O(N255) );
xor2 gate7( .a(N49), .b(N53), .O(N256) );
xor2 gate8( .a(N57), .b(N61), .O(N257) );

  xor2  gate343(.a(N69), .b(N65), .O(gate9inter0));
  nand2 gate344(.a(gate9inter0), .b(s_20), .O(gate9inter1));
  and2  gate345(.a(N69), .b(N65), .O(gate9inter2));
  inv1  gate346(.a(s_20), .O(gate9inter3));
  inv1  gate347(.a(s_21), .O(gate9inter4));
  nand2 gate348(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate349(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate350(.a(N65), .O(gate9inter7));
  inv1  gate351(.a(N69), .O(gate9inter8));
  nand2 gate352(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate353(.a(s_21), .b(gate9inter3), .O(gate9inter10));
  nor2  gate354(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate355(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate356(.a(gate9inter12), .b(gate9inter1), .O(N258));
xor2 gate10( .a(N73), .b(N77), .O(N259) );
xor2 gate11( .a(N81), .b(N85), .O(N260) );

  xor2  gate497(.a(N93), .b(N89), .O(gate12inter0));
  nand2 gate498(.a(gate12inter0), .b(s_42), .O(gate12inter1));
  and2  gate499(.a(N93), .b(N89), .O(gate12inter2));
  inv1  gate500(.a(s_42), .O(gate12inter3));
  inv1  gate501(.a(s_43), .O(gate12inter4));
  nand2 gate502(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate503(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate504(.a(N89), .O(gate12inter7));
  inv1  gate505(.a(N93), .O(gate12inter8));
  nand2 gate506(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate507(.a(s_43), .b(gate12inter3), .O(gate12inter10));
  nor2  gate508(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate509(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate510(.a(gate12inter12), .b(gate12inter1), .O(N261));
xor2 gate13( .a(N97), .b(N101), .O(N262) );
xor2 gate14( .a(N105), .b(N109), .O(N263) );
xor2 gate15( .a(N113), .b(N117), .O(N264) );
xor2 gate16( .a(N121), .b(N125), .O(N265) );
and2 gate17( .a(N129), .b(N137), .O(N266) );
and2 gate18( .a(N130), .b(N137), .O(N267) );
and2 gate19( .a(N131), .b(N137), .O(N268) );
and2 gate20( .a(N132), .b(N137), .O(N269) );
and2 gate21( .a(N133), .b(N137), .O(N270) );
and2 gate22( .a(N134), .b(N137), .O(N271) );
and2 gate23( .a(N135), .b(N137), .O(N272) );
and2 gate24( .a(N136), .b(N137), .O(N273) );
xor2 gate25( .a(N1), .b(N17), .O(N274) );
xor2 gate26( .a(N33), .b(N49), .O(N275) );
xor2 gate27( .a(N5), .b(N21), .O(N276) );
xor2 gate28( .a(N37), .b(N53), .O(N277) );
xor2 gate29( .a(N9), .b(N25), .O(N278) );
xor2 gate30( .a(N41), .b(N57), .O(N279) );
xor2 gate31( .a(N13), .b(N29), .O(N280) );

  xor2  gate329(.a(N61), .b(N45), .O(gate32inter0));
  nand2 gate330(.a(gate32inter0), .b(s_18), .O(gate32inter1));
  and2  gate331(.a(N61), .b(N45), .O(gate32inter2));
  inv1  gate332(.a(s_18), .O(gate32inter3));
  inv1  gate333(.a(s_19), .O(gate32inter4));
  nand2 gate334(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate335(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate336(.a(N45), .O(gate32inter7));
  inv1  gate337(.a(N61), .O(gate32inter8));
  nand2 gate338(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate339(.a(s_19), .b(gate32inter3), .O(gate32inter10));
  nor2  gate340(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate341(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate342(.a(gate32inter12), .b(gate32inter1), .O(N281));
xor2 gate33( .a(N65), .b(N81), .O(N282) );
xor2 gate34( .a(N97), .b(N113), .O(N283) );
xor2 gate35( .a(N69), .b(N85), .O(N284) );
xor2 gate36( .a(N101), .b(N117), .O(N285) );

  xor2  gate483(.a(N89), .b(N73), .O(gate37inter0));
  nand2 gate484(.a(gate37inter0), .b(s_40), .O(gate37inter1));
  and2  gate485(.a(N89), .b(N73), .O(gate37inter2));
  inv1  gate486(.a(s_40), .O(gate37inter3));
  inv1  gate487(.a(s_41), .O(gate37inter4));
  nand2 gate488(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate489(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate490(.a(N73), .O(gate37inter7));
  inv1  gate491(.a(N89), .O(gate37inter8));
  nand2 gate492(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate493(.a(s_41), .b(gate37inter3), .O(gate37inter10));
  nor2  gate494(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate495(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate496(.a(gate37inter12), .b(gate37inter1), .O(N286));

  xor2  gate203(.a(N121), .b(N105), .O(gate38inter0));
  nand2 gate204(.a(gate38inter0), .b(s_0), .O(gate38inter1));
  and2  gate205(.a(N121), .b(N105), .O(gate38inter2));
  inv1  gate206(.a(s_0), .O(gate38inter3));
  inv1  gate207(.a(s_1), .O(gate38inter4));
  nand2 gate208(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate209(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate210(.a(N105), .O(gate38inter7));
  inv1  gate211(.a(N121), .O(gate38inter8));
  nand2 gate212(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate213(.a(s_1), .b(gate38inter3), .O(gate38inter10));
  nor2  gate214(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate215(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate216(.a(gate38inter12), .b(gate38inter1), .O(N287));
xor2 gate39( .a(N77), .b(N93), .O(N288) );
xor2 gate40( .a(N109), .b(N125), .O(N289) );
xor2 gate41( .a(N250), .b(N251), .O(N290) );
xor2 gate42( .a(N252), .b(N253), .O(N293) );
xor2 gate43( .a(N254), .b(N255), .O(N296) );
xor2 gate44( .a(N256), .b(N257), .O(N299) );
xor2 gate45( .a(N258), .b(N259), .O(N302) );
xor2 gate46( .a(N260), .b(N261), .O(N305) );
xor2 gate47( .a(N262), .b(N263), .O(N308) );
xor2 gate48( .a(N264), .b(N265), .O(N311) );

  xor2  gate553(.a(N275), .b(N274), .O(gate49inter0));
  nand2 gate554(.a(gate49inter0), .b(s_50), .O(gate49inter1));
  and2  gate555(.a(N275), .b(N274), .O(gate49inter2));
  inv1  gate556(.a(s_50), .O(gate49inter3));
  inv1  gate557(.a(s_51), .O(gate49inter4));
  nand2 gate558(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate559(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate560(.a(N274), .O(gate49inter7));
  inv1  gate561(.a(N275), .O(gate49inter8));
  nand2 gate562(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate563(.a(s_51), .b(gate49inter3), .O(gate49inter10));
  nor2  gate564(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate565(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate566(.a(gate49inter12), .b(gate49inter1), .O(N314));
xor2 gate50( .a(N276), .b(N277), .O(N315) );

  xor2  gate441(.a(N279), .b(N278), .O(gate51inter0));
  nand2 gate442(.a(gate51inter0), .b(s_34), .O(gate51inter1));
  and2  gate443(.a(N279), .b(N278), .O(gate51inter2));
  inv1  gate444(.a(s_34), .O(gate51inter3));
  inv1  gate445(.a(s_35), .O(gate51inter4));
  nand2 gate446(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate447(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate448(.a(N278), .O(gate51inter7));
  inv1  gate449(.a(N279), .O(gate51inter8));
  nand2 gate450(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate451(.a(s_35), .b(gate51inter3), .O(gate51inter10));
  nor2  gate452(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate453(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate454(.a(gate51inter12), .b(gate51inter1), .O(N316));
xor2 gate52( .a(N280), .b(N281), .O(N317) );
xor2 gate53( .a(N282), .b(N283), .O(N318) );
xor2 gate54( .a(N284), .b(N285), .O(N319) );

  xor2  gate413(.a(N287), .b(N286), .O(gate55inter0));
  nand2 gate414(.a(gate55inter0), .b(s_30), .O(gate55inter1));
  and2  gate415(.a(N287), .b(N286), .O(gate55inter2));
  inv1  gate416(.a(s_30), .O(gate55inter3));
  inv1  gate417(.a(s_31), .O(gate55inter4));
  nand2 gate418(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate419(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate420(.a(N286), .O(gate55inter7));
  inv1  gate421(.a(N287), .O(gate55inter8));
  nand2 gate422(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate423(.a(s_31), .b(gate55inter3), .O(gate55inter10));
  nor2  gate424(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate425(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate426(.a(gate55inter12), .b(gate55inter1), .O(N320));
xor2 gate56( .a(N288), .b(N289), .O(N321) );
xor2 gate57( .a(N290), .b(N293), .O(N338) );
xor2 gate58( .a(N296), .b(N299), .O(N339) );
xor2 gate59( .a(N290), .b(N296), .O(N340) );
xor2 gate60( .a(N293), .b(N299), .O(N341) );

  xor2  gate371(.a(N305), .b(N302), .O(gate61inter0));
  nand2 gate372(.a(gate61inter0), .b(s_24), .O(gate61inter1));
  and2  gate373(.a(N305), .b(N302), .O(gate61inter2));
  inv1  gate374(.a(s_24), .O(gate61inter3));
  inv1  gate375(.a(s_25), .O(gate61inter4));
  nand2 gate376(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate377(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate378(.a(N302), .O(gate61inter7));
  inv1  gate379(.a(N305), .O(gate61inter8));
  nand2 gate380(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate381(.a(s_25), .b(gate61inter3), .O(gate61inter10));
  nor2  gate382(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate383(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate384(.a(gate61inter12), .b(gate61inter1), .O(N342));
xor2 gate62( .a(N308), .b(N311), .O(N343) );

  xor2  gate245(.a(N308), .b(N302), .O(gate63inter0));
  nand2 gate246(.a(gate63inter0), .b(s_6), .O(gate63inter1));
  and2  gate247(.a(N308), .b(N302), .O(gate63inter2));
  inv1  gate248(.a(s_6), .O(gate63inter3));
  inv1  gate249(.a(s_7), .O(gate63inter4));
  nand2 gate250(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate251(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate252(.a(N302), .O(gate63inter7));
  inv1  gate253(.a(N308), .O(gate63inter8));
  nand2 gate254(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate255(.a(s_7), .b(gate63inter3), .O(gate63inter10));
  nor2  gate256(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate257(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate258(.a(gate63inter12), .b(gate63inter1), .O(N344));
xor2 gate64( .a(N305), .b(N311), .O(N345) );
xor2 gate65( .a(N266), .b(N342), .O(N346) );
xor2 gate66( .a(N267), .b(N343), .O(N347) );

  xor2  gate455(.a(N344), .b(N268), .O(gate67inter0));
  nand2 gate456(.a(gate67inter0), .b(s_36), .O(gate67inter1));
  and2  gate457(.a(N344), .b(N268), .O(gate67inter2));
  inv1  gate458(.a(s_36), .O(gate67inter3));
  inv1  gate459(.a(s_37), .O(gate67inter4));
  nand2 gate460(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate461(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate462(.a(N268), .O(gate67inter7));
  inv1  gate463(.a(N344), .O(gate67inter8));
  nand2 gate464(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate465(.a(s_37), .b(gate67inter3), .O(gate67inter10));
  nor2  gate466(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate467(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate468(.a(gate67inter12), .b(gate67inter1), .O(N348));
xor2 gate68( .a(N269), .b(N345), .O(N349) );
xor2 gate69( .a(N270), .b(N338), .O(N350) );
xor2 gate70( .a(N271), .b(N339), .O(N351) );
xor2 gate71( .a(N272), .b(N340), .O(N352) );

  xor2  gate511(.a(N341), .b(N273), .O(gate72inter0));
  nand2 gate512(.a(gate72inter0), .b(s_44), .O(gate72inter1));
  and2  gate513(.a(N341), .b(N273), .O(gate72inter2));
  inv1  gate514(.a(s_44), .O(gate72inter3));
  inv1  gate515(.a(s_45), .O(gate72inter4));
  nand2 gate516(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate517(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate518(.a(N273), .O(gate72inter7));
  inv1  gate519(.a(N341), .O(gate72inter8));
  nand2 gate520(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate521(.a(s_45), .b(gate72inter3), .O(gate72inter10));
  nor2  gate522(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate523(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate524(.a(gate72inter12), .b(gate72inter1), .O(N353));
xor2 gate73( .a(N314), .b(N346), .O(N354) );
xor2 gate74( .a(N315), .b(N347), .O(N367) );

  xor2  gate357(.a(N348), .b(N316), .O(gate75inter0));
  nand2 gate358(.a(gate75inter0), .b(s_22), .O(gate75inter1));
  and2  gate359(.a(N348), .b(N316), .O(gate75inter2));
  inv1  gate360(.a(s_22), .O(gate75inter3));
  inv1  gate361(.a(s_23), .O(gate75inter4));
  nand2 gate362(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate363(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate364(.a(N316), .O(gate75inter7));
  inv1  gate365(.a(N348), .O(gate75inter8));
  nand2 gate366(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate367(.a(s_23), .b(gate75inter3), .O(gate75inter10));
  nor2  gate368(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate369(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate370(.a(gate75inter12), .b(gate75inter1), .O(N380));

  xor2  gate525(.a(N349), .b(N317), .O(gate76inter0));
  nand2 gate526(.a(gate76inter0), .b(s_46), .O(gate76inter1));
  and2  gate527(.a(N349), .b(N317), .O(gate76inter2));
  inv1  gate528(.a(s_46), .O(gate76inter3));
  inv1  gate529(.a(s_47), .O(gate76inter4));
  nand2 gate530(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate531(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate532(.a(N317), .O(gate76inter7));
  inv1  gate533(.a(N349), .O(gate76inter8));
  nand2 gate534(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate535(.a(s_47), .b(gate76inter3), .O(gate76inter10));
  nor2  gate536(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate537(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate538(.a(gate76inter12), .b(gate76inter1), .O(N393));

  xor2  gate231(.a(N350), .b(N318), .O(gate77inter0));
  nand2 gate232(.a(gate77inter0), .b(s_4), .O(gate77inter1));
  and2  gate233(.a(N350), .b(N318), .O(gate77inter2));
  inv1  gate234(.a(s_4), .O(gate77inter3));
  inv1  gate235(.a(s_5), .O(gate77inter4));
  nand2 gate236(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate237(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate238(.a(N318), .O(gate77inter7));
  inv1  gate239(.a(N350), .O(gate77inter8));
  nand2 gate240(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate241(.a(s_5), .b(gate77inter3), .O(gate77inter10));
  nor2  gate242(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate243(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate244(.a(gate77inter12), .b(gate77inter1), .O(N406));

  xor2  gate469(.a(N351), .b(N319), .O(gate78inter0));
  nand2 gate470(.a(gate78inter0), .b(s_38), .O(gate78inter1));
  and2  gate471(.a(N351), .b(N319), .O(gate78inter2));
  inv1  gate472(.a(s_38), .O(gate78inter3));
  inv1  gate473(.a(s_39), .O(gate78inter4));
  nand2 gate474(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate475(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate476(.a(N319), .O(gate78inter7));
  inv1  gate477(.a(N351), .O(gate78inter8));
  nand2 gate478(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate479(.a(s_39), .b(gate78inter3), .O(gate78inter10));
  nor2  gate480(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate481(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate482(.a(gate78inter12), .b(gate78inter1), .O(N419));
xor2 gate79( .a(N320), .b(N352), .O(N432) );

  xor2  gate287(.a(N353), .b(N321), .O(gate80inter0));
  nand2 gate288(.a(gate80inter0), .b(s_12), .O(gate80inter1));
  and2  gate289(.a(N353), .b(N321), .O(gate80inter2));
  inv1  gate290(.a(s_12), .O(gate80inter3));
  inv1  gate291(.a(s_13), .O(gate80inter4));
  nand2 gate292(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate293(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate294(.a(N321), .O(gate80inter7));
  inv1  gate295(.a(N353), .O(gate80inter8));
  nand2 gate296(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate297(.a(s_13), .b(gate80inter3), .O(gate80inter10));
  nor2  gate298(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate299(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate300(.a(gate80inter12), .b(gate80inter1), .O(N445));
inv1 gate81( .a(N354), .O(N554) );
inv1 gate82( .a(N367), .O(N555) );
inv1 gate83( .a(N380), .O(N556) );
inv1 gate84( .a(N354), .O(N557) );
inv1 gate85( .a(N367), .O(N558) );
inv1 gate86( .a(N393), .O(N559) );
inv1 gate87( .a(N354), .O(N560) );
inv1 gate88( .a(N380), .O(N561) );
inv1 gate89( .a(N393), .O(N562) );
inv1 gate90( .a(N367), .O(N563) );
inv1 gate91( .a(N380), .O(N564) );
inv1 gate92( .a(N393), .O(N565) );
inv1 gate93( .a(N419), .O(N566) );
inv1 gate94( .a(N445), .O(N567) );
inv1 gate95( .a(N419), .O(N568) );
inv1 gate96( .a(N432), .O(N569) );
inv1 gate97( .a(N406), .O(N570) );
inv1 gate98( .a(N445), .O(N571) );
inv1 gate99( .a(N406), .O(N572) );
inv1 gate100( .a(N432), .O(N573) );
inv1 gate101( .a(N406), .O(N574) );
inv1 gate102( .a(N419), .O(N575) );
inv1 gate103( .a(N432), .O(N576) );
inv1 gate104( .a(N406), .O(N577) );
inv1 gate105( .a(N419), .O(N578) );
inv1 gate106( .a(N445), .O(N579) );
inv1 gate107( .a(N406), .O(N580) );
inv1 gate108( .a(N432), .O(N581) );
inv1 gate109( .a(N445), .O(N582) );
inv1 gate110( .a(N419), .O(N583) );
inv1 gate111( .a(N432), .O(N584) );
inv1 gate112( .a(N445), .O(N585) );
inv1 gate113( .a(N367), .O(N586) );
inv1 gate114( .a(N393), .O(N587) );
inv1 gate115( .a(N367), .O(N588) );
inv1 gate116( .a(N380), .O(N589) );
inv1 gate117( .a(N354), .O(N590) );
inv1 gate118( .a(N393), .O(N591) );
inv1 gate119( .a(N354), .O(N592) );
inv1 gate120( .a(N380), .O(N593) );
and4 gate121( .a(N554), .b(N555), .c(N556), .d(N393), .O(N594) );
and4 gate122( .a(N557), .b(N558), .c(N380), .d(N559), .O(N595) );
and4 gate123( .a(N560), .b(N367), .c(N561), .d(N562), .O(N596) );
and4 gate124( .a(N354), .b(N563), .c(N564), .d(N565), .O(N597) );
and4 gate125( .a(N574), .b(N575), .c(N576), .d(N445), .O(N598) );
and4 gate126( .a(N577), .b(N578), .c(N432), .d(N579), .O(N599) );
and4 gate127( .a(N580), .b(N419), .c(N581), .d(N582), .O(N600) );
and4 gate128( .a(N406), .b(N583), .c(N584), .d(N585), .O(N601) );
or4 gate129( .a(N594), .b(N595), .c(N596), .d(N597), .O(N602) );
or4 gate130( .a(N598), .b(N599), .c(N600), .d(N601), .O(N607) );
and5 gate131( .a(N406), .b(N566), .c(N432), .d(N567), .e(N602), .O(N620) );
and5 gate132( .a(N406), .b(N568), .c(N569), .d(N445), .e(N602), .O(N625) );
and5 gate133( .a(N570), .b(N419), .c(N432), .d(N571), .e(N602), .O(N630) );
and5 gate134( .a(N572), .b(N419), .c(N573), .d(N445), .e(N602), .O(N635) );
and5 gate135( .a(N354), .b(N586), .c(N380), .d(N587), .e(N607), .O(N640) );
and5 gate136( .a(N354), .b(N588), .c(N589), .d(N393), .e(N607), .O(N645) );
and5 gate137( .a(N590), .b(N367), .c(N380), .d(N591), .e(N607), .O(N650) );
and5 gate138( .a(N592), .b(N367), .c(N593), .d(N393), .e(N607), .O(N655) );
and2 gate139( .a(N354), .b(N620), .O(N692) );
and2 gate140( .a(N367), .b(N620), .O(N693) );
and2 gate141( .a(N380), .b(N620), .O(N694) );
and2 gate142( .a(N393), .b(N620), .O(N695) );
and2 gate143( .a(N354), .b(N625), .O(N696) );
and2 gate144( .a(N367), .b(N625), .O(N697) );
and2 gate145( .a(N380), .b(N625), .O(N698) );
and2 gate146( .a(N393), .b(N625), .O(N699) );
and2 gate147( .a(N354), .b(N630), .O(N700) );
and2 gate148( .a(N367), .b(N630), .O(N701) );
and2 gate149( .a(N380), .b(N630), .O(N702) );
and2 gate150( .a(N393), .b(N630), .O(N703) );
and2 gate151( .a(N354), .b(N635), .O(N704) );
and2 gate152( .a(N367), .b(N635), .O(N705) );
and2 gate153( .a(N380), .b(N635), .O(N706) );
and2 gate154( .a(N393), .b(N635), .O(N707) );
and2 gate155( .a(N406), .b(N640), .O(N708) );
and2 gate156( .a(N419), .b(N640), .O(N709) );
and2 gate157( .a(N432), .b(N640), .O(N710) );
and2 gate158( .a(N445), .b(N640), .O(N711) );
and2 gate159( .a(N406), .b(N645), .O(N712) );
and2 gate160( .a(N419), .b(N645), .O(N713) );
and2 gate161( .a(N432), .b(N645), .O(N714) );
and2 gate162( .a(N445), .b(N645), .O(N715) );
and2 gate163( .a(N406), .b(N650), .O(N716) );
and2 gate164( .a(N419), .b(N650), .O(N717) );
and2 gate165( .a(N432), .b(N650), .O(N718) );
and2 gate166( .a(N445), .b(N650), .O(N719) );
and2 gate167( .a(N406), .b(N655), .O(N720) );
and2 gate168( .a(N419), .b(N655), .O(N721) );
and2 gate169( .a(N432), .b(N655), .O(N722) );
and2 gate170( .a(N445), .b(N655), .O(N723) );
xor2 gate171( .a(N1), .b(N692), .O(N724) );
xor2 gate172( .a(N5), .b(N693), .O(N725) );

  xor2  gate217(.a(N694), .b(N9), .O(gate173inter0));
  nand2 gate218(.a(gate173inter0), .b(s_2), .O(gate173inter1));
  and2  gate219(.a(N694), .b(N9), .O(gate173inter2));
  inv1  gate220(.a(s_2), .O(gate173inter3));
  inv1  gate221(.a(s_3), .O(gate173inter4));
  nand2 gate222(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate223(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate224(.a(N9), .O(gate173inter7));
  inv1  gate225(.a(N694), .O(gate173inter8));
  nand2 gate226(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate227(.a(s_3), .b(gate173inter3), .O(gate173inter10));
  nor2  gate228(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate229(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate230(.a(gate173inter12), .b(gate173inter1), .O(N726));
xor2 gate174( .a(N13), .b(N695), .O(N727) );
xor2 gate175( .a(N17), .b(N696), .O(N728) );
xor2 gate176( .a(N21), .b(N697), .O(N729) );

  xor2  gate427(.a(N698), .b(N25), .O(gate177inter0));
  nand2 gate428(.a(gate177inter0), .b(s_32), .O(gate177inter1));
  and2  gate429(.a(N698), .b(N25), .O(gate177inter2));
  inv1  gate430(.a(s_32), .O(gate177inter3));
  inv1  gate431(.a(s_33), .O(gate177inter4));
  nand2 gate432(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate433(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate434(.a(N25), .O(gate177inter7));
  inv1  gate435(.a(N698), .O(gate177inter8));
  nand2 gate436(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate437(.a(s_33), .b(gate177inter3), .O(gate177inter10));
  nor2  gate438(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate439(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate440(.a(gate177inter12), .b(gate177inter1), .O(N730));

  xor2  gate399(.a(N699), .b(N29), .O(gate178inter0));
  nand2 gate400(.a(gate178inter0), .b(s_28), .O(gate178inter1));
  and2  gate401(.a(N699), .b(N29), .O(gate178inter2));
  inv1  gate402(.a(s_28), .O(gate178inter3));
  inv1  gate403(.a(s_29), .O(gate178inter4));
  nand2 gate404(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate405(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate406(.a(N29), .O(gate178inter7));
  inv1  gate407(.a(N699), .O(gate178inter8));
  nand2 gate408(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate409(.a(s_29), .b(gate178inter3), .O(gate178inter10));
  nor2  gate410(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate411(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate412(.a(gate178inter12), .b(gate178inter1), .O(N731));
xor2 gate179( .a(N33), .b(N700), .O(N732) );

  xor2  gate539(.a(N701), .b(N37), .O(gate180inter0));
  nand2 gate540(.a(gate180inter0), .b(s_48), .O(gate180inter1));
  and2  gate541(.a(N701), .b(N37), .O(gate180inter2));
  inv1  gate542(.a(s_48), .O(gate180inter3));
  inv1  gate543(.a(s_49), .O(gate180inter4));
  nand2 gate544(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate545(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate546(.a(N37), .O(gate180inter7));
  inv1  gate547(.a(N701), .O(gate180inter8));
  nand2 gate548(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate549(.a(s_49), .b(gate180inter3), .O(gate180inter10));
  nor2  gate550(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate551(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate552(.a(gate180inter12), .b(gate180inter1), .O(N733));

  xor2  gate315(.a(N702), .b(N41), .O(gate181inter0));
  nand2 gate316(.a(gate181inter0), .b(s_16), .O(gate181inter1));
  and2  gate317(.a(N702), .b(N41), .O(gate181inter2));
  inv1  gate318(.a(s_16), .O(gate181inter3));
  inv1  gate319(.a(s_17), .O(gate181inter4));
  nand2 gate320(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate321(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate322(.a(N41), .O(gate181inter7));
  inv1  gate323(.a(N702), .O(gate181inter8));
  nand2 gate324(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate325(.a(s_17), .b(gate181inter3), .O(gate181inter10));
  nor2  gate326(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate327(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate328(.a(gate181inter12), .b(gate181inter1), .O(N734));

  xor2  gate385(.a(N703), .b(N45), .O(gate182inter0));
  nand2 gate386(.a(gate182inter0), .b(s_26), .O(gate182inter1));
  and2  gate387(.a(N703), .b(N45), .O(gate182inter2));
  inv1  gate388(.a(s_26), .O(gate182inter3));
  inv1  gate389(.a(s_27), .O(gate182inter4));
  nand2 gate390(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate391(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate392(.a(N45), .O(gate182inter7));
  inv1  gate393(.a(N703), .O(gate182inter8));
  nand2 gate394(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate395(.a(s_27), .b(gate182inter3), .O(gate182inter10));
  nor2  gate396(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate397(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate398(.a(gate182inter12), .b(gate182inter1), .O(N735));
xor2 gate183( .a(N49), .b(N704), .O(N736) );

  xor2  gate273(.a(N705), .b(N53), .O(gate184inter0));
  nand2 gate274(.a(gate184inter0), .b(s_10), .O(gate184inter1));
  and2  gate275(.a(N705), .b(N53), .O(gate184inter2));
  inv1  gate276(.a(s_10), .O(gate184inter3));
  inv1  gate277(.a(s_11), .O(gate184inter4));
  nand2 gate278(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate279(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate280(.a(N53), .O(gate184inter7));
  inv1  gate281(.a(N705), .O(gate184inter8));
  nand2 gate282(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate283(.a(s_11), .b(gate184inter3), .O(gate184inter10));
  nor2  gate284(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate285(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate286(.a(gate184inter12), .b(gate184inter1), .O(N737));
xor2 gate185( .a(N57), .b(N706), .O(N738) );
xor2 gate186( .a(N61), .b(N707), .O(N739) );
xor2 gate187( .a(N65), .b(N708), .O(N740) );
xor2 gate188( .a(N69), .b(N709), .O(N741) );
xor2 gate189( .a(N73), .b(N710), .O(N742) );

  xor2  gate301(.a(N711), .b(N77), .O(gate190inter0));
  nand2 gate302(.a(gate190inter0), .b(s_14), .O(gate190inter1));
  and2  gate303(.a(N711), .b(N77), .O(gate190inter2));
  inv1  gate304(.a(s_14), .O(gate190inter3));
  inv1  gate305(.a(s_15), .O(gate190inter4));
  nand2 gate306(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate307(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate308(.a(N77), .O(gate190inter7));
  inv1  gate309(.a(N711), .O(gate190inter8));
  nand2 gate310(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate311(.a(s_15), .b(gate190inter3), .O(gate190inter10));
  nor2  gate312(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate313(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate314(.a(gate190inter12), .b(gate190inter1), .O(N743));
xor2 gate191( .a(N81), .b(N712), .O(N744) );
xor2 gate192( .a(N85), .b(N713), .O(N745) );
xor2 gate193( .a(N89), .b(N714), .O(N746) );
xor2 gate194( .a(N93), .b(N715), .O(N747) );
xor2 gate195( .a(N97), .b(N716), .O(N748) );
xor2 gate196( .a(N101), .b(N717), .O(N749) );
xor2 gate197( .a(N105), .b(N718), .O(N750) );
xor2 gate198( .a(N109), .b(N719), .O(N751) );
xor2 gate199( .a(N113), .b(N720), .O(N752) );
xor2 gate200( .a(N117), .b(N721), .O(N753) );
xor2 gate201( .a(N121), .b(N722), .O(N754) );
xor2 gate202( .a(N125), .b(N723), .O(N755) );

endmodule