module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281, s_282, s_283, s_284, s_285, s_286, s_287, s_288, s_289, s_290, s_291, s_292, s_293, s_294, s_295, s_296, s_297, s_298, s_299, s_300, s_301, s_302, s_303, s_304, s_305, s_306, s_307, s_308, s_309, s_310, s_311, s_312, s_313, s_314, s_315, s_316, s_317, s_318, s_319, s_320, s_321, s_322, s_323, s_324, s_325, s_326, s_327, s_328, s_329, s_330, s_331, s_332, s_333, s_334, s_335, s_336, s_337, s_338, s_339, s_340, s_341, s_342, s_343, s_344, s_345, s_346, s_347, s_348, s_349, s_350, s_351, s_352, s_353, s_354, s_355, s_356, s_357, s_358, s_359, s_360, s_361;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate454inter0, gate454inter1, gate454inter2, gate454inter3, gate454inter4, gate454inter5, gate454inter6, gate454inter7, gate454inter8, gate454inter9, gate454inter10, gate454inter11, gate454inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );

  xor2  gate1373(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate1374(.a(gate10inter0), .b(s_118), .O(gate10inter1));
  and2  gate1375(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate1376(.a(s_118), .O(gate10inter3));
  inv1  gate1377(.a(s_119), .O(gate10inter4));
  nand2 gate1378(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate1379(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate1380(.a(G3), .O(gate10inter7));
  inv1  gate1381(.a(G4), .O(gate10inter8));
  nand2 gate1382(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate1383(.a(s_119), .b(gate10inter3), .O(gate10inter10));
  nor2  gate1384(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate1385(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate1386(.a(gate10inter12), .b(gate10inter1), .O(G269));

  xor2  gate1177(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate1178(.a(gate11inter0), .b(s_90), .O(gate11inter1));
  and2  gate1179(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate1180(.a(s_90), .O(gate11inter3));
  inv1  gate1181(.a(s_91), .O(gate11inter4));
  nand2 gate1182(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate1183(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate1184(.a(G5), .O(gate11inter7));
  inv1  gate1185(.a(G6), .O(gate11inter8));
  nand2 gate1186(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate1187(.a(s_91), .b(gate11inter3), .O(gate11inter10));
  nor2  gate1188(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate1189(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate1190(.a(gate11inter12), .b(gate11inter1), .O(G272));

  xor2  gate1863(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate1864(.a(gate12inter0), .b(s_188), .O(gate12inter1));
  and2  gate1865(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate1866(.a(s_188), .O(gate12inter3));
  inv1  gate1867(.a(s_189), .O(gate12inter4));
  nand2 gate1868(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate1869(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate1870(.a(G7), .O(gate12inter7));
  inv1  gate1871(.a(G8), .O(gate12inter8));
  nand2 gate1872(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate1873(.a(s_189), .b(gate12inter3), .O(gate12inter10));
  nor2  gate1874(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate1875(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate1876(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate2409(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate2410(.a(gate15inter0), .b(s_266), .O(gate15inter1));
  and2  gate2411(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate2412(.a(s_266), .O(gate15inter3));
  inv1  gate2413(.a(s_267), .O(gate15inter4));
  nand2 gate2414(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate2415(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate2416(.a(G13), .O(gate15inter7));
  inv1  gate2417(.a(G14), .O(gate15inter8));
  nand2 gate2418(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate2419(.a(s_267), .b(gate15inter3), .O(gate15inter10));
  nor2  gate2420(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate2421(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate2422(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate1429(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate1430(.a(gate17inter0), .b(s_126), .O(gate17inter1));
  and2  gate1431(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate1432(.a(s_126), .O(gate17inter3));
  inv1  gate1433(.a(s_127), .O(gate17inter4));
  nand2 gate1434(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate1435(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate1436(.a(G17), .O(gate17inter7));
  inv1  gate1437(.a(G18), .O(gate17inter8));
  nand2 gate1438(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate1439(.a(s_127), .b(gate17inter3), .O(gate17inter10));
  nor2  gate1440(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate1441(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate1442(.a(gate17inter12), .b(gate17inter1), .O(G290));

  xor2  gate967(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate968(.a(gate18inter0), .b(s_60), .O(gate18inter1));
  and2  gate969(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate970(.a(s_60), .O(gate18inter3));
  inv1  gate971(.a(s_61), .O(gate18inter4));
  nand2 gate972(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate973(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate974(.a(G19), .O(gate18inter7));
  inv1  gate975(.a(G20), .O(gate18inter8));
  nand2 gate976(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate977(.a(s_61), .b(gate18inter3), .O(gate18inter10));
  nor2  gate978(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate979(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate980(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate841(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate842(.a(gate21inter0), .b(s_42), .O(gate21inter1));
  and2  gate843(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate844(.a(s_42), .O(gate21inter3));
  inv1  gate845(.a(s_43), .O(gate21inter4));
  nand2 gate846(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate847(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate848(.a(G25), .O(gate21inter7));
  inv1  gate849(.a(G26), .O(gate21inter8));
  nand2 gate850(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate851(.a(s_43), .b(gate21inter3), .O(gate21inter10));
  nor2  gate852(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate853(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate854(.a(gate21inter12), .b(gate21inter1), .O(G302));

  xor2  gate2801(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate2802(.a(gate22inter0), .b(s_322), .O(gate22inter1));
  and2  gate2803(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate2804(.a(s_322), .O(gate22inter3));
  inv1  gate2805(.a(s_323), .O(gate22inter4));
  nand2 gate2806(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate2807(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate2808(.a(G27), .O(gate22inter7));
  inv1  gate2809(.a(G28), .O(gate22inter8));
  nand2 gate2810(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate2811(.a(s_323), .b(gate22inter3), .O(gate22inter10));
  nor2  gate2812(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate2813(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate2814(.a(gate22inter12), .b(gate22inter1), .O(G305));
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate2157(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate2158(.a(gate24inter0), .b(s_230), .O(gate24inter1));
  and2  gate2159(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate2160(.a(s_230), .O(gate24inter3));
  inv1  gate2161(.a(s_231), .O(gate24inter4));
  nand2 gate2162(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate2163(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate2164(.a(G31), .O(gate24inter7));
  inv1  gate2165(.a(G32), .O(gate24inter8));
  nand2 gate2166(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate2167(.a(s_231), .b(gate24inter3), .O(gate24inter10));
  nor2  gate2168(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate2169(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate2170(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate1653(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate1654(.a(gate27inter0), .b(s_158), .O(gate27inter1));
  and2  gate1655(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate1656(.a(s_158), .O(gate27inter3));
  inv1  gate1657(.a(s_159), .O(gate27inter4));
  nand2 gate1658(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate1659(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate1660(.a(G2), .O(gate27inter7));
  inv1  gate1661(.a(G6), .O(gate27inter8));
  nand2 gate1662(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate1663(.a(s_159), .b(gate27inter3), .O(gate27inter10));
  nor2  gate1664(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate1665(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate1666(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate3053(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate3054(.a(gate29inter0), .b(s_358), .O(gate29inter1));
  and2  gate3055(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate3056(.a(s_358), .O(gate29inter3));
  inv1  gate3057(.a(s_359), .O(gate29inter4));
  nand2 gate3058(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate3059(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate3060(.a(G3), .O(gate29inter7));
  inv1  gate3061(.a(G7), .O(gate29inter8));
  nand2 gate3062(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate3063(.a(s_359), .b(gate29inter3), .O(gate29inter10));
  nor2  gate3064(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate3065(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate3066(.a(gate29inter12), .b(gate29inter1), .O(G326));

  xor2  gate813(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate814(.a(gate30inter0), .b(s_38), .O(gate30inter1));
  and2  gate815(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate816(.a(s_38), .O(gate30inter3));
  inv1  gate817(.a(s_39), .O(gate30inter4));
  nand2 gate818(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate819(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate820(.a(G11), .O(gate30inter7));
  inv1  gate821(.a(G15), .O(gate30inter8));
  nand2 gate822(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate823(.a(s_39), .b(gate30inter3), .O(gate30inter10));
  nor2  gate824(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate825(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate826(.a(gate30inter12), .b(gate30inter1), .O(G329));
nand2 gate31( .a(G4), .b(G8), .O(G332) );

  xor2  gate729(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate730(.a(gate32inter0), .b(s_26), .O(gate32inter1));
  and2  gate731(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate732(.a(s_26), .O(gate32inter3));
  inv1  gate733(.a(s_27), .O(gate32inter4));
  nand2 gate734(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate735(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate736(.a(G12), .O(gate32inter7));
  inv1  gate737(.a(G16), .O(gate32inter8));
  nand2 gate738(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate739(.a(s_27), .b(gate32inter3), .O(gate32inter10));
  nor2  gate740(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate741(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate742(.a(gate32inter12), .b(gate32inter1), .O(G335));

  xor2  gate2199(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate2200(.a(gate33inter0), .b(s_236), .O(gate33inter1));
  and2  gate2201(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate2202(.a(s_236), .O(gate33inter3));
  inv1  gate2203(.a(s_237), .O(gate33inter4));
  nand2 gate2204(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate2205(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate2206(.a(G17), .O(gate33inter7));
  inv1  gate2207(.a(G21), .O(gate33inter8));
  nand2 gate2208(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate2209(.a(s_237), .b(gate33inter3), .O(gate33inter10));
  nor2  gate2210(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate2211(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate2212(.a(gate33inter12), .b(gate33inter1), .O(G338));
nand2 gate34( .a(G25), .b(G29), .O(G341) );

  xor2  gate1723(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate1724(.a(gate35inter0), .b(s_168), .O(gate35inter1));
  and2  gate1725(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate1726(.a(s_168), .O(gate35inter3));
  inv1  gate1727(.a(s_169), .O(gate35inter4));
  nand2 gate1728(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate1729(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate1730(.a(G18), .O(gate35inter7));
  inv1  gate1731(.a(G22), .O(gate35inter8));
  nand2 gate1732(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate1733(.a(s_169), .b(gate35inter3), .O(gate35inter10));
  nor2  gate1734(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate1735(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate1736(.a(gate35inter12), .b(gate35inter1), .O(G344));
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate659(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate660(.a(gate37inter0), .b(s_16), .O(gate37inter1));
  and2  gate661(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate662(.a(s_16), .O(gate37inter3));
  inv1  gate663(.a(s_17), .O(gate37inter4));
  nand2 gate664(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate665(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate666(.a(G19), .O(gate37inter7));
  inv1  gate667(.a(G23), .O(gate37inter8));
  nand2 gate668(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate669(.a(s_17), .b(gate37inter3), .O(gate37inter10));
  nor2  gate670(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate671(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate672(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate1765(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate1766(.a(gate39inter0), .b(s_174), .O(gate39inter1));
  and2  gate1767(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate1768(.a(s_174), .O(gate39inter3));
  inv1  gate1769(.a(s_175), .O(gate39inter4));
  nand2 gate1770(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate1771(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate1772(.a(G20), .O(gate39inter7));
  inv1  gate1773(.a(G24), .O(gate39inter8));
  nand2 gate1774(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate1775(.a(s_175), .b(gate39inter3), .O(gate39inter10));
  nor2  gate1776(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate1777(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate1778(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate2395(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate2396(.a(gate41inter0), .b(s_264), .O(gate41inter1));
  and2  gate2397(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate2398(.a(s_264), .O(gate41inter3));
  inv1  gate2399(.a(s_265), .O(gate41inter4));
  nand2 gate2400(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate2401(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate2402(.a(G1), .O(gate41inter7));
  inv1  gate2403(.a(G266), .O(gate41inter8));
  nand2 gate2404(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate2405(.a(s_265), .b(gate41inter3), .O(gate41inter10));
  nor2  gate2406(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate2407(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate2408(.a(gate41inter12), .b(gate41inter1), .O(G362));

  xor2  gate2913(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate2914(.a(gate42inter0), .b(s_338), .O(gate42inter1));
  and2  gate2915(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate2916(.a(s_338), .O(gate42inter3));
  inv1  gate2917(.a(s_339), .O(gate42inter4));
  nand2 gate2918(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate2919(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate2920(.a(G2), .O(gate42inter7));
  inv1  gate2921(.a(G266), .O(gate42inter8));
  nand2 gate2922(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate2923(.a(s_339), .b(gate42inter3), .O(gate42inter10));
  nor2  gate2924(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate2925(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate2926(.a(gate42inter12), .b(gate42inter1), .O(G363));

  xor2  gate2367(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate2368(.a(gate43inter0), .b(s_260), .O(gate43inter1));
  and2  gate2369(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate2370(.a(s_260), .O(gate43inter3));
  inv1  gate2371(.a(s_261), .O(gate43inter4));
  nand2 gate2372(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate2373(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate2374(.a(G3), .O(gate43inter7));
  inv1  gate2375(.a(G269), .O(gate43inter8));
  nand2 gate2376(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate2377(.a(s_261), .b(gate43inter3), .O(gate43inter10));
  nor2  gate2378(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate2379(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate2380(.a(gate43inter12), .b(gate43inter1), .O(G364));
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );

  xor2  gate2353(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate2354(.a(gate47inter0), .b(s_258), .O(gate47inter1));
  and2  gate2355(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate2356(.a(s_258), .O(gate47inter3));
  inv1  gate2357(.a(s_259), .O(gate47inter4));
  nand2 gate2358(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate2359(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate2360(.a(G7), .O(gate47inter7));
  inv1  gate2361(.a(G275), .O(gate47inter8));
  nand2 gate2362(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate2363(.a(s_259), .b(gate47inter3), .O(gate47inter10));
  nor2  gate2364(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate2365(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate2366(.a(gate47inter12), .b(gate47inter1), .O(G368));

  xor2  gate1471(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate1472(.a(gate48inter0), .b(s_132), .O(gate48inter1));
  and2  gate1473(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate1474(.a(s_132), .O(gate48inter3));
  inv1  gate1475(.a(s_133), .O(gate48inter4));
  nand2 gate1476(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate1477(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate1478(.a(G8), .O(gate48inter7));
  inv1  gate1479(.a(G275), .O(gate48inter8));
  nand2 gate1480(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate1481(.a(s_133), .b(gate48inter3), .O(gate48inter10));
  nor2  gate1482(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate1483(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate1484(.a(gate48inter12), .b(gate48inter1), .O(G369));

  xor2  gate1849(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate1850(.a(gate49inter0), .b(s_186), .O(gate49inter1));
  and2  gate1851(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate1852(.a(s_186), .O(gate49inter3));
  inv1  gate1853(.a(s_187), .O(gate49inter4));
  nand2 gate1854(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate1855(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate1856(.a(G9), .O(gate49inter7));
  inv1  gate1857(.a(G278), .O(gate49inter8));
  nand2 gate1858(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate1859(.a(s_187), .b(gate49inter3), .O(gate49inter10));
  nor2  gate1860(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate1861(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate1862(.a(gate49inter12), .b(gate49inter1), .O(G370));

  xor2  gate2297(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate2298(.a(gate50inter0), .b(s_250), .O(gate50inter1));
  and2  gate2299(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate2300(.a(s_250), .O(gate50inter3));
  inv1  gate2301(.a(s_251), .O(gate50inter4));
  nand2 gate2302(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate2303(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate2304(.a(G10), .O(gate50inter7));
  inv1  gate2305(.a(G278), .O(gate50inter8));
  nand2 gate2306(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate2307(.a(s_251), .b(gate50inter3), .O(gate50inter10));
  nor2  gate2308(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate2309(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate2310(.a(gate50inter12), .b(gate50inter1), .O(G371));

  xor2  gate883(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate884(.a(gate51inter0), .b(s_48), .O(gate51inter1));
  and2  gate885(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate886(.a(s_48), .O(gate51inter3));
  inv1  gate887(.a(s_49), .O(gate51inter4));
  nand2 gate888(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate889(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate890(.a(G11), .O(gate51inter7));
  inv1  gate891(.a(G281), .O(gate51inter8));
  nand2 gate892(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate893(.a(s_49), .b(gate51inter3), .O(gate51inter10));
  nor2  gate894(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate895(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate896(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );

  xor2  gate2871(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate2872(.a(gate56inter0), .b(s_332), .O(gate56inter1));
  and2  gate2873(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate2874(.a(s_332), .O(gate56inter3));
  inv1  gate2875(.a(s_333), .O(gate56inter4));
  nand2 gate2876(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate2877(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate2878(.a(G16), .O(gate56inter7));
  inv1  gate2879(.a(G287), .O(gate56inter8));
  nand2 gate2880(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate2881(.a(s_333), .b(gate56inter3), .O(gate56inter10));
  nor2  gate2882(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate2883(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate2884(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate2703(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate2704(.a(gate59inter0), .b(s_308), .O(gate59inter1));
  and2  gate2705(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate2706(.a(s_308), .O(gate59inter3));
  inv1  gate2707(.a(s_309), .O(gate59inter4));
  nand2 gate2708(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate2709(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate2710(.a(G19), .O(gate59inter7));
  inv1  gate2711(.a(G293), .O(gate59inter8));
  nand2 gate2712(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate2713(.a(s_309), .b(gate59inter3), .O(gate59inter10));
  nor2  gate2714(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate2715(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate2716(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate1219(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate1220(.a(gate62inter0), .b(s_96), .O(gate62inter1));
  and2  gate1221(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate1222(.a(s_96), .O(gate62inter3));
  inv1  gate1223(.a(s_97), .O(gate62inter4));
  nand2 gate1224(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate1225(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate1226(.a(G22), .O(gate62inter7));
  inv1  gate1227(.a(G296), .O(gate62inter8));
  nand2 gate1228(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate1229(.a(s_97), .b(gate62inter3), .O(gate62inter10));
  nor2  gate1230(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate1231(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate1232(.a(gate62inter12), .b(gate62inter1), .O(G383));

  xor2  gate2927(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate2928(.a(gate63inter0), .b(s_340), .O(gate63inter1));
  and2  gate2929(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate2930(.a(s_340), .O(gate63inter3));
  inv1  gate2931(.a(s_341), .O(gate63inter4));
  nand2 gate2932(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate2933(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate2934(.a(G23), .O(gate63inter7));
  inv1  gate2935(.a(G299), .O(gate63inter8));
  nand2 gate2936(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate2937(.a(s_341), .b(gate63inter3), .O(gate63inter10));
  nor2  gate2938(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate2939(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate2940(.a(gate63inter12), .b(gate63inter1), .O(G384));

  xor2  gate2101(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate2102(.a(gate64inter0), .b(s_222), .O(gate64inter1));
  and2  gate2103(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate2104(.a(s_222), .O(gate64inter3));
  inv1  gate2105(.a(s_223), .O(gate64inter4));
  nand2 gate2106(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate2107(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate2108(.a(G24), .O(gate64inter7));
  inv1  gate2109(.a(G299), .O(gate64inter8));
  nand2 gate2110(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate2111(.a(s_223), .b(gate64inter3), .O(gate64inter10));
  nor2  gate2112(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate2113(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate2114(.a(gate64inter12), .b(gate64inter1), .O(G385));

  xor2  gate1989(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate1990(.a(gate65inter0), .b(s_206), .O(gate65inter1));
  and2  gate1991(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate1992(.a(s_206), .O(gate65inter3));
  inv1  gate1993(.a(s_207), .O(gate65inter4));
  nand2 gate1994(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate1995(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate1996(.a(G25), .O(gate65inter7));
  inv1  gate1997(.a(G302), .O(gate65inter8));
  nand2 gate1998(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate1999(.a(s_207), .b(gate65inter3), .O(gate65inter10));
  nor2  gate2000(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate2001(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate2002(.a(gate65inter12), .b(gate65inter1), .O(G386));

  xor2  gate2969(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate2970(.a(gate66inter0), .b(s_346), .O(gate66inter1));
  and2  gate2971(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate2972(.a(s_346), .O(gate66inter3));
  inv1  gate2973(.a(s_347), .O(gate66inter4));
  nand2 gate2974(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate2975(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate2976(.a(G26), .O(gate66inter7));
  inv1  gate2977(.a(G302), .O(gate66inter8));
  nand2 gate2978(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate2979(.a(s_347), .b(gate66inter3), .O(gate66inter10));
  nor2  gate2980(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate2981(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate2982(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate1709(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate1710(.a(gate71inter0), .b(s_166), .O(gate71inter1));
  and2  gate1711(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate1712(.a(s_166), .O(gate71inter3));
  inv1  gate1713(.a(s_167), .O(gate71inter4));
  nand2 gate1714(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate1715(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate1716(.a(G31), .O(gate71inter7));
  inv1  gate1717(.a(G311), .O(gate71inter8));
  nand2 gate1718(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate1719(.a(s_167), .b(gate71inter3), .O(gate71inter10));
  nor2  gate1720(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate1721(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate1722(.a(gate71inter12), .b(gate71inter1), .O(G392));

  xor2  gate2717(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate2718(.a(gate72inter0), .b(s_310), .O(gate72inter1));
  and2  gate2719(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate2720(.a(s_310), .O(gate72inter3));
  inv1  gate2721(.a(s_311), .O(gate72inter4));
  nand2 gate2722(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate2723(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate2724(.a(G32), .O(gate72inter7));
  inv1  gate2725(.a(G311), .O(gate72inter8));
  nand2 gate2726(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate2727(.a(s_311), .b(gate72inter3), .O(gate72inter10));
  nor2  gate2728(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate2729(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate2730(.a(gate72inter12), .b(gate72inter1), .O(G393));
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate2549(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate2550(.a(gate74inter0), .b(s_286), .O(gate74inter1));
  and2  gate2551(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate2552(.a(s_286), .O(gate74inter3));
  inv1  gate2553(.a(s_287), .O(gate74inter4));
  nand2 gate2554(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate2555(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate2556(.a(G5), .O(gate74inter7));
  inv1  gate2557(.a(G314), .O(gate74inter8));
  nand2 gate2558(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate2559(.a(s_287), .b(gate74inter3), .O(gate74inter10));
  nor2  gate2560(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate2561(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate2562(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );

  xor2  gate2059(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate2060(.a(gate76inter0), .b(s_216), .O(gate76inter1));
  and2  gate2061(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate2062(.a(s_216), .O(gate76inter3));
  inv1  gate2063(.a(s_217), .O(gate76inter4));
  nand2 gate2064(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate2065(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate2066(.a(G13), .O(gate76inter7));
  inv1  gate2067(.a(G317), .O(gate76inter8));
  nand2 gate2068(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate2069(.a(s_217), .b(gate76inter3), .O(gate76inter10));
  nor2  gate2070(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate2071(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate2072(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate757(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate758(.a(gate78inter0), .b(s_30), .O(gate78inter1));
  and2  gate759(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate760(.a(s_30), .O(gate78inter3));
  inv1  gate761(.a(s_31), .O(gate78inter4));
  nand2 gate762(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate763(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate764(.a(G6), .O(gate78inter7));
  inv1  gate765(.a(G320), .O(gate78inter8));
  nand2 gate766(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate767(.a(s_31), .b(gate78inter3), .O(gate78inter10));
  nor2  gate768(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate769(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate770(.a(gate78inter12), .b(gate78inter1), .O(G399));

  xor2  gate2143(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate2144(.a(gate79inter0), .b(s_228), .O(gate79inter1));
  and2  gate2145(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate2146(.a(s_228), .O(gate79inter3));
  inv1  gate2147(.a(s_229), .O(gate79inter4));
  nand2 gate2148(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate2149(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate2150(.a(G10), .O(gate79inter7));
  inv1  gate2151(.a(G323), .O(gate79inter8));
  nand2 gate2152(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate2153(.a(s_229), .b(gate79inter3), .O(gate79inter10));
  nor2  gate2154(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate2155(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate2156(.a(gate79inter12), .b(gate79inter1), .O(G400));

  xor2  gate1457(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate1458(.a(gate80inter0), .b(s_130), .O(gate80inter1));
  and2  gate1459(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate1460(.a(s_130), .O(gate80inter3));
  inv1  gate1461(.a(s_131), .O(gate80inter4));
  nand2 gate1462(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate1463(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate1464(.a(G14), .O(gate80inter7));
  inv1  gate1465(.a(G323), .O(gate80inter8));
  nand2 gate1466(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate1467(.a(s_131), .b(gate80inter3), .O(gate80inter10));
  nor2  gate1468(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate1469(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate1470(.a(gate80inter12), .b(gate80inter1), .O(G401));

  xor2  gate589(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate590(.a(gate81inter0), .b(s_6), .O(gate81inter1));
  and2  gate591(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate592(.a(s_6), .O(gate81inter3));
  inv1  gate593(.a(s_7), .O(gate81inter4));
  nand2 gate594(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate595(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate596(.a(G3), .O(gate81inter7));
  inv1  gate597(.a(G326), .O(gate81inter8));
  nand2 gate598(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate599(.a(s_7), .b(gate81inter3), .O(gate81inter10));
  nor2  gate600(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate601(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate602(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate771(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate772(.a(gate85inter0), .b(s_32), .O(gate85inter1));
  and2  gate773(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate774(.a(s_32), .O(gate85inter3));
  inv1  gate775(.a(s_33), .O(gate85inter4));
  nand2 gate776(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate777(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate778(.a(G4), .O(gate85inter7));
  inv1  gate779(.a(G332), .O(gate85inter8));
  nand2 gate780(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate781(.a(s_33), .b(gate85inter3), .O(gate85inter10));
  nor2  gate782(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate783(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate784(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );

  xor2  gate1331(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate1332(.a(gate87inter0), .b(s_112), .O(gate87inter1));
  and2  gate1333(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate1334(.a(s_112), .O(gate87inter3));
  inv1  gate1335(.a(s_113), .O(gate87inter4));
  nand2 gate1336(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate1337(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate1338(.a(G12), .O(gate87inter7));
  inv1  gate1339(.a(G335), .O(gate87inter8));
  nand2 gate1340(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate1341(.a(s_113), .b(gate87inter3), .O(gate87inter10));
  nor2  gate1342(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate1343(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate1344(.a(gate87inter12), .b(gate87inter1), .O(G408));

  xor2  gate1401(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate1402(.a(gate88inter0), .b(s_122), .O(gate88inter1));
  and2  gate1403(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate1404(.a(s_122), .O(gate88inter3));
  inv1  gate1405(.a(s_123), .O(gate88inter4));
  nand2 gate1406(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate1407(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate1408(.a(G16), .O(gate88inter7));
  inv1  gate1409(.a(G335), .O(gate88inter8));
  nand2 gate1410(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate1411(.a(s_123), .b(gate88inter3), .O(gate88inter10));
  nor2  gate1412(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate1413(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate1414(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate1149(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate1150(.a(gate91inter0), .b(s_86), .O(gate91inter1));
  and2  gate1151(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate1152(.a(s_86), .O(gate91inter3));
  inv1  gate1153(.a(s_87), .O(gate91inter4));
  nand2 gate1154(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate1155(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate1156(.a(G25), .O(gate91inter7));
  inv1  gate1157(.a(G341), .O(gate91inter8));
  nand2 gate1158(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate1159(.a(s_87), .b(gate91inter3), .O(gate91inter10));
  nor2  gate1160(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate1161(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate1162(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );

  xor2  gate2017(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate2018(.a(gate93inter0), .b(s_210), .O(gate93inter1));
  and2  gate2019(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate2020(.a(s_210), .O(gate93inter3));
  inv1  gate2021(.a(s_211), .O(gate93inter4));
  nand2 gate2022(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate2023(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate2024(.a(G18), .O(gate93inter7));
  inv1  gate2025(.a(G344), .O(gate93inter8));
  nand2 gate2026(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate2027(.a(s_211), .b(gate93inter3), .O(gate93inter10));
  nor2  gate2028(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate2029(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate2030(.a(gate93inter12), .b(gate93inter1), .O(G414));

  xor2  gate1793(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate1794(.a(gate94inter0), .b(s_178), .O(gate94inter1));
  and2  gate1795(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate1796(.a(s_178), .O(gate94inter3));
  inv1  gate1797(.a(s_179), .O(gate94inter4));
  nand2 gate1798(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate1799(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate1800(.a(G22), .O(gate94inter7));
  inv1  gate1801(.a(G344), .O(gate94inter8));
  nand2 gate1802(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate1803(.a(s_179), .b(gate94inter3), .O(gate94inter10));
  nor2  gate1804(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate1805(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate1806(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate2241(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate2242(.a(gate96inter0), .b(s_242), .O(gate96inter1));
  and2  gate2243(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate2244(.a(s_242), .O(gate96inter3));
  inv1  gate2245(.a(s_243), .O(gate96inter4));
  nand2 gate2246(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate2247(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate2248(.a(G30), .O(gate96inter7));
  inv1  gate2249(.a(G347), .O(gate96inter8));
  nand2 gate2250(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate2251(.a(s_243), .b(gate96inter3), .O(gate96inter10));
  nor2  gate2252(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate2253(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate2254(.a(gate96inter12), .b(gate96inter1), .O(G417));
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate1037(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate1038(.a(gate98inter0), .b(s_70), .O(gate98inter1));
  and2  gate1039(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate1040(.a(s_70), .O(gate98inter3));
  inv1  gate1041(.a(s_71), .O(gate98inter4));
  nand2 gate1042(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1043(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1044(.a(G23), .O(gate98inter7));
  inv1  gate1045(.a(G350), .O(gate98inter8));
  nand2 gate1046(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1047(.a(s_71), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1048(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1049(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1050(.a(gate98inter12), .b(gate98inter1), .O(G419));

  xor2  gate1527(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate1528(.a(gate99inter0), .b(s_140), .O(gate99inter1));
  and2  gate1529(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate1530(.a(s_140), .O(gate99inter3));
  inv1  gate1531(.a(s_141), .O(gate99inter4));
  nand2 gate1532(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate1533(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate1534(.a(G27), .O(gate99inter7));
  inv1  gate1535(.a(G353), .O(gate99inter8));
  nand2 gate1536(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate1537(.a(s_141), .b(gate99inter3), .O(gate99inter10));
  nor2  gate1538(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate1539(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate1540(.a(gate99inter12), .b(gate99inter1), .O(G420));

  xor2  gate1107(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate1108(.a(gate100inter0), .b(s_80), .O(gate100inter1));
  and2  gate1109(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate1110(.a(s_80), .O(gate100inter3));
  inv1  gate1111(.a(s_81), .O(gate100inter4));
  nand2 gate1112(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate1113(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate1114(.a(G31), .O(gate100inter7));
  inv1  gate1115(.a(G353), .O(gate100inter8));
  nand2 gate1116(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate1117(.a(s_81), .b(gate100inter3), .O(gate100inter10));
  nor2  gate1118(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate1119(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate1120(.a(gate100inter12), .b(gate100inter1), .O(G421));

  xor2  gate1751(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate1752(.a(gate101inter0), .b(s_172), .O(gate101inter1));
  and2  gate1753(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate1754(.a(s_172), .O(gate101inter3));
  inv1  gate1755(.a(s_173), .O(gate101inter4));
  nand2 gate1756(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate1757(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate1758(.a(G20), .O(gate101inter7));
  inv1  gate1759(.a(G356), .O(gate101inter8));
  nand2 gate1760(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate1761(.a(s_173), .b(gate101inter3), .O(gate101inter10));
  nor2  gate1762(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate1763(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate1764(.a(gate101inter12), .b(gate101inter1), .O(G422));

  xor2  gate1555(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate1556(.a(gate102inter0), .b(s_144), .O(gate102inter1));
  and2  gate1557(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate1558(.a(s_144), .O(gate102inter3));
  inv1  gate1559(.a(s_145), .O(gate102inter4));
  nand2 gate1560(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate1561(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate1562(.a(G24), .O(gate102inter7));
  inv1  gate1563(.a(G356), .O(gate102inter8));
  nand2 gate1564(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate1565(.a(s_145), .b(gate102inter3), .O(gate102inter10));
  nor2  gate1566(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate1567(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate1568(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate2465(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate2466(.a(gate104inter0), .b(s_274), .O(gate104inter1));
  and2  gate2467(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate2468(.a(s_274), .O(gate104inter3));
  inv1  gate2469(.a(s_275), .O(gate104inter4));
  nand2 gate2470(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate2471(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate2472(.a(G32), .O(gate104inter7));
  inv1  gate2473(.a(G359), .O(gate104inter8));
  nand2 gate2474(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate2475(.a(s_275), .b(gate104inter3), .O(gate104inter10));
  nor2  gate2476(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate2477(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate2478(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate1261(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate1262(.a(gate106inter0), .b(s_102), .O(gate106inter1));
  and2  gate1263(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate1264(.a(s_102), .O(gate106inter3));
  inv1  gate1265(.a(s_103), .O(gate106inter4));
  nand2 gate1266(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate1267(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate1268(.a(G364), .O(gate106inter7));
  inv1  gate1269(.a(G365), .O(gate106inter8));
  nand2 gate1270(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate1271(.a(s_103), .b(gate106inter3), .O(gate106inter10));
  nor2  gate1272(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate1273(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate1274(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate1891(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate1892(.a(gate108inter0), .b(s_192), .O(gate108inter1));
  and2  gate1893(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate1894(.a(s_192), .O(gate108inter3));
  inv1  gate1895(.a(s_193), .O(gate108inter4));
  nand2 gate1896(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate1897(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate1898(.a(G368), .O(gate108inter7));
  inv1  gate1899(.a(G369), .O(gate108inter8));
  nand2 gate1900(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate1901(.a(s_193), .b(gate108inter3), .O(gate108inter10));
  nor2  gate1902(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate1903(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate1904(.a(gate108inter12), .b(gate108inter1), .O(G435));
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate1611(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate1612(.a(gate112inter0), .b(s_152), .O(gate112inter1));
  and2  gate1613(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate1614(.a(s_152), .O(gate112inter3));
  inv1  gate1615(.a(s_153), .O(gate112inter4));
  nand2 gate1616(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate1617(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate1618(.a(G376), .O(gate112inter7));
  inv1  gate1619(.a(G377), .O(gate112inter8));
  nand2 gate1620(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate1621(.a(s_153), .b(gate112inter3), .O(gate112inter10));
  nor2  gate1622(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate1623(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate1624(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );

  xor2  gate2605(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate2606(.a(gate114inter0), .b(s_294), .O(gate114inter1));
  and2  gate2607(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate2608(.a(s_294), .O(gate114inter3));
  inv1  gate2609(.a(s_295), .O(gate114inter4));
  nand2 gate2610(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate2611(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate2612(.a(G380), .O(gate114inter7));
  inv1  gate2613(.a(G381), .O(gate114inter8));
  nand2 gate2614(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate2615(.a(s_295), .b(gate114inter3), .O(gate114inter10));
  nor2  gate2616(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate2617(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate2618(.a(gate114inter12), .b(gate114inter1), .O(G453));
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate2255(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate2256(.a(gate117inter0), .b(s_244), .O(gate117inter1));
  and2  gate2257(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate2258(.a(s_244), .O(gate117inter3));
  inv1  gate2259(.a(s_245), .O(gate117inter4));
  nand2 gate2260(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate2261(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate2262(.a(G386), .O(gate117inter7));
  inv1  gate2263(.a(G387), .O(gate117inter8));
  nand2 gate2264(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate2265(.a(s_245), .b(gate117inter3), .O(gate117inter10));
  nor2  gate2266(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate2267(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate2268(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate631(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate632(.a(gate119inter0), .b(s_12), .O(gate119inter1));
  and2  gate633(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate634(.a(s_12), .O(gate119inter3));
  inv1  gate635(.a(s_13), .O(gate119inter4));
  nand2 gate636(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate637(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate638(.a(G390), .O(gate119inter7));
  inv1  gate639(.a(G391), .O(gate119inter8));
  nand2 gate640(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate641(.a(s_13), .b(gate119inter3), .O(gate119inter10));
  nor2  gate642(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate643(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate644(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );

  xor2  gate1583(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate1584(.a(gate122inter0), .b(s_148), .O(gate122inter1));
  and2  gate1585(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate1586(.a(s_148), .O(gate122inter3));
  inv1  gate1587(.a(s_149), .O(gate122inter4));
  nand2 gate1588(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate1589(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate1590(.a(G396), .O(gate122inter7));
  inv1  gate1591(.a(G397), .O(gate122inter8));
  nand2 gate1592(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate1593(.a(s_149), .b(gate122inter3), .O(gate122inter10));
  nor2  gate1594(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate1595(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate1596(.a(gate122inter12), .b(gate122inter1), .O(G477));
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate1009(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate1010(.a(gate126inter0), .b(s_66), .O(gate126inter1));
  and2  gate1011(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate1012(.a(s_66), .O(gate126inter3));
  inv1  gate1013(.a(s_67), .O(gate126inter4));
  nand2 gate1014(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate1015(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate1016(.a(G404), .O(gate126inter7));
  inv1  gate1017(.a(G405), .O(gate126inter8));
  nand2 gate1018(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate1019(.a(s_67), .b(gate126inter3), .O(gate126inter10));
  nor2  gate1020(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate1021(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate1022(.a(gate126inter12), .b(gate126inter1), .O(G489));

  xor2  gate2087(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate2088(.a(gate127inter0), .b(s_220), .O(gate127inter1));
  and2  gate2089(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate2090(.a(s_220), .O(gate127inter3));
  inv1  gate2091(.a(s_221), .O(gate127inter4));
  nand2 gate2092(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate2093(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate2094(.a(G406), .O(gate127inter7));
  inv1  gate2095(.a(G407), .O(gate127inter8));
  nand2 gate2096(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate2097(.a(s_221), .b(gate127inter3), .O(gate127inter10));
  nor2  gate2098(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate2099(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate2100(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate2185(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate2186(.a(gate131inter0), .b(s_234), .O(gate131inter1));
  and2  gate2187(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate2188(.a(s_234), .O(gate131inter3));
  inv1  gate2189(.a(s_235), .O(gate131inter4));
  nand2 gate2190(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate2191(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate2192(.a(G414), .O(gate131inter7));
  inv1  gate2193(.a(G415), .O(gate131inter8));
  nand2 gate2194(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate2195(.a(s_235), .b(gate131inter3), .O(gate131inter10));
  nor2  gate2196(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate2197(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate2198(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );

  xor2  gate953(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate954(.a(gate134inter0), .b(s_58), .O(gate134inter1));
  and2  gate955(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate956(.a(s_58), .O(gate134inter3));
  inv1  gate957(.a(s_59), .O(gate134inter4));
  nand2 gate958(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate959(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate960(.a(G420), .O(gate134inter7));
  inv1  gate961(.a(G421), .O(gate134inter8));
  nand2 gate962(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate963(.a(s_59), .b(gate134inter3), .O(gate134inter10));
  nor2  gate964(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate965(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate966(.a(gate134inter12), .b(gate134inter1), .O(G513));

  xor2  gate2689(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate2690(.a(gate135inter0), .b(s_306), .O(gate135inter1));
  and2  gate2691(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate2692(.a(s_306), .O(gate135inter3));
  inv1  gate2693(.a(s_307), .O(gate135inter4));
  nand2 gate2694(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate2695(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate2696(.a(G422), .O(gate135inter7));
  inv1  gate2697(.a(G423), .O(gate135inter8));
  nand2 gate2698(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate2699(.a(s_307), .b(gate135inter3), .O(gate135inter10));
  nor2  gate2700(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate2701(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate2702(.a(gate135inter12), .b(gate135inter1), .O(G516));

  xor2  gate1975(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate1976(.a(gate136inter0), .b(s_204), .O(gate136inter1));
  and2  gate1977(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate1978(.a(s_204), .O(gate136inter3));
  inv1  gate1979(.a(s_205), .O(gate136inter4));
  nand2 gate1980(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate1981(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate1982(.a(G424), .O(gate136inter7));
  inv1  gate1983(.a(G425), .O(gate136inter8));
  nand2 gate1984(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate1985(.a(s_205), .b(gate136inter3), .O(gate136inter10));
  nor2  gate1986(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate1987(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate1988(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate827(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate828(.a(gate138inter0), .b(s_40), .O(gate138inter1));
  and2  gate829(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate830(.a(s_40), .O(gate138inter3));
  inv1  gate831(.a(s_41), .O(gate138inter4));
  nand2 gate832(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate833(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate834(.a(G432), .O(gate138inter7));
  inv1  gate835(.a(G435), .O(gate138inter8));
  nand2 gate836(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate837(.a(s_41), .b(gate138inter3), .O(gate138inter10));
  nor2  gate838(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate839(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate840(.a(gate138inter12), .b(gate138inter1), .O(G525));

  xor2  gate1485(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate1486(.a(gate139inter0), .b(s_134), .O(gate139inter1));
  and2  gate1487(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate1488(.a(s_134), .O(gate139inter3));
  inv1  gate1489(.a(s_135), .O(gate139inter4));
  nand2 gate1490(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate1491(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate1492(.a(G438), .O(gate139inter7));
  inv1  gate1493(.a(G441), .O(gate139inter8));
  nand2 gate1494(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate1495(.a(s_135), .b(gate139inter3), .O(gate139inter10));
  nor2  gate1496(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate1497(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate1498(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate2941(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate2942(.a(gate142inter0), .b(s_342), .O(gate142inter1));
  and2  gate2943(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate2944(.a(s_342), .O(gate142inter3));
  inv1  gate2945(.a(s_343), .O(gate142inter4));
  nand2 gate2946(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate2947(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate2948(.a(G456), .O(gate142inter7));
  inv1  gate2949(.a(G459), .O(gate142inter8));
  nand2 gate2950(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate2951(.a(s_343), .b(gate142inter3), .O(gate142inter10));
  nor2  gate2952(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate2953(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate2954(.a(gate142inter12), .b(gate142inter1), .O(G537));

  xor2  gate1821(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate1822(.a(gate143inter0), .b(s_182), .O(gate143inter1));
  and2  gate1823(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate1824(.a(s_182), .O(gate143inter3));
  inv1  gate1825(.a(s_183), .O(gate143inter4));
  nand2 gate1826(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate1827(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate1828(.a(G462), .O(gate143inter7));
  inv1  gate1829(.a(G465), .O(gate143inter8));
  nand2 gate1830(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate1831(.a(s_183), .b(gate143inter3), .O(gate143inter10));
  nor2  gate1832(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate1833(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate1834(.a(gate143inter12), .b(gate143inter1), .O(G540));
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate1625(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate1626(.a(gate147inter0), .b(s_154), .O(gate147inter1));
  and2  gate1627(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate1628(.a(s_154), .O(gate147inter3));
  inv1  gate1629(.a(s_155), .O(gate147inter4));
  nand2 gate1630(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate1631(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate1632(.a(G486), .O(gate147inter7));
  inv1  gate1633(.a(G489), .O(gate147inter8));
  nand2 gate1634(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate1635(.a(s_155), .b(gate147inter3), .O(gate147inter10));
  nor2  gate1636(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate1637(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate1638(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate1597(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate1598(.a(gate150inter0), .b(s_150), .O(gate150inter1));
  and2  gate1599(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate1600(.a(s_150), .O(gate150inter3));
  inv1  gate1601(.a(s_151), .O(gate150inter4));
  nand2 gate1602(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate1603(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate1604(.a(G504), .O(gate150inter7));
  inv1  gate1605(.a(G507), .O(gate150inter8));
  nand2 gate1606(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate1607(.a(s_151), .b(gate150inter3), .O(gate150inter10));
  nor2  gate1608(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate1609(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate1610(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate1317(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate1318(.a(gate156inter0), .b(s_110), .O(gate156inter1));
  and2  gate1319(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate1320(.a(s_110), .O(gate156inter3));
  inv1  gate1321(.a(s_111), .O(gate156inter4));
  nand2 gate1322(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate1323(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate1324(.a(G435), .O(gate156inter7));
  inv1  gate1325(.a(G525), .O(gate156inter8));
  nand2 gate1326(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate1327(.a(s_111), .b(gate156inter3), .O(gate156inter10));
  nor2  gate1328(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate1329(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate1330(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate2381(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate2382(.a(gate158inter0), .b(s_262), .O(gate158inter1));
  and2  gate2383(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate2384(.a(s_262), .O(gate158inter3));
  inv1  gate2385(.a(s_263), .O(gate158inter4));
  nand2 gate2386(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate2387(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate2388(.a(G441), .O(gate158inter7));
  inv1  gate2389(.a(G528), .O(gate158inter8));
  nand2 gate2390(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate2391(.a(s_263), .b(gate158inter3), .O(gate158inter10));
  nor2  gate2392(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate2393(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate2394(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate1695(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate1696(.a(gate164inter0), .b(s_164), .O(gate164inter1));
  and2  gate1697(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate1698(.a(s_164), .O(gate164inter3));
  inv1  gate1699(.a(s_165), .O(gate164inter4));
  nand2 gate1700(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate1701(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate1702(.a(G459), .O(gate164inter7));
  inv1  gate1703(.a(G537), .O(gate164inter8));
  nand2 gate1704(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate1705(.a(s_165), .b(gate164inter3), .O(gate164inter10));
  nor2  gate1706(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate1707(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate1708(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );

  xor2  gate785(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate786(.a(gate166inter0), .b(s_34), .O(gate166inter1));
  and2  gate787(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate788(.a(s_34), .O(gate166inter3));
  inv1  gate789(.a(s_35), .O(gate166inter4));
  nand2 gate790(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate791(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate792(.a(G465), .O(gate166inter7));
  inv1  gate793(.a(G540), .O(gate166inter8));
  nand2 gate794(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate795(.a(s_35), .b(gate166inter3), .O(gate166inter10));
  nor2  gate796(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate797(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate798(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );

  xor2  gate2311(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate2312(.a(gate171inter0), .b(s_252), .O(gate171inter1));
  and2  gate2313(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate2314(.a(s_252), .O(gate171inter3));
  inv1  gate2315(.a(s_253), .O(gate171inter4));
  nand2 gate2316(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate2317(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate2318(.a(G480), .O(gate171inter7));
  inv1  gate2319(.a(G549), .O(gate171inter8));
  nand2 gate2320(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate2321(.a(s_253), .b(gate171inter3), .O(gate171inter10));
  nor2  gate2322(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate2323(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate2324(.a(gate171inter12), .b(gate171inter1), .O(G588));

  xor2  gate701(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate702(.a(gate172inter0), .b(s_22), .O(gate172inter1));
  and2  gate703(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate704(.a(s_22), .O(gate172inter3));
  inv1  gate705(.a(s_23), .O(gate172inter4));
  nand2 gate706(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate707(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate708(.a(G483), .O(gate172inter7));
  inv1  gate709(.a(G549), .O(gate172inter8));
  nand2 gate710(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate711(.a(s_23), .b(gate172inter3), .O(gate172inter10));
  nor2  gate712(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate713(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate714(.a(gate172inter12), .b(gate172inter1), .O(G589));

  xor2  gate2731(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate2732(.a(gate173inter0), .b(s_312), .O(gate173inter1));
  and2  gate2733(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate2734(.a(s_312), .O(gate173inter3));
  inv1  gate2735(.a(s_313), .O(gate173inter4));
  nand2 gate2736(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate2737(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate2738(.a(G486), .O(gate173inter7));
  inv1  gate2739(.a(G552), .O(gate173inter8));
  nand2 gate2740(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate2741(.a(s_313), .b(gate173inter3), .O(gate173inter10));
  nor2  gate2742(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate2743(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate2744(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate2339(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate2340(.a(gate175inter0), .b(s_256), .O(gate175inter1));
  and2  gate2341(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate2342(.a(s_256), .O(gate175inter3));
  inv1  gate2343(.a(s_257), .O(gate175inter4));
  nand2 gate2344(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate2345(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate2346(.a(G492), .O(gate175inter7));
  inv1  gate2347(.a(G555), .O(gate175inter8));
  nand2 gate2348(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate2349(.a(s_257), .b(gate175inter3), .O(gate175inter10));
  nor2  gate2350(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate2351(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate2352(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );

  xor2  gate1233(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate1234(.a(gate177inter0), .b(s_98), .O(gate177inter1));
  and2  gate1235(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate1236(.a(s_98), .O(gate177inter3));
  inv1  gate1237(.a(s_99), .O(gate177inter4));
  nand2 gate1238(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate1239(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate1240(.a(G498), .O(gate177inter7));
  inv1  gate1241(.a(G558), .O(gate177inter8));
  nand2 gate1242(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate1243(.a(s_99), .b(gate177inter3), .O(gate177inter10));
  nor2  gate1244(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate1245(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate1246(.a(gate177inter12), .b(gate177inter1), .O(G594));
nand2 gate178( .a(G501), .b(G558), .O(G595) );

  xor2  gate2843(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate2844(.a(gate179inter0), .b(s_328), .O(gate179inter1));
  and2  gate2845(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate2846(.a(s_328), .O(gate179inter3));
  inv1  gate2847(.a(s_329), .O(gate179inter4));
  nand2 gate2848(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate2849(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate2850(.a(G504), .O(gate179inter7));
  inv1  gate2851(.a(G561), .O(gate179inter8));
  nand2 gate2852(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate2853(.a(s_329), .b(gate179inter3), .O(gate179inter10));
  nor2  gate2854(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate2855(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate2856(.a(gate179inter12), .b(gate179inter1), .O(G596));
nand2 gate180( .a(G507), .b(G561), .O(G597) );

  xor2  gate995(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate996(.a(gate181inter0), .b(s_64), .O(gate181inter1));
  and2  gate997(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate998(.a(s_64), .O(gate181inter3));
  inv1  gate999(.a(s_65), .O(gate181inter4));
  nand2 gate1000(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate1001(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate1002(.a(G510), .O(gate181inter7));
  inv1  gate1003(.a(G564), .O(gate181inter8));
  nand2 gate1004(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate1005(.a(s_65), .b(gate181inter3), .O(gate181inter10));
  nor2  gate1006(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate1007(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate1008(.a(gate181inter12), .b(gate181inter1), .O(G598));

  xor2  gate603(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate604(.a(gate182inter0), .b(s_8), .O(gate182inter1));
  and2  gate605(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate606(.a(s_8), .O(gate182inter3));
  inv1  gate607(.a(s_9), .O(gate182inter4));
  nand2 gate608(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate609(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate610(.a(G513), .O(gate182inter7));
  inv1  gate611(.a(G564), .O(gate182inter8));
  nand2 gate612(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate613(.a(s_9), .b(gate182inter3), .O(gate182inter10));
  nor2  gate614(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate615(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate616(.a(gate182inter12), .b(gate182inter1), .O(G599));

  xor2  gate1667(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate1668(.a(gate183inter0), .b(s_160), .O(gate183inter1));
  and2  gate1669(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate1670(.a(s_160), .O(gate183inter3));
  inv1  gate1671(.a(s_161), .O(gate183inter4));
  nand2 gate1672(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate1673(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate1674(.a(G516), .O(gate183inter7));
  inv1  gate1675(.a(G567), .O(gate183inter8));
  nand2 gate1676(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate1677(.a(s_161), .b(gate183inter3), .O(gate183inter10));
  nor2  gate1678(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate1679(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate1680(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate1919(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate1920(.a(gate185inter0), .b(s_196), .O(gate185inter1));
  and2  gate1921(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate1922(.a(s_196), .O(gate185inter3));
  inv1  gate1923(.a(s_197), .O(gate185inter4));
  nand2 gate1924(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate1925(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate1926(.a(G570), .O(gate185inter7));
  inv1  gate1927(.a(G571), .O(gate185inter8));
  nand2 gate1928(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate1929(.a(s_197), .b(gate185inter3), .O(gate185inter10));
  nor2  gate1930(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate1931(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate1932(.a(gate185inter12), .b(gate185inter1), .O(G602));
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );

  xor2  gate2577(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate2578(.a(gate189inter0), .b(s_290), .O(gate189inter1));
  and2  gate2579(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate2580(.a(s_290), .O(gate189inter3));
  inv1  gate2581(.a(s_291), .O(gate189inter4));
  nand2 gate2582(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate2583(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate2584(.a(G578), .O(gate189inter7));
  inv1  gate2585(.a(G579), .O(gate189inter8));
  nand2 gate2586(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate2587(.a(s_291), .b(gate189inter3), .O(gate189inter10));
  nor2  gate2588(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate2589(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate2590(.a(gate189inter12), .b(gate189inter1), .O(G622));
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate1779(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate1780(.a(gate193inter0), .b(s_176), .O(gate193inter1));
  and2  gate1781(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate1782(.a(s_176), .O(gate193inter3));
  inv1  gate1783(.a(s_177), .O(gate193inter4));
  nand2 gate1784(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate1785(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate1786(.a(G586), .O(gate193inter7));
  inv1  gate1787(.a(G587), .O(gate193inter8));
  nand2 gate1788(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate1789(.a(s_177), .b(gate193inter3), .O(gate193inter10));
  nor2  gate1790(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate1791(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate1792(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate2983(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate2984(.a(gate195inter0), .b(s_348), .O(gate195inter1));
  and2  gate2985(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate2986(.a(s_348), .O(gate195inter3));
  inv1  gate2987(.a(s_349), .O(gate195inter4));
  nand2 gate2988(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate2989(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate2990(.a(G590), .O(gate195inter7));
  inv1  gate2991(.a(G591), .O(gate195inter8));
  nand2 gate2992(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate2993(.a(s_349), .b(gate195inter3), .O(gate195inter10));
  nor2  gate2994(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate2995(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate2996(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate2073(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate2074(.a(gate198inter0), .b(s_218), .O(gate198inter1));
  and2  gate2075(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate2076(.a(s_218), .O(gate198inter3));
  inv1  gate2077(.a(s_219), .O(gate198inter4));
  nand2 gate2078(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate2079(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate2080(.a(G596), .O(gate198inter7));
  inv1  gate2081(.a(G597), .O(gate198inter8));
  nand2 gate2082(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate2083(.a(s_219), .b(gate198inter3), .O(gate198inter10));
  nor2  gate2084(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate2085(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate2086(.a(gate198inter12), .b(gate198inter1), .O(G657));

  xor2  gate2591(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate2592(.a(gate199inter0), .b(s_292), .O(gate199inter1));
  and2  gate2593(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate2594(.a(s_292), .O(gate199inter3));
  inv1  gate2595(.a(s_293), .O(gate199inter4));
  nand2 gate2596(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate2597(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate2598(.a(G598), .O(gate199inter7));
  inv1  gate2599(.a(G599), .O(gate199inter8));
  nand2 gate2600(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate2601(.a(s_293), .b(gate199inter3), .O(gate199inter10));
  nor2  gate2602(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate2603(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate2604(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate2325(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate2326(.a(gate206inter0), .b(s_254), .O(gate206inter1));
  and2  gate2327(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate2328(.a(s_254), .O(gate206inter3));
  inv1  gate2329(.a(s_255), .O(gate206inter4));
  nand2 gate2330(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate2331(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate2332(.a(G632), .O(gate206inter7));
  inv1  gate2333(.a(G637), .O(gate206inter8));
  nand2 gate2334(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate2335(.a(s_255), .b(gate206inter3), .O(gate206inter10));
  nor2  gate2336(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate2337(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate2338(.a(gate206inter12), .b(gate206inter1), .O(G681));

  xor2  gate869(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate870(.a(gate207inter0), .b(s_46), .O(gate207inter1));
  and2  gate871(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate872(.a(s_46), .O(gate207inter3));
  inv1  gate873(.a(s_47), .O(gate207inter4));
  nand2 gate874(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate875(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate876(.a(G622), .O(gate207inter7));
  inv1  gate877(.a(G632), .O(gate207inter8));
  nand2 gate878(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate879(.a(s_47), .b(gate207inter3), .O(gate207inter10));
  nor2  gate880(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate881(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate882(.a(gate207inter12), .b(gate207inter1), .O(G684));

  xor2  gate3067(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate3068(.a(gate208inter0), .b(s_360), .O(gate208inter1));
  and2  gate3069(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate3070(.a(s_360), .O(gate208inter3));
  inv1  gate3071(.a(s_361), .O(gate208inter4));
  nand2 gate3072(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate3073(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate3074(.a(G627), .O(gate208inter7));
  inv1  gate3075(.a(G637), .O(gate208inter8));
  nand2 gate3076(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate3077(.a(s_361), .b(gate208inter3), .O(gate208inter10));
  nor2  gate3078(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate3079(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate3080(.a(gate208inter12), .b(gate208inter1), .O(G687));
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate2563(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate2564(.a(gate213inter0), .b(s_288), .O(gate213inter1));
  and2  gate2565(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate2566(.a(s_288), .O(gate213inter3));
  inv1  gate2567(.a(s_289), .O(gate213inter4));
  nand2 gate2568(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate2569(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate2570(.a(G602), .O(gate213inter7));
  inv1  gate2571(.a(G672), .O(gate213inter8));
  nand2 gate2572(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate2573(.a(s_289), .b(gate213inter3), .O(gate213inter10));
  nor2  gate2574(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate2575(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate2576(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate2675(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate2676(.a(gate215inter0), .b(s_304), .O(gate215inter1));
  and2  gate2677(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate2678(.a(s_304), .O(gate215inter3));
  inv1  gate2679(.a(s_305), .O(gate215inter4));
  nand2 gate2680(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate2681(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate2682(.a(G607), .O(gate215inter7));
  inv1  gate2683(.a(G675), .O(gate215inter8));
  nand2 gate2684(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate2685(.a(s_305), .b(gate215inter3), .O(gate215inter10));
  nor2  gate2686(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate2687(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate2688(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );

  xor2  gate2535(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate2536(.a(gate217inter0), .b(s_284), .O(gate217inter1));
  and2  gate2537(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate2538(.a(s_284), .O(gate217inter3));
  inv1  gate2539(.a(s_285), .O(gate217inter4));
  nand2 gate2540(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate2541(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate2542(.a(G622), .O(gate217inter7));
  inv1  gate2543(.a(G678), .O(gate217inter8));
  nand2 gate2544(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate2545(.a(s_285), .b(gate217inter3), .O(gate217inter10));
  nor2  gate2546(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate2547(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate2548(.a(gate217inter12), .b(gate217inter1), .O(G698));

  xor2  gate1191(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate1192(.a(gate218inter0), .b(s_92), .O(gate218inter1));
  and2  gate1193(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate1194(.a(s_92), .O(gate218inter3));
  inv1  gate1195(.a(s_93), .O(gate218inter4));
  nand2 gate1196(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate1197(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate1198(.a(G627), .O(gate218inter7));
  inv1  gate1199(.a(G678), .O(gate218inter8));
  nand2 gate1200(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate1201(.a(s_93), .b(gate218inter3), .O(gate218inter10));
  nor2  gate1202(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate1203(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate1204(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate2885(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate2886(.a(gate220inter0), .b(s_334), .O(gate220inter1));
  and2  gate2887(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate2888(.a(s_334), .O(gate220inter3));
  inv1  gate2889(.a(s_335), .O(gate220inter4));
  nand2 gate2890(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate2891(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate2892(.a(G637), .O(gate220inter7));
  inv1  gate2893(.a(G681), .O(gate220inter8));
  nand2 gate2894(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate2895(.a(s_335), .b(gate220inter3), .O(gate220inter10));
  nor2  gate2896(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate2897(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate2898(.a(gate220inter12), .b(gate220inter1), .O(G701));

  xor2  gate1947(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate1948(.a(gate221inter0), .b(s_200), .O(gate221inter1));
  and2  gate1949(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate1950(.a(s_200), .O(gate221inter3));
  inv1  gate1951(.a(s_201), .O(gate221inter4));
  nand2 gate1952(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate1953(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate1954(.a(G622), .O(gate221inter7));
  inv1  gate1955(.a(G684), .O(gate221inter8));
  nand2 gate1956(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate1957(.a(s_201), .b(gate221inter3), .O(gate221inter10));
  nor2  gate1958(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate1959(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate1960(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate2479(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate2480(.a(gate223inter0), .b(s_276), .O(gate223inter1));
  and2  gate2481(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate2482(.a(s_276), .O(gate223inter3));
  inv1  gate2483(.a(s_277), .O(gate223inter4));
  nand2 gate2484(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate2485(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate2486(.a(G627), .O(gate223inter7));
  inv1  gate2487(.a(G687), .O(gate223inter8));
  nand2 gate2488(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate2489(.a(s_277), .b(gate223inter3), .O(gate223inter10));
  nor2  gate2490(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate2491(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate2492(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate1275(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate1276(.a(gate226inter0), .b(s_104), .O(gate226inter1));
  and2  gate1277(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate1278(.a(s_104), .O(gate226inter3));
  inv1  gate1279(.a(s_105), .O(gate226inter4));
  nand2 gate1280(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate1281(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate1282(.a(G692), .O(gate226inter7));
  inv1  gate1283(.a(G693), .O(gate226inter8));
  nand2 gate1284(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate1285(.a(s_105), .b(gate226inter3), .O(gate226inter10));
  nor2  gate1286(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate1287(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate1288(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate575(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate576(.a(gate228inter0), .b(s_4), .O(gate228inter1));
  and2  gate577(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate578(.a(s_4), .O(gate228inter3));
  inv1  gate579(.a(s_5), .O(gate228inter4));
  nand2 gate580(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate581(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate582(.a(G696), .O(gate228inter7));
  inv1  gate583(.a(G697), .O(gate228inter8));
  nand2 gate584(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate585(.a(s_5), .b(gate228inter3), .O(gate228inter10));
  nor2  gate586(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate587(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate588(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );

  xor2  gate3011(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate3012(.a(gate232inter0), .b(s_352), .O(gate232inter1));
  and2  gate3013(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate3014(.a(s_352), .O(gate232inter3));
  inv1  gate3015(.a(s_353), .O(gate232inter4));
  nand2 gate3016(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate3017(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate3018(.a(G704), .O(gate232inter7));
  inv1  gate3019(.a(G705), .O(gate232inter8));
  nand2 gate3020(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate3021(.a(s_353), .b(gate232inter3), .O(gate232inter10));
  nor2  gate3022(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate3023(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate3024(.a(gate232inter12), .b(gate232inter1), .O(G727));
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate1415(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate1416(.a(gate237inter0), .b(s_124), .O(gate237inter1));
  and2  gate1417(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate1418(.a(s_124), .O(gate237inter3));
  inv1  gate1419(.a(s_125), .O(gate237inter4));
  nand2 gate1420(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1421(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1422(.a(G254), .O(gate237inter7));
  inv1  gate1423(.a(G706), .O(gate237inter8));
  nand2 gate1424(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1425(.a(s_125), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1426(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1427(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1428(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate2283(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate2284(.a(gate240inter0), .b(s_248), .O(gate240inter1));
  and2  gate2285(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate2286(.a(s_248), .O(gate240inter3));
  inv1  gate2287(.a(s_249), .O(gate240inter4));
  nand2 gate2288(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate2289(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate2290(.a(G263), .O(gate240inter7));
  inv1  gate2291(.a(G715), .O(gate240inter8));
  nand2 gate2292(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate2293(.a(s_249), .b(gate240inter3), .O(gate240inter10));
  nor2  gate2294(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate2295(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate2296(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate2031(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate2032(.a(gate245inter0), .b(s_212), .O(gate245inter1));
  and2  gate2033(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate2034(.a(s_212), .O(gate245inter3));
  inv1  gate2035(.a(s_213), .O(gate245inter4));
  nand2 gate2036(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate2037(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate2038(.a(G248), .O(gate245inter7));
  inv1  gate2039(.a(G736), .O(gate245inter8));
  nand2 gate2040(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate2041(.a(s_213), .b(gate245inter3), .O(gate245inter10));
  nor2  gate2042(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate2043(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate2044(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );

  xor2  gate1639(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate1640(.a(gate247inter0), .b(s_156), .O(gate247inter1));
  and2  gate1641(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate1642(.a(s_156), .O(gate247inter3));
  inv1  gate1643(.a(s_157), .O(gate247inter4));
  nand2 gate1644(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate1645(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate1646(.a(G251), .O(gate247inter7));
  inv1  gate1647(.a(G739), .O(gate247inter8));
  nand2 gate1648(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate1649(.a(s_157), .b(gate247inter3), .O(gate247inter10));
  nor2  gate1650(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate1651(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate1652(.a(gate247inter12), .b(gate247inter1), .O(G760));

  xor2  gate2129(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate2130(.a(gate248inter0), .b(s_226), .O(gate248inter1));
  and2  gate2131(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate2132(.a(s_226), .O(gate248inter3));
  inv1  gate2133(.a(s_227), .O(gate248inter4));
  nand2 gate2134(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate2135(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate2136(.a(G727), .O(gate248inter7));
  inv1  gate2137(.a(G739), .O(gate248inter8));
  nand2 gate2138(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate2139(.a(s_227), .b(gate248inter3), .O(gate248inter10));
  nor2  gate2140(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate2141(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate2142(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate1135(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate1136(.a(gate256inter0), .b(s_84), .O(gate256inter1));
  and2  gate1137(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate1138(.a(s_84), .O(gate256inter3));
  inv1  gate1139(.a(s_85), .O(gate256inter4));
  nand2 gate1140(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate1141(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate1142(.a(G715), .O(gate256inter7));
  inv1  gate1143(.a(G751), .O(gate256inter8));
  nand2 gate1144(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate1145(.a(s_85), .b(gate256inter3), .O(gate256inter10));
  nor2  gate1146(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate1147(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate1148(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate2647(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate2648(.a(gate258inter0), .b(s_300), .O(gate258inter1));
  and2  gate2649(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate2650(.a(s_300), .O(gate258inter3));
  inv1  gate2651(.a(s_301), .O(gate258inter4));
  nand2 gate2652(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate2653(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate2654(.a(G756), .O(gate258inter7));
  inv1  gate2655(.a(G757), .O(gate258inter8));
  nand2 gate2656(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate2657(.a(s_301), .b(gate258inter3), .O(gate258inter10));
  nor2  gate2658(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate2659(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate2660(.a(gate258inter12), .b(gate258inter1), .O(G773));

  xor2  gate2745(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate2746(.a(gate259inter0), .b(s_314), .O(gate259inter1));
  and2  gate2747(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate2748(.a(s_314), .O(gate259inter3));
  inv1  gate2749(.a(s_315), .O(gate259inter4));
  nand2 gate2750(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate2751(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate2752(.a(G758), .O(gate259inter7));
  inv1  gate2753(.a(G759), .O(gate259inter8));
  nand2 gate2754(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate2755(.a(s_315), .b(gate259inter3), .O(gate259inter10));
  nor2  gate2756(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate2757(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate2758(.a(gate259inter12), .b(gate259inter1), .O(G776));

  xor2  gate1835(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate1836(.a(gate260inter0), .b(s_184), .O(gate260inter1));
  and2  gate1837(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate1838(.a(s_184), .O(gate260inter3));
  inv1  gate1839(.a(s_185), .O(gate260inter4));
  nand2 gate1840(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate1841(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate1842(.a(G760), .O(gate260inter7));
  inv1  gate1843(.a(G761), .O(gate260inter8));
  nand2 gate1844(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate1845(.a(s_185), .b(gate260inter3), .O(gate260inter10));
  nor2  gate1846(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate1847(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate1848(.a(gate260inter12), .b(gate260inter1), .O(G779));

  xor2  gate1303(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate1304(.a(gate261inter0), .b(s_108), .O(gate261inter1));
  and2  gate1305(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate1306(.a(s_108), .O(gate261inter3));
  inv1  gate1307(.a(s_109), .O(gate261inter4));
  nand2 gate1308(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate1309(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate1310(.a(G762), .O(gate261inter7));
  inv1  gate1311(.a(G763), .O(gate261inter8));
  nand2 gate1312(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate1313(.a(s_109), .b(gate261inter3), .O(gate261inter10));
  nor2  gate1314(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate1315(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate1316(.a(gate261inter12), .b(gate261inter1), .O(G782));
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate2115(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate2116(.a(gate265inter0), .b(s_224), .O(gate265inter1));
  and2  gate2117(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate2118(.a(s_224), .O(gate265inter3));
  inv1  gate2119(.a(s_225), .O(gate265inter4));
  nand2 gate2120(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate2121(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate2122(.a(G642), .O(gate265inter7));
  inv1  gate2123(.a(G770), .O(gate265inter8));
  nand2 gate2124(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate2125(.a(s_225), .b(gate265inter3), .O(gate265inter10));
  nor2  gate2126(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate2127(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate2128(.a(gate265inter12), .b(gate265inter1), .O(G794));

  xor2  gate2269(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate2270(.a(gate266inter0), .b(s_246), .O(gate266inter1));
  and2  gate2271(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate2272(.a(s_246), .O(gate266inter3));
  inv1  gate2273(.a(s_247), .O(gate266inter4));
  nand2 gate2274(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate2275(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate2276(.a(G645), .O(gate266inter7));
  inv1  gate2277(.a(G773), .O(gate266inter8));
  nand2 gate2278(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate2279(.a(s_247), .b(gate266inter3), .O(gate266inter10));
  nor2  gate2280(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate2281(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate2282(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate1961(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate1962(.a(gate274inter0), .b(s_202), .O(gate274inter1));
  and2  gate1963(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate1964(.a(s_202), .O(gate274inter3));
  inv1  gate1965(.a(s_203), .O(gate274inter4));
  nand2 gate1966(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate1967(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate1968(.a(G770), .O(gate274inter7));
  inv1  gate1969(.a(G794), .O(gate274inter8));
  nand2 gate1970(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate1971(.a(s_203), .b(gate274inter3), .O(gate274inter10));
  nor2  gate1972(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate1973(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate1974(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate1051(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate1052(.a(gate276inter0), .b(s_72), .O(gate276inter1));
  and2  gate1053(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate1054(.a(s_72), .O(gate276inter3));
  inv1  gate1055(.a(s_73), .O(gate276inter4));
  nand2 gate1056(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate1057(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate1058(.a(G773), .O(gate276inter7));
  inv1  gate1059(.a(G797), .O(gate276inter8));
  nand2 gate1060(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate1061(.a(s_73), .b(gate276inter3), .O(gate276inter10));
  nor2  gate1062(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate1063(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate1064(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate2829(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate2830(.a(gate278inter0), .b(s_326), .O(gate278inter1));
  and2  gate2831(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate2832(.a(s_326), .O(gate278inter3));
  inv1  gate2833(.a(s_327), .O(gate278inter4));
  nand2 gate2834(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate2835(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate2836(.a(G776), .O(gate278inter7));
  inv1  gate2837(.a(G800), .O(gate278inter8));
  nand2 gate2838(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate2839(.a(s_327), .b(gate278inter3), .O(gate278inter10));
  nor2  gate2840(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate2841(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate2842(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate1541(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate1542(.a(gate280inter0), .b(s_142), .O(gate280inter1));
  and2  gate1543(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate1544(.a(s_142), .O(gate280inter3));
  inv1  gate1545(.a(s_143), .O(gate280inter4));
  nand2 gate1546(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate1547(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate1548(.a(G779), .O(gate280inter7));
  inv1  gate1549(.a(G803), .O(gate280inter8));
  nand2 gate1550(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate1551(.a(s_143), .b(gate280inter3), .O(gate280inter10));
  nor2  gate1552(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate1553(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate1554(.a(gate280inter12), .b(gate280inter1), .O(G825));

  xor2  gate1737(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate1738(.a(gate281inter0), .b(s_170), .O(gate281inter1));
  and2  gate1739(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate1740(.a(s_170), .O(gate281inter3));
  inv1  gate1741(.a(s_171), .O(gate281inter4));
  nand2 gate1742(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate1743(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate1744(.a(G654), .O(gate281inter7));
  inv1  gate1745(.a(G806), .O(gate281inter8));
  nand2 gate1746(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate1747(.a(s_171), .b(gate281inter3), .O(gate281inter10));
  nor2  gate1748(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate1749(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate1750(.a(gate281inter12), .b(gate281inter1), .O(G826));

  xor2  gate2899(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate2900(.a(gate282inter0), .b(s_336), .O(gate282inter1));
  and2  gate2901(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate2902(.a(s_336), .O(gate282inter3));
  inv1  gate2903(.a(s_337), .O(gate282inter4));
  nand2 gate2904(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate2905(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate2906(.a(G782), .O(gate282inter7));
  inv1  gate2907(.a(G806), .O(gate282inter8));
  nand2 gate2908(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate2909(.a(s_337), .b(gate282inter3), .O(gate282inter10));
  nor2  gate2910(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate2911(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate2912(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate561(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate562(.a(gate285inter0), .b(s_2), .O(gate285inter1));
  and2  gate563(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate564(.a(s_2), .O(gate285inter3));
  inv1  gate565(.a(s_3), .O(gate285inter4));
  nand2 gate566(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate567(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate568(.a(G660), .O(gate285inter7));
  inv1  gate569(.a(G812), .O(gate285inter8));
  nand2 gate570(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate571(.a(s_3), .b(gate285inter3), .O(gate285inter10));
  nor2  gate572(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate573(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate574(.a(gate285inter12), .b(gate285inter1), .O(G830));

  xor2  gate547(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate548(.a(gate286inter0), .b(s_0), .O(gate286inter1));
  and2  gate549(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate550(.a(s_0), .O(gate286inter3));
  inv1  gate551(.a(s_1), .O(gate286inter4));
  nand2 gate552(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate553(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate554(.a(G788), .O(gate286inter7));
  inv1  gate555(.a(G812), .O(gate286inter8));
  nand2 gate556(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate557(.a(s_1), .b(gate286inter3), .O(gate286inter10));
  nor2  gate558(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate559(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate560(.a(gate286inter12), .b(gate286inter1), .O(G831));
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate715(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate716(.a(gate288inter0), .b(s_24), .O(gate288inter1));
  and2  gate717(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate718(.a(s_24), .O(gate288inter3));
  inv1  gate719(.a(s_25), .O(gate288inter4));
  nand2 gate720(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate721(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate722(.a(G791), .O(gate288inter7));
  inv1  gate723(.a(G815), .O(gate288inter8));
  nand2 gate724(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate725(.a(s_25), .b(gate288inter3), .O(gate288inter10));
  nor2  gate726(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate727(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate728(.a(gate288inter12), .b(gate288inter1), .O(G833));

  xor2  gate1905(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate1906(.a(gate289inter0), .b(s_194), .O(gate289inter1));
  and2  gate1907(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate1908(.a(s_194), .O(gate289inter3));
  inv1  gate1909(.a(s_195), .O(gate289inter4));
  nand2 gate1910(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate1911(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate1912(.a(G818), .O(gate289inter7));
  inv1  gate1913(.a(G819), .O(gate289inter8));
  nand2 gate1914(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate1915(.a(s_195), .b(gate289inter3), .O(gate289inter10));
  nor2  gate1916(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate1917(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate1918(.a(gate289inter12), .b(gate289inter1), .O(G834));

  xor2  gate2493(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate2494(.a(gate290inter0), .b(s_278), .O(gate290inter1));
  and2  gate2495(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate2496(.a(s_278), .O(gate290inter3));
  inv1  gate2497(.a(s_279), .O(gate290inter4));
  nand2 gate2498(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate2499(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate2500(.a(G820), .O(gate290inter7));
  inv1  gate2501(.a(G821), .O(gate290inter8));
  nand2 gate2502(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate2503(.a(s_279), .b(gate290inter3), .O(gate290inter10));
  nor2  gate2504(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate2505(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate2506(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate2857(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate2858(.a(gate294inter0), .b(s_330), .O(gate294inter1));
  and2  gate2859(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate2860(.a(s_330), .O(gate294inter3));
  inv1  gate2861(.a(s_331), .O(gate294inter4));
  nand2 gate2862(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate2863(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate2864(.a(G832), .O(gate294inter7));
  inv1  gate2865(.a(G833), .O(gate294inter8));
  nand2 gate2866(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate2867(.a(s_331), .b(gate294inter3), .O(gate294inter10));
  nor2  gate2868(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate2869(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate2870(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate897(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate898(.a(gate296inter0), .b(s_50), .O(gate296inter1));
  and2  gate899(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate900(.a(s_50), .O(gate296inter3));
  inv1  gate901(.a(s_51), .O(gate296inter4));
  nand2 gate902(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate903(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate904(.a(G826), .O(gate296inter7));
  inv1  gate905(.a(G827), .O(gate296inter8));
  nand2 gate906(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate907(.a(s_51), .b(gate296inter3), .O(gate296inter10));
  nor2  gate908(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate909(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate910(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate3039(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate3040(.a(gate388inter0), .b(s_356), .O(gate388inter1));
  and2  gate3041(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate3042(.a(s_356), .O(gate388inter3));
  inv1  gate3043(.a(s_357), .O(gate388inter4));
  nand2 gate3044(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate3045(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate3046(.a(G2), .O(gate388inter7));
  inv1  gate3047(.a(G1039), .O(gate388inter8));
  nand2 gate3048(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate3049(.a(s_357), .b(gate388inter3), .O(gate388inter10));
  nor2  gate3050(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate3051(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate3052(.a(gate388inter12), .b(gate388inter1), .O(G1135));

  xor2  gate2997(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate2998(.a(gate389inter0), .b(s_350), .O(gate389inter1));
  and2  gate2999(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate3000(.a(s_350), .O(gate389inter3));
  inv1  gate3001(.a(s_351), .O(gate389inter4));
  nand2 gate3002(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate3003(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate3004(.a(G3), .O(gate389inter7));
  inv1  gate3005(.a(G1042), .O(gate389inter8));
  nand2 gate3006(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate3007(.a(s_351), .b(gate389inter3), .O(gate389inter10));
  nor2  gate3008(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate3009(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate3010(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );

  xor2  gate1877(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate1878(.a(gate392inter0), .b(s_190), .O(gate392inter1));
  and2  gate1879(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate1880(.a(s_190), .O(gate392inter3));
  inv1  gate1881(.a(s_191), .O(gate392inter4));
  nand2 gate1882(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate1883(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate1884(.a(G6), .O(gate392inter7));
  inv1  gate1885(.a(G1051), .O(gate392inter8));
  nand2 gate1886(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate1887(.a(s_191), .b(gate392inter3), .O(gate392inter10));
  nor2  gate1888(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate1889(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate1890(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate799(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate800(.a(gate394inter0), .b(s_36), .O(gate394inter1));
  and2  gate801(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate802(.a(s_36), .O(gate394inter3));
  inv1  gate803(.a(s_37), .O(gate394inter4));
  nand2 gate804(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate805(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate806(.a(G8), .O(gate394inter7));
  inv1  gate807(.a(G1057), .O(gate394inter8));
  nand2 gate808(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate809(.a(s_37), .b(gate394inter3), .O(gate394inter10));
  nor2  gate810(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate811(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate812(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate1387(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate1388(.a(gate397inter0), .b(s_120), .O(gate397inter1));
  and2  gate1389(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate1390(.a(s_120), .O(gate397inter3));
  inv1  gate1391(.a(s_121), .O(gate397inter4));
  nand2 gate1392(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate1393(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate1394(.a(G11), .O(gate397inter7));
  inv1  gate1395(.a(G1066), .O(gate397inter8));
  nand2 gate1396(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate1397(.a(s_121), .b(gate397inter3), .O(gate397inter10));
  nor2  gate1398(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate1399(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate1400(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate1079(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate1080(.a(gate400inter0), .b(s_76), .O(gate400inter1));
  and2  gate1081(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate1082(.a(s_76), .O(gate400inter3));
  inv1  gate1083(.a(s_77), .O(gate400inter4));
  nand2 gate1084(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate1085(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate1086(.a(G14), .O(gate400inter7));
  inv1  gate1087(.a(G1075), .O(gate400inter8));
  nand2 gate1088(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate1089(.a(s_77), .b(gate400inter3), .O(gate400inter10));
  nor2  gate1090(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate1091(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate1092(.a(gate400inter12), .b(gate400inter1), .O(G1171));

  xor2  gate1359(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate1360(.a(gate401inter0), .b(s_116), .O(gate401inter1));
  and2  gate1361(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate1362(.a(s_116), .O(gate401inter3));
  inv1  gate1363(.a(s_117), .O(gate401inter4));
  nand2 gate1364(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate1365(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate1366(.a(G15), .O(gate401inter7));
  inv1  gate1367(.a(G1078), .O(gate401inter8));
  nand2 gate1368(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate1369(.a(s_117), .b(gate401inter3), .O(gate401inter10));
  nor2  gate1370(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate1371(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate1372(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );

  xor2  gate1933(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate1934(.a(gate404inter0), .b(s_198), .O(gate404inter1));
  and2  gate1935(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate1936(.a(s_198), .O(gate404inter3));
  inv1  gate1937(.a(s_199), .O(gate404inter4));
  nand2 gate1938(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate1939(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate1940(.a(G18), .O(gate404inter7));
  inv1  gate1941(.a(G1087), .O(gate404inter8));
  nand2 gate1942(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate1943(.a(s_199), .b(gate404inter3), .O(gate404inter10));
  nor2  gate1944(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate1945(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate1946(.a(gate404inter12), .b(gate404inter1), .O(G1183));
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate2815(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate2816(.a(gate406inter0), .b(s_324), .O(gate406inter1));
  and2  gate2817(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate2818(.a(s_324), .O(gate406inter3));
  inv1  gate2819(.a(s_325), .O(gate406inter4));
  nand2 gate2820(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate2821(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate2822(.a(G20), .O(gate406inter7));
  inv1  gate2823(.a(G1093), .O(gate406inter8));
  nand2 gate2824(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate2825(.a(s_325), .b(gate406inter3), .O(gate406inter10));
  nor2  gate2826(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate2827(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate2828(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate2759(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate2760(.a(gate410inter0), .b(s_316), .O(gate410inter1));
  and2  gate2761(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate2762(.a(s_316), .O(gate410inter3));
  inv1  gate2763(.a(s_317), .O(gate410inter4));
  nand2 gate2764(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate2765(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate2766(.a(G24), .O(gate410inter7));
  inv1  gate2767(.a(G1105), .O(gate410inter8));
  nand2 gate2768(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate2769(.a(s_317), .b(gate410inter3), .O(gate410inter10));
  nor2  gate2770(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate2771(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate2772(.a(gate410inter12), .b(gate410inter1), .O(G1201));

  xor2  gate2787(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate2788(.a(gate411inter0), .b(s_320), .O(gate411inter1));
  and2  gate2789(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate2790(.a(s_320), .O(gate411inter3));
  inv1  gate2791(.a(s_321), .O(gate411inter4));
  nand2 gate2792(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate2793(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate2794(.a(G25), .O(gate411inter7));
  inv1  gate2795(.a(G1108), .O(gate411inter8));
  nand2 gate2796(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate2797(.a(s_321), .b(gate411inter3), .O(gate411inter10));
  nor2  gate2798(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate2799(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate2800(.a(gate411inter12), .b(gate411inter1), .O(G1204));

  xor2  gate2451(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate2452(.a(gate412inter0), .b(s_272), .O(gate412inter1));
  and2  gate2453(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate2454(.a(s_272), .O(gate412inter3));
  inv1  gate2455(.a(s_273), .O(gate412inter4));
  nand2 gate2456(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate2457(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate2458(.a(G26), .O(gate412inter7));
  inv1  gate2459(.a(G1111), .O(gate412inter8));
  nand2 gate2460(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate2461(.a(s_273), .b(gate412inter3), .O(gate412inter10));
  nor2  gate2462(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate2463(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate2464(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );

  xor2  gate855(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate856(.a(gate414inter0), .b(s_44), .O(gate414inter1));
  and2  gate857(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate858(.a(s_44), .O(gate414inter3));
  inv1  gate859(.a(s_45), .O(gate414inter4));
  nand2 gate860(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate861(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate862(.a(G28), .O(gate414inter7));
  inv1  gate863(.a(G1117), .O(gate414inter8));
  nand2 gate864(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate865(.a(s_45), .b(gate414inter3), .O(gate414inter10));
  nor2  gate866(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate867(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate868(.a(gate414inter12), .b(gate414inter1), .O(G1213));
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );

  xor2  gate673(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate674(.a(gate416inter0), .b(s_18), .O(gate416inter1));
  and2  gate675(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate676(.a(s_18), .O(gate416inter3));
  inv1  gate677(.a(s_19), .O(gate416inter4));
  nand2 gate678(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate679(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate680(.a(G30), .O(gate416inter7));
  inv1  gate681(.a(G1123), .O(gate416inter8));
  nand2 gate682(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate683(.a(s_19), .b(gate416inter3), .O(gate416inter10));
  nor2  gate684(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate685(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate686(.a(gate416inter12), .b(gate416inter1), .O(G1219));
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate2227(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate2228(.a(gate419inter0), .b(s_240), .O(gate419inter1));
  and2  gate2229(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate2230(.a(s_240), .O(gate419inter3));
  inv1  gate2231(.a(s_241), .O(gate419inter4));
  nand2 gate2232(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate2233(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate2234(.a(G1), .O(gate419inter7));
  inv1  gate2235(.a(G1132), .O(gate419inter8));
  nand2 gate2236(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate2237(.a(s_241), .b(gate419inter3), .O(gate419inter10));
  nor2  gate2238(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate2239(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate2240(.a(gate419inter12), .b(gate419inter1), .O(G1228));

  xor2  gate1247(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1248(.a(gate420inter0), .b(s_100), .O(gate420inter1));
  and2  gate1249(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1250(.a(s_100), .O(gate420inter3));
  inv1  gate1251(.a(s_101), .O(gate420inter4));
  nand2 gate1252(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1253(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1254(.a(G1036), .O(gate420inter7));
  inv1  gate1255(.a(G1132), .O(gate420inter8));
  nand2 gate1256(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1257(.a(s_101), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1258(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1259(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1260(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate1443(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate1444(.a(gate422inter0), .b(s_128), .O(gate422inter1));
  and2  gate1445(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate1446(.a(s_128), .O(gate422inter3));
  inv1  gate1447(.a(s_129), .O(gate422inter4));
  nand2 gate1448(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate1449(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate1450(.a(G1039), .O(gate422inter7));
  inv1  gate1451(.a(G1135), .O(gate422inter8));
  nand2 gate1452(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate1453(.a(s_129), .b(gate422inter3), .O(gate422inter10));
  nor2  gate1454(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate1455(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate1456(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );

  xor2  gate1023(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate1024(.a(gate427inter0), .b(s_68), .O(gate427inter1));
  and2  gate1025(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate1026(.a(s_68), .O(gate427inter3));
  inv1  gate1027(.a(s_69), .O(gate427inter4));
  nand2 gate1028(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate1029(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate1030(.a(G5), .O(gate427inter7));
  inv1  gate1031(.a(G1144), .O(gate427inter8));
  nand2 gate1032(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate1033(.a(s_69), .b(gate427inter3), .O(gate427inter10));
  nor2  gate1034(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate1035(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate1036(.a(gate427inter12), .b(gate427inter1), .O(G1236));

  xor2  gate1807(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate1808(.a(gate428inter0), .b(s_180), .O(gate428inter1));
  and2  gate1809(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate1810(.a(s_180), .O(gate428inter3));
  inv1  gate1811(.a(s_181), .O(gate428inter4));
  nand2 gate1812(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate1813(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate1814(.a(G1048), .O(gate428inter7));
  inv1  gate1815(.a(G1144), .O(gate428inter8));
  nand2 gate1816(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate1817(.a(s_181), .b(gate428inter3), .O(gate428inter10));
  nor2  gate1818(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate1819(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate1820(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate1681(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate1682(.a(gate431inter0), .b(s_162), .O(gate431inter1));
  and2  gate1683(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate1684(.a(s_162), .O(gate431inter3));
  inv1  gate1685(.a(s_163), .O(gate431inter4));
  nand2 gate1686(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate1687(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate1688(.a(G7), .O(gate431inter7));
  inv1  gate1689(.a(G1150), .O(gate431inter8));
  nand2 gate1690(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate1691(.a(s_163), .b(gate431inter3), .O(gate431inter10));
  nor2  gate1692(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate1693(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate1694(.a(gate431inter12), .b(gate431inter1), .O(G1240));

  xor2  gate2213(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate2214(.a(gate432inter0), .b(s_238), .O(gate432inter1));
  and2  gate2215(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate2216(.a(s_238), .O(gate432inter3));
  inv1  gate2217(.a(s_239), .O(gate432inter4));
  nand2 gate2218(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate2219(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate2220(.a(G1054), .O(gate432inter7));
  inv1  gate2221(.a(G1150), .O(gate432inter8));
  nand2 gate2222(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate2223(.a(s_239), .b(gate432inter3), .O(gate432inter10));
  nor2  gate2224(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate2225(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate2226(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate981(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate982(.a(gate435inter0), .b(s_62), .O(gate435inter1));
  and2  gate983(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate984(.a(s_62), .O(gate435inter3));
  inv1  gate985(.a(s_63), .O(gate435inter4));
  nand2 gate986(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate987(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate988(.a(G9), .O(gate435inter7));
  inv1  gate989(.a(G1156), .O(gate435inter8));
  nand2 gate990(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate991(.a(s_63), .b(gate435inter3), .O(gate435inter10));
  nor2  gate992(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate993(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate994(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate911(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate912(.a(gate439inter0), .b(s_52), .O(gate439inter1));
  and2  gate913(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate914(.a(s_52), .O(gate439inter3));
  inv1  gate915(.a(s_53), .O(gate439inter4));
  nand2 gate916(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate917(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate918(.a(G11), .O(gate439inter7));
  inv1  gate919(.a(G1162), .O(gate439inter8));
  nand2 gate920(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate921(.a(s_53), .b(gate439inter3), .O(gate439inter10));
  nor2  gate922(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate923(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate924(.a(gate439inter12), .b(gate439inter1), .O(G1248));

  xor2  gate2003(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate2004(.a(gate440inter0), .b(s_208), .O(gate440inter1));
  and2  gate2005(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate2006(.a(s_208), .O(gate440inter3));
  inv1  gate2007(.a(s_209), .O(gate440inter4));
  nand2 gate2008(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate2009(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate2010(.a(G1066), .O(gate440inter7));
  inv1  gate2011(.a(G1162), .O(gate440inter8));
  nand2 gate2012(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate2013(.a(s_209), .b(gate440inter3), .O(gate440inter10));
  nor2  gate2014(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate2015(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate2016(.a(gate440inter12), .b(gate440inter1), .O(G1249));

  xor2  gate2507(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate2508(.a(gate441inter0), .b(s_280), .O(gate441inter1));
  and2  gate2509(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate2510(.a(s_280), .O(gate441inter3));
  inv1  gate2511(.a(s_281), .O(gate441inter4));
  nand2 gate2512(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate2513(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate2514(.a(G12), .O(gate441inter7));
  inv1  gate2515(.a(G1165), .O(gate441inter8));
  nand2 gate2516(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate2517(.a(s_281), .b(gate441inter3), .O(gate441inter10));
  nor2  gate2518(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate2519(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate2520(.a(gate441inter12), .b(gate441inter1), .O(G1250));

  xor2  gate2955(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate2956(.a(gate442inter0), .b(s_344), .O(gate442inter1));
  and2  gate2957(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate2958(.a(s_344), .O(gate442inter3));
  inv1  gate2959(.a(s_345), .O(gate442inter4));
  nand2 gate2960(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate2961(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate2962(.a(G1069), .O(gate442inter7));
  inv1  gate2963(.a(G1165), .O(gate442inter8));
  nand2 gate2964(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate2965(.a(s_345), .b(gate442inter3), .O(gate442inter10));
  nor2  gate2966(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate2967(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate2968(.a(gate442inter12), .b(gate442inter1), .O(G1251));

  xor2  gate3025(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate3026(.a(gate443inter0), .b(s_354), .O(gate443inter1));
  and2  gate3027(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate3028(.a(s_354), .O(gate443inter3));
  inv1  gate3029(.a(s_355), .O(gate443inter4));
  nand2 gate3030(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate3031(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate3032(.a(G13), .O(gate443inter7));
  inv1  gate3033(.a(G1168), .O(gate443inter8));
  nand2 gate3034(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate3035(.a(s_355), .b(gate443inter3), .O(gate443inter10));
  nor2  gate3036(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate3037(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate3038(.a(gate443inter12), .b(gate443inter1), .O(G1252));

  xor2  gate2773(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate2774(.a(gate444inter0), .b(s_318), .O(gate444inter1));
  and2  gate2775(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate2776(.a(s_318), .O(gate444inter3));
  inv1  gate2777(.a(s_319), .O(gate444inter4));
  nand2 gate2778(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate2779(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate2780(.a(G1072), .O(gate444inter7));
  inv1  gate2781(.a(G1168), .O(gate444inter8));
  nand2 gate2782(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate2783(.a(s_319), .b(gate444inter3), .O(gate444inter10));
  nor2  gate2784(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate2785(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate2786(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );

  xor2  gate1065(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate1066(.a(gate446inter0), .b(s_74), .O(gate446inter1));
  and2  gate1067(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate1068(.a(s_74), .O(gate446inter3));
  inv1  gate1069(.a(s_75), .O(gate446inter4));
  nand2 gate1070(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate1071(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate1072(.a(G1075), .O(gate446inter7));
  inv1  gate1073(.a(G1171), .O(gate446inter8));
  nand2 gate1074(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate1075(.a(s_75), .b(gate446inter3), .O(gate446inter10));
  nor2  gate1076(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate1077(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate1078(.a(gate446inter12), .b(gate446inter1), .O(G1255));
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );

  xor2  gate1163(.a(G1183), .b(G1087), .O(gate454inter0));
  nand2 gate1164(.a(gate454inter0), .b(s_88), .O(gate454inter1));
  and2  gate1165(.a(G1183), .b(G1087), .O(gate454inter2));
  inv1  gate1166(.a(s_88), .O(gate454inter3));
  inv1  gate1167(.a(s_89), .O(gate454inter4));
  nand2 gate1168(.a(gate454inter4), .b(gate454inter3), .O(gate454inter5));
  nor2  gate1169(.a(gate454inter5), .b(gate454inter2), .O(gate454inter6));
  inv1  gate1170(.a(G1087), .O(gate454inter7));
  inv1  gate1171(.a(G1183), .O(gate454inter8));
  nand2 gate1172(.a(gate454inter8), .b(gate454inter7), .O(gate454inter9));
  nand2 gate1173(.a(s_89), .b(gate454inter3), .O(gate454inter10));
  nor2  gate1174(.a(gate454inter10), .b(gate454inter9), .O(gate454inter11));
  nor2  gate1175(.a(gate454inter11), .b(gate454inter6), .O(gate454inter12));
  nand2 gate1176(.a(gate454inter12), .b(gate454inter1), .O(G1263));

  xor2  gate2619(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate2620(.a(gate455inter0), .b(s_296), .O(gate455inter1));
  and2  gate2621(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate2622(.a(s_296), .O(gate455inter3));
  inv1  gate2623(.a(s_297), .O(gate455inter4));
  nand2 gate2624(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate2625(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate2626(.a(G19), .O(gate455inter7));
  inv1  gate2627(.a(G1186), .O(gate455inter8));
  nand2 gate2628(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate2629(.a(s_297), .b(gate455inter3), .O(gate455inter10));
  nor2  gate2630(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate2631(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate2632(.a(gate455inter12), .b(gate455inter1), .O(G1264));
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate1569(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate1570(.a(gate463inter0), .b(s_146), .O(gate463inter1));
  and2  gate1571(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate1572(.a(s_146), .O(gate463inter3));
  inv1  gate1573(.a(s_147), .O(gate463inter4));
  nand2 gate1574(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate1575(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate1576(.a(G23), .O(gate463inter7));
  inv1  gate1577(.a(G1198), .O(gate463inter8));
  nand2 gate1578(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate1579(.a(s_147), .b(gate463inter3), .O(gate463inter10));
  nor2  gate1580(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate1581(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate1582(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate1513(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate1514(.a(gate465inter0), .b(s_138), .O(gate465inter1));
  and2  gate1515(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate1516(.a(s_138), .O(gate465inter3));
  inv1  gate1517(.a(s_139), .O(gate465inter4));
  nand2 gate1518(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate1519(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate1520(.a(G24), .O(gate465inter7));
  inv1  gate1521(.a(G1201), .O(gate465inter8));
  nand2 gate1522(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate1523(.a(s_139), .b(gate465inter3), .O(gate465inter10));
  nor2  gate1524(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate1525(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate1526(.a(gate465inter12), .b(gate465inter1), .O(G1274));

  xor2  gate2171(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate2172(.a(gate466inter0), .b(s_232), .O(gate466inter1));
  and2  gate2173(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate2174(.a(s_232), .O(gate466inter3));
  inv1  gate2175(.a(s_233), .O(gate466inter4));
  nand2 gate2176(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate2177(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate2178(.a(G1105), .O(gate466inter7));
  inv1  gate2179(.a(G1201), .O(gate466inter8));
  nand2 gate2180(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate2181(.a(s_233), .b(gate466inter3), .O(gate466inter10));
  nor2  gate2182(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate2183(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate2184(.a(gate466inter12), .b(gate466inter1), .O(G1275));

  xor2  gate1499(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate1500(.a(gate467inter0), .b(s_136), .O(gate467inter1));
  and2  gate1501(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate1502(.a(s_136), .O(gate467inter3));
  inv1  gate1503(.a(s_137), .O(gate467inter4));
  nand2 gate1504(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate1505(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate1506(.a(G25), .O(gate467inter7));
  inv1  gate1507(.a(G1204), .O(gate467inter8));
  nand2 gate1508(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate1509(.a(s_137), .b(gate467inter3), .O(gate467inter10));
  nor2  gate1510(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate1511(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate1512(.a(gate467inter12), .b(gate467inter1), .O(G1276));

  xor2  gate1093(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate1094(.a(gate468inter0), .b(s_78), .O(gate468inter1));
  and2  gate1095(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate1096(.a(s_78), .O(gate468inter3));
  inv1  gate1097(.a(s_79), .O(gate468inter4));
  nand2 gate1098(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate1099(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate1100(.a(G1108), .O(gate468inter7));
  inv1  gate1101(.a(G1204), .O(gate468inter8));
  nand2 gate1102(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate1103(.a(s_79), .b(gate468inter3), .O(gate468inter10));
  nor2  gate1104(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate1105(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate1106(.a(gate468inter12), .b(gate468inter1), .O(G1277));

  xor2  gate687(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate688(.a(gate469inter0), .b(s_20), .O(gate469inter1));
  and2  gate689(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate690(.a(s_20), .O(gate469inter3));
  inv1  gate691(.a(s_21), .O(gate469inter4));
  nand2 gate692(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate693(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate694(.a(G26), .O(gate469inter7));
  inv1  gate695(.a(G1207), .O(gate469inter8));
  nand2 gate696(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate697(.a(s_21), .b(gate469inter3), .O(gate469inter10));
  nor2  gate698(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate699(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate700(.a(gate469inter12), .b(gate469inter1), .O(G1278));
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate617(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate618(.a(gate472inter0), .b(s_10), .O(gate472inter1));
  and2  gate619(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate620(.a(s_10), .O(gate472inter3));
  inv1  gate621(.a(s_11), .O(gate472inter4));
  nand2 gate622(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate623(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate624(.a(G1114), .O(gate472inter7));
  inv1  gate625(.a(G1210), .O(gate472inter8));
  nand2 gate626(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate627(.a(s_11), .b(gate472inter3), .O(gate472inter10));
  nor2  gate628(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate629(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate630(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate2437(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate2438(.a(gate476inter0), .b(s_270), .O(gate476inter1));
  and2  gate2439(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate2440(.a(s_270), .O(gate476inter3));
  inv1  gate2441(.a(s_271), .O(gate476inter4));
  nand2 gate2442(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate2443(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate2444(.a(G1120), .O(gate476inter7));
  inv1  gate2445(.a(G1216), .O(gate476inter8));
  nand2 gate2446(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate2447(.a(s_271), .b(gate476inter3), .O(gate476inter10));
  nor2  gate2448(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate2449(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate2450(.a(gate476inter12), .b(gate476inter1), .O(G1285));

  xor2  gate2521(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate2522(.a(gate477inter0), .b(s_282), .O(gate477inter1));
  and2  gate2523(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate2524(.a(s_282), .O(gate477inter3));
  inv1  gate2525(.a(s_283), .O(gate477inter4));
  nand2 gate2526(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate2527(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate2528(.a(G30), .O(gate477inter7));
  inv1  gate2529(.a(G1219), .O(gate477inter8));
  nand2 gate2530(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate2531(.a(s_283), .b(gate477inter3), .O(gate477inter10));
  nor2  gate2532(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate2533(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate2534(.a(gate477inter12), .b(gate477inter1), .O(G1286));

  xor2  gate925(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate926(.a(gate478inter0), .b(s_54), .O(gate478inter1));
  and2  gate927(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate928(.a(s_54), .O(gate478inter3));
  inv1  gate929(.a(s_55), .O(gate478inter4));
  nand2 gate930(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate931(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate932(.a(G1123), .O(gate478inter7));
  inv1  gate933(.a(G1219), .O(gate478inter8));
  nand2 gate934(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate935(.a(s_55), .b(gate478inter3), .O(gate478inter10));
  nor2  gate936(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate937(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate938(.a(gate478inter12), .b(gate478inter1), .O(G1287));

  xor2  gate1345(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate1346(.a(gate479inter0), .b(s_114), .O(gate479inter1));
  and2  gate1347(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate1348(.a(s_114), .O(gate479inter3));
  inv1  gate1349(.a(s_115), .O(gate479inter4));
  nand2 gate1350(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate1351(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate1352(.a(G31), .O(gate479inter7));
  inv1  gate1353(.a(G1222), .O(gate479inter8));
  nand2 gate1354(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate1355(.a(s_115), .b(gate479inter3), .O(gate479inter10));
  nor2  gate1356(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate1357(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate1358(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate2661(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate2662(.a(gate486inter0), .b(s_302), .O(gate486inter1));
  and2  gate2663(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate2664(.a(s_302), .O(gate486inter3));
  inv1  gate2665(.a(s_303), .O(gate486inter4));
  nand2 gate2666(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate2667(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate2668(.a(G1234), .O(gate486inter7));
  inv1  gate2669(.a(G1235), .O(gate486inter8));
  nand2 gate2670(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate2671(.a(s_303), .b(gate486inter3), .O(gate486inter10));
  nor2  gate2672(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate2673(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate2674(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate645(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate646(.a(gate488inter0), .b(s_14), .O(gate488inter1));
  and2  gate647(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate648(.a(s_14), .O(gate488inter3));
  inv1  gate649(.a(s_15), .O(gate488inter4));
  nand2 gate650(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate651(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate652(.a(G1238), .O(gate488inter7));
  inv1  gate653(.a(G1239), .O(gate488inter8));
  nand2 gate654(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate655(.a(s_15), .b(gate488inter3), .O(gate488inter10));
  nor2  gate656(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate657(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate658(.a(gate488inter12), .b(gate488inter1), .O(G1297));

  xor2  gate939(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate940(.a(gate489inter0), .b(s_56), .O(gate489inter1));
  and2  gate941(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate942(.a(s_56), .O(gate489inter3));
  inv1  gate943(.a(s_57), .O(gate489inter4));
  nand2 gate944(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate945(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate946(.a(G1240), .O(gate489inter7));
  inv1  gate947(.a(G1241), .O(gate489inter8));
  nand2 gate948(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate949(.a(s_57), .b(gate489inter3), .O(gate489inter10));
  nor2  gate950(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate951(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate952(.a(gate489inter12), .b(gate489inter1), .O(G1298));

  xor2  gate1289(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate1290(.a(gate490inter0), .b(s_106), .O(gate490inter1));
  and2  gate1291(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate1292(.a(s_106), .O(gate490inter3));
  inv1  gate1293(.a(s_107), .O(gate490inter4));
  nand2 gate1294(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate1295(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate1296(.a(G1242), .O(gate490inter7));
  inv1  gate1297(.a(G1243), .O(gate490inter8));
  nand2 gate1298(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate1299(.a(s_107), .b(gate490inter3), .O(gate490inter10));
  nor2  gate1300(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate1301(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate1302(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate2633(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate2634(.a(gate494inter0), .b(s_298), .O(gate494inter1));
  and2  gate2635(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate2636(.a(s_298), .O(gate494inter3));
  inv1  gate2637(.a(s_299), .O(gate494inter4));
  nand2 gate2638(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate2639(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate2640(.a(G1250), .O(gate494inter7));
  inv1  gate2641(.a(G1251), .O(gate494inter8));
  nand2 gate2642(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate2643(.a(s_299), .b(gate494inter3), .O(gate494inter10));
  nor2  gate2644(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate2645(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate2646(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate743(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate744(.a(gate497inter0), .b(s_28), .O(gate497inter1));
  and2  gate745(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate746(.a(s_28), .O(gate497inter3));
  inv1  gate747(.a(s_29), .O(gate497inter4));
  nand2 gate748(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate749(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate750(.a(G1256), .O(gate497inter7));
  inv1  gate751(.a(G1257), .O(gate497inter8));
  nand2 gate752(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate753(.a(s_29), .b(gate497inter3), .O(gate497inter10));
  nor2  gate754(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate755(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate756(.a(gate497inter12), .b(gate497inter1), .O(G1306));

  xor2  gate2423(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate2424(.a(gate498inter0), .b(s_268), .O(gate498inter1));
  and2  gate2425(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate2426(.a(s_268), .O(gate498inter3));
  inv1  gate2427(.a(s_269), .O(gate498inter4));
  nand2 gate2428(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate2429(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate2430(.a(G1258), .O(gate498inter7));
  inv1  gate2431(.a(G1259), .O(gate498inter8));
  nand2 gate2432(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate2433(.a(s_269), .b(gate498inter3), .O(gate498inter10));
  nor2  gate2434(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate2435(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate2436(.a(gate498inter12), .b(gate498inter1), .O(G1307));
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );

  xor2  gate2045(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate2046(.a(gate507inter0), .b(s_214), .O(gate507inter1));
  and2  gate2047(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate2048(.a(s_214), .O(gate507inter3));
  inv1  gate2049(.a(s_215), .O(gate507inter4));
  nand2 gate2050(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate2051(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate2052(.a(G1276), .O(gate507inter7));
  inv1  gate2053(.a(G1277), .O(gate507inter8));
  nand2 gate2054(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate2055(.a(s_215), .b(gate507inter3), .O(gate507inter10));
  nor2  gate2056(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate2057(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate2058(.a(gate507inter12), .b(gate507inter1), .O(G1316));
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate1121(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate1122(.a(gate509inter0), .b(s_82), .O(gate509inter1));
  and2  gate1123(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate1124(.a(s_82), .O(gate509inter3));
  inv1  gate1125(.a(s_83), .O(gate509inter4));
  nand2 gate1126(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate1127(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate1128(.a(G1280), .O(gate509inter7));
  inv1  gate1129(.a(G1281), .O(gate509inter8));
  nand2 gate1130(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate1131(.a(s_83), .b(gate509inter3), .O(gate509inter10));
  nor2  gate1132(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate1133(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate1134(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate1205(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate1206(.a(gate514inter0), .b(s_94), .O(gate514inter1));
  and2  gate1207(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate1208(.a(s_94), .O(gate514inter3));
  inv1  gate1209(.a(s_95), .O(gate514inter4));
  nand2 gate1210(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate1211(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate1212(.a(G1290), .O(gate514inter7));
  inv1  gate1213(.a(G1291), .O(gate514inter8));
  nand2 gate1214(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate1215(.a(s_95), .b(gate514inter3), .O(gate514inter10));
  nor2  gate1216(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate1217(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate1218(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule