module c432 (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
             N430,N431,N432);
input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
      N99,N102,N105,N108,N112,N115;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141;
output N223,N329,N370,N421,N430,N431,N432;
wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12;


inv1 gate1( .a(N1), .O(N118) );
inv1 gate2( .a(N4), .O(N119) );
inv1 gate3( .a(N11), .O(N122) );
inv1 gate4( .a(N17), .O(N123) );
inv1 gate5( .a(N24), .O(N126) );
inv1 gate6( .a(N30), .O(N127) );
inv1 gate7( .a(N37), .O(N130) );
inv1 gate8( .a(N43), .O(N131) );
inv1 gate9( .a(N50), .O(N134) );
inv1 gate10( .a(N56), .O(N135) );
inv1 gate11( .a(N63), .O(N138) );
inv1 gate12( .a(N69), .O(N139) );
inv1 gate13( .a(N76), .O(N142) );
inv1 gate14( .a(N82), .O(N143) );
inv1 gate15( .a(N89), .O(N146) );
inv1 gate16( .a(N95), .O(N147) );
inv1 gate17( .a(N102), .O(N150) );
inv1 gate18( .a(N108), .O(N151) );
nand2 gate19( .a(N118), .b(N4), .O(N154) );

  xor2  gate945(.a(N119), .b(N8), .O(gate20inter0));
  nand2 gate946(.a(gate20inter0), .b(s_112), .O(gate20inter1));
  and2  gate947(.a(N119), .b(N8), .O(gate20inter2));
  inv1  gate948(.a(s_112), .O(gate20inter3));
  inv1  gate949(.a(s_113), .O(gate20inter4));
  nand2 gate950(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate951(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate952(.a(N8), .O(gate20inter7));
  inv1  gate953(.a(N119), .O(gate20inter8));
  nand2 gate954(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate955(.a(s_113), .b(gate20inter3), .O(gate20inter10));
  nor2  gate956(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate957(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate958(.a(gate20inter12), .b(gate20inter1), .O(N157));

  xor2  gate455(.a(N119), .b(N14), .O(gate21inter0));
  nand2 gate456(.a(gate21inter0), .b(s_42), .O(gate21inter1));
  and2  gate457(.a(N119), .b(N14), .O(gate21inter2));
  inv1  gate458(.a(s_42), .O(gate21inter3));
  inv1  gate459(.a(s_43), .O(gate21inter4));
  nand2 gate460(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate461(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate462(.a(N14), .O(gate21inter7));
  inv1  gate463(.a(N119), .O(gate21inter8));
  nand2 gate464(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate465(.a(s_43), .b(gate21inter3), .O(gate21inter10));
  nor2  gate466(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate467(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate468(.a(gate21inter12), .b(gate21inter1), .O(N158));

  xor2  gate651(.a(N17), .b(N122), .O(gate22inter0));
  nand2 gate652(.a(gate22inter0), .b(s_70), .O(gate22inter1));
  and2  gate653(.a(N17), .b(N122), .O(gate22inter2));
  inv1  gate654(.a(s_70), .O(gate22inter3));
  inv1  gate655(.a(s_71), .O(gate22inter4));
  nand2 gate656(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate657(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate658(.a(N122), .O(gate22inter7));
  inv1  gate659(.a(N17), .O(gate22inter8));
  nand2 gate660(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate661(.a(s_71), .b(gate22inter3), .O(gate22inter10));
  nor2  gate662(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate663(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate664(.a(gate22inter12), .b(gate22inter1), .O(N159));
nand2 gate23( .a(N126), .b(N30), .O(N162) );

  xor2  gate357(.a(N43), .b(N130), .O(gate24inter0));
  nand2 gate358(.a(gate24inter0), .b(s_28), .O(gate24inter1));
  and2  gate359(.a(N43), .b(N130), .O(gate24inter2));
  inv1  gate360(.a(s_28), .O(gate24inter3));
  inv1  gate361(.a(s_29), .O(gate24inter4));
  nand2 gate362(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate363(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate364(.a(N130), .O(gate24inter7));
  inv1  gate365(.a(N43), .O(gate24inter8));
  nand2 gate366(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate367(.a(s_29), .b(gate24inter3), .O(gate24inter10));
  nor2  gate368(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate369(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate370(.a(gate24inter12), .b(gate24inter1), .O(N165));
nand2 gate25( .a(N134), .b(N56), .O(N168) );

  xor2  gate553(.a(N69), .b(N138), .O(gate26inter0));
  nand2 gate554(.a(gate26inter0), .b(s_56), .O(gate26inter1));
  and2  gate555(.a(N69), .b(N138), .O(gate26inter2));
  inv1  gate556(.a(s_56), .O(gate26inter3));
  inv1  gate557(.a(s_57), .O(gate26inter4));
  nand2 gate558(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate559(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate560(.a(N138), .O(gate26inter7));
  inv1  gate561(.a(N69), .O(gate26inter8));
  nand2 gate562(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate563(.a(s_57), .b(gate26inter3), .O(gate26inter10));
  nor2  gate564(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate565(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate566(.a(gate26inter12), .b(gate26inter1), .O(N171));

  xor2  gate763(.a(N82), .b(N142), .O(gate27inter0));
  nand2 gate764(.a(gate27inter0), .b(s_86), .O(gate27inter1));
  and2  gate765(.a(N82), .b(N142), .O(gate27inter2));
  inv1  gate766(.a(s_86), .O(gate27inter3));
  inv1  gate767(.a(s_87), .O(gate27inter4));
  nand2 gate768(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate769(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate770(.a(N142), .O(gate27inter7));
  inv1  gate771(.a(N82), .O(gate27inter8));
  nand2 gate772(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate773(.a(s_87), .b(gate27inter3), .O(gate27inter10));
  nor2  gate774(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate775(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate776(.a(gate27inter12), .b(gate27inter1), .O(N174));

  xor2  gate1057(.a(N95), .b(N146), .O(gate28inter0));
  nand2 gate1058(.a(gate28inter0), .b(s_128), .O(gate28inter1));
  and2  gate1059(.a(N95), .b(N146), .O(gate28inter2));
  inv1  gate1060(.a(s_128), .O(gate28inter3));
  inv1  gate1061(.a(s_129), .O(gate28inter4));
  nand2 gate1062(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate1063(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate1064(.a(N146), .O(gate28inter7));
  inv1  gate1065(.a(N95), .O(gate28inter8));
  nand2 gate1066(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate1067(.a(s_129), .b(gate28inter3), .O(gate28inter10));
  nor2  gate1068(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate1069(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate1070(.a(gate28inter12), .b(gate28inter1), .O(N177));
nand2 gate29( .a(N150), .b(N108), .O(N180) );

  xor2  gate217(.a(N123), .b(N21), .O(gate30inter0));
  nand2 gate218(.a(gate30inter0), .b(s_8), .O(gate30inter1));
  and2  gate219(.a(N123), .b(N21), .O(gate30inter2));
  inv1  gate220(.a(s_8), .O(gate30inter3));
  inv1  gate221(.a(s_9), .O(gate30inter4));
  nand2 gate222(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate223(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate224(.a(N21), .O(gate30inter7));
  inv1  gate225(.a(N123), .O(gate30inter8));
  nand2 gate226(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate227(.a(s_9), .b(gate30inter3), .O(gate30inter10));
  nor2  gate228(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate229(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate230(.a(gate30inter12), .b(gate30inter1), .O(N183));

  xor2  gate889(.a(N123), .b(N27), .O(gate31inter0));
  nand2 gate890(.a(gate31inter0), .b(s_104), .O(gate31inter1));
  and2  gate891(.a(N123), .b(N27), .O(gate31inter2));
  inv1  gate892(.a(s_104), .O(gate31inter3));
  inv1  gate893(.a(s_105), .O(gate31inter4));
  nand2 gate894(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate895(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate896(.a(N27), .O(gate31inter7));
  inv1  gate897(.a(N123), .O(gate31inter8));
  nand2 gate898(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate899(.a(s_105), .b(gate31inter3), .O(gate31inter10));
  nor2  gate900(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate901(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate902(.a(gate31inter12), .b(gate31inter1), .O(N184));

  xor2  gate917(.a(N127), .b(N34), .O(gate32inter0));
  nand2 gate918(.a(gate32inter0), .b(s_108), .O(gate32inter1));
  and2  gate919(.a(N127), .b(N34), .O(gate32inter2));
  inv1  gate920(.a(s_108), .O(gate32inter3));
  inv1  gate921(.a(s_109), .O(gate32inter4));
  nand2 gate922(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate923(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate924(.a(N34), .O(gate32inter7));
  inv1  gate925(.a(N127), .O(gate32inter8));
  nand2 gate926(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate927(.a(s_109), .b(gate32inter3), .O(gate32inter10));
  nor2  gate928(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate929(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate930(.a(gate32inter12), .b(gate32inter1), .O(N185));
nor2 gate33( .a(N40), .b(N127), .O(N186) );

  xor2  gate1141(.a(N131), .b(N47), .O(gate34inter0));
  nand2 gate1142(.a(gate34inter0), .b(s_140), .O(gate34inter1));
  and2  gate1143(.a(N131), .b(N47), .O(gate34inter2));
  inv1  gate1144(.a(s_140), .O(gate34inter3));
  inv1  gate1145(.a(s_141), .O(gate34inter4));
  nand2 gate1146(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate1147(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate1148(.a(N47), .O(gate34inter7));
  inv1  gate1149(.a(N131), .O(gate34inter8));
  nand2 gate1150(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate1151(.a(s_141), .b(gate34inter3), .O(gate34inter10));
  nor2  gate1152(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate1153(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate1154(.a(gate34inter12), .b(gate34inter1), .O(N187));
nor2 gate35( .a(N53), .b(N131), .O(N188) );

  xor2  gate203(.a(N135), .b(N60), .O(gate36inter0));
  nand2 gate204(.a(gate36inter0), .b(s_6), .O(gate36inter1));
  and2  gate205(.a(N135), .b(N60), .O(gate36inter2));
  inv1  gate206(.a(s_6), .O(gate36inter3));
  inv1  gate207(.a(s_7), .O(gate36inter4));
  nand2 gate208(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate209(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate210(.a(N60), .O(gate36inter7));
  inv1  gate211(.a(N135), .O(gate36inter8));
  nand2 gate212(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate213(.a(s_7), .b(gate36inter3), .O(gate36inter10));
  nor2  gate214(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate215(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate216(.a(gate36inter12), .b(gate36inter1), .O(N189));

  xor2  gate973(.a(N135), .b(N66), .O(gate37inter0));
  nand2 gate974(.a(gate37inter0), .b(s_116), .O(gate37inter1));
  and2  gate975(.a(N135), .b(N66), .O(gate37inter2));
  inv1  gate976(.a(s_116), .O(gate37inter3));
  inv1  gate977(.a(s_117), .O(gate37inter4));
  nand2 gate978(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate979(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate980(.a(N66), .O(gate37inter7));
  inv1  gate981(.a(N135), .O(gate37inter8));
  nand2 gate982(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate983(.a(s_117), .b(gate37inter3), .O(gate37inter10));
  nor2  gate984(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate985(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate986(.a(gate37inter12), .b(gate37inter1), .O(N190));

  xor2  gate427(.a(N139), .b(N73), .O(gate38inter0));
  nand2 gate428(.a(gate38inter0), .b(s_38), .O(gate38inter1));
  and2  gate429(.a(N139), .b(N73), .O(gate38inter2));
  inv1  gate430(.a(s_38), .O(gate38inter3));
  inv1  gate431(.a(s_39), .O(gate38inter4));
  nand2 gate432(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate433(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate434(.a(N73), .O(gate38inter7));
  inv1  gate435(.a(N139), .O(gate38inter8));
  nand2 gate436(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate437(.a(s_39), .b(gate38inter3), .O(gate38inter10));
  nor2  gate438(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate439(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate440(.a(gate38inter12), .b(gate38inter1), .O(N191));
nor2 gate39( .a(N79), .b(N139), .O(N192) );

  xor2  gate315(.a(N143), .b(N86), .O(gate40inter0));
  nand2 gate316(.a(gate40inter0), .b(s_22), .O(gate40inter1));
  and2  gate317(.a(N143), .b(N86), .O(gate40inter2));
  inv1  gate318(.a(s_22), .O(gate40inter3));
  inv1  gate319(.a(s_23), .O(gate40inter4));
  nand2 gate320(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate321(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate322(.a(N86), .O(gate40inter7));
  inv1  gate323(.a(N143), .O(gate40inter8));
  nand2 gate324(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate325(.a(s_23), .b(gate40inter3), .O(gate40inter10));
  nor2  gate326(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate327(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate328(.a(gate40inter12), .b(gate40inter1), .O(N193));

  xor2  gate1015(.a(N143), .b(N92), .O(gate41inter0));
  nand2 gate1016(.a(gate41inter0), .b(s_122), .O(gate41inter1));
  and2  gate1017(.a(N143), .b(N92), .O(gate41inter2));
  inv1  gate1018(.a(s_122), .O(gate41inter3));
  inv1  gate1019(.a(s_123), .O(gate41inter4));
  nand2 gate1020(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate1021(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate1022(.a(N92), .O(gate41inter7));
  inv1  gate1023(.a(N143), .O(gate41inter8));
  nand2 gate1024(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate1025(.a(s_123), .b(gate41inter3), .O(gate41inter10));
  nor2  gate1026(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate1027(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate1028(.a(gate41inter12), .b(gate41inter1), .O(N194));

  xor2  gate1001(.a(N147), .b(N99), .O(gate42inter0));
  nand2 gate1002(.a(gate42inter0), .b(s_120), .O(gate42inter1));
  and2  gate1003(.a(N147), .b(N99), .O(gate42inter2));
  inv1  gate1004(.a(s_120), .O(gate42inter3));
  inv1  gate1005(.a(s_121), .O(gate42inter4));
  nand2 gate1006(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate1007(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate1008(.a(N99), .O(gate42inter7));
  inv1  gate1009(.a(N147), .O(gate42inter8));
  nand2 gate1010(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate1011(.a(s_121), .b(gate42inter3), .O(gate42inter10));
  nor2  gate1012(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate1013(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate1014(.a(gate42inter12), .b(gate42inter1), .O(N195));

  xor2  gate805(.a(N147), .b(N105), .O(gate43inter0));
  nand2 gate806(.a(gate43inter0), .b(s_92), .O(gate43inter1));
  and2  gate807(.a(N147), .b(N105), .O(gate43inter2));
  inv1  gate808(.a(s_92), .O(gate43inter3));
  inv1  gate809(.a(s_93), .O(gate43inter4));
  nand2 gate810(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate811(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate812(.a(N105), .O(gate43inter7));
  inv1  gate813(.a(N147), .O(gate43inter8));
  nand2 gate814(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate815(.a(s_93), .b(gate43inter3), .O(gate43inter10));
  nor2  gate816(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate817(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate818(.a(gate43inter12), .b(gate43inter1), .O(N196));

  xor2  gate1099(.a(N151), .b(N112), .O(gate44inter0));
  nand2 gate1100(.a(gate44inter0), .b(s_134), .O(gate44inter1));
  and2  gate1101(.a(N151), .b(N112), .O(gate44inter2));
  inv1  gate1102(.a(s_134), .O(gate44inter3));
  inv1  gate1103(.a(s_135), .O(gate44inter4));
  nand2 gate1104(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate1105(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate1106(.a(N112), .O(gate44inter7));
  inv1  gate1107(.a(N151), .O(gate44inter8));
  nand2 gate1108(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate1109(.a(s_135), .b(gate44inter3), .O(gate44inter10));
  nor2  gate1110(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate1111(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate1112(.a(gate44inter12), .b(gate44inter1), .O(N197));

  xor2  gate847(.a(N151), .b(N115), .O(gate45inter0));
  nand2 gate848(.a(gate45inter0), .b(s_98), .O(gate45inter1));
  and2  gate849(.a(N151), .b(N115), .O(gate45inter2));
  inv1  gate850(.a(s_98), .O(gate45inter3));
  inv1  gate851(.a(s_99), .O(gate45inter4));
  nand2 gate852(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate853(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate854(.a(N115), .O(gate45inter7));
  inv1  gate855(.a(N151), .O(gate45inter8));
  nand2 gate856(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate857(.a(s_99), .b(gate45inter3), .O(gate45inter10));
  nor2  gate858(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate859(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate860(.a(gate45inter12), .b(gate45inter1), .O(N198));
and9 gate46( .a(N154), .b(N159), .c(N162), .d(N165), .e(N168), .f(N171), .g(N174), .h(N177), .i(N180), .O(N199) );
inv1 gate47( .a(N199), .O(N203) );
inv1 gate48( .a(N199), .O(N213) );
inv1 gate49( .a(N199), .O(N223) );

  xor2  gate581(.a(N154), .b(N203), .O(gate50inter0));
  nand2 gate582(.a(gate50inter0), .b(s_60), .O(gate50inter1));
  and2  gate583(.a(N154), .b(N203), .O(gate50inter2));
  inv1  gate584(.a(s_60), .O(gate50inter3));
  inv1  gate585(.a(s_61), .O(gate50inter4));
  nand2 gate586(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate587(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate588(.a(N203), .O(gate50inter7));
  inv1  gate589(.a(N154), .O(gate50inter8));
  nand2 gate590(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate591(.a(s_61), .b(gate50inter3), .O(gate50inter10));
  nor2  gate592(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate593(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate594(.a(gate50inter12), .b(gate50inter1), .O(N224));

  xor2  gate385(.a(N159), .b(N203), .O(gate51inter0));
  nand2 gate386(.a(gate51inter0), .b(s_32), .O(gate51inter1));
  and2  gate387(.a(N159), .b(N203), .O(gate51inter2));
  inv1  gate388(.a(s_32), .O(gate51inter3));
  inv1  gate389(.a(s_33), .O(gate51inter4));
  nand2 gate390(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate391(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate392(.a(N203), .O(gate51inter7));
  inv1  gate393(.a(N159), .O(gate51inter8));
  nand2 gate394(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate395(.a(s_33), .b(gate51inter3), .O(gate51inter10));
  nor2  gate396(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate397(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate398(.a(gate51inter12), .b(gate51inter1), .O(N227));

  xor2  gate371(.a(N162), .b(N203), .O(gate52inter0));
  nand2 gate372(.a(gate52inter0), .b(s_30), .O(gate52inter1));
  and2  gate373(.a(N162), .b(N203), .O(gate52inter2));
  inv1  gate374(.a(s_30), .O(gate52inter3));
  inv1  gate375(.a(s_31), .O(gate52inter4));
  nand2 gate376(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate377(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate378(.a(N203), .O(gate52inter7));
  inv1  gate379(.a(N162), .O(gate52inter8));
  nand2 gate380(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate381(.a(s_31), .b(gate52inter3), .O(gate52inter10));
  nor2  gate382(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate383(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate384(.a(gate52inter12), .b(gate52inter1), .O(N230));
xor2 gate53( .a(N203), .b(N165), .O(N233) );

  xor2  gate735(.a(N168), .b(N203), .O(gate54inter0));
  nand2 gate736(.a(gate54inter0), .b(s_82), .O(gate54inter1));
  and2  gate737(.a(N168), .b(N203), .O(gate54inter2));
  inv1  gate738(.a(s_82), .O(gate54inter3));
  inv1  gate739(.a(s_83), .O(gate54inter4));
  nand2 gate740(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate741(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate742(.a(N203), .O(gate54inter7));
  inv1  gate743(.a(N168), .O(gate54inter8));
  nand2 gate744(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate745(.a(s_83), .b(gate54inter3), .O(gate54inter10));
  nor2  gate746(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate747(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate748(.a(gate54inter12), .b(gate54inter1), .O(N236));

  xor2  gate721(.a(N171), .b(N203), .O(gate55inter0));
  nand2 gate722(.a(gate55inter0), .b(s_80), .O(gate55inter1));
  and2  gate723(.a(N171), .b(N203), .O(gate55inter2));
  inv1  gate724(.a(s_80), .O(gate55inter3));
  inv1  gate725(.a(s_81), .O(gate55inter4));
  nand2 gate726(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate727(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate728(.a(N203), .O(gate55inter7));
  inv1  gate729(.a(N171), .O(gate55inter8));
  nand2 gate730(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate731(.a(s_81), .b(gate55inter3), .O(gate55inter10));
  nor2  gate732(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate733(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate734(.a(gate55inter12), .b(gate55inter1), .O(N239));

  xor2  gate441(.a(N213), .b(N1), .O(gate56inter0));
  nand2 gate442(.a(gate56inter0), .b(s_40), .O(gate56inter1));
  and2  gate443(.a(N213), .b(N1), .O(gate56inter2));
  inv1  gate444(.a(s_40), .O(gate56inter3));
  inv1  gate445(.a(s_41), .O(gate56inter4));
  nand2 gate446(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate447(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate448(.a(N1), .O(gate56inter7));
  inv1  gate449(.a(N213), .O(gate56inter8));
  nand2 gate450(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate451(.a(s_41), .b(gate56inter3), .O(gate56inter10));
  nor2  gate452(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate453(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate454(.a(gate56inter12), .b(gate56inter1), .O(N242));
xor2 gate57( .a(N203), .b(N174), .O(N243) );

  xor2  gate595(.a(N11), .b(N213), .O(gate58inter0));
  nand2 gate596(.a(gate58inter0), .b(s_62), .O(gate58inter1));
  and2  gate597(.a(N11), .b(N213), .O(gate58inter2));
  inv1  gate598(.a(s_62), .O(gate58inter3));
  inv1  gate599(.a(s_63), .O(gate58inter4));
  nand2 gate600(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate601(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate602(.a(N213), .O(gate58inter7));
  inv1  gate603(.a(N11), .O(gate58inter8));
  nand2 gate604(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate605(.a(s_63), .b(gate58inter3), .O(gate58inter10));
  nor2  gate606(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate607(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate608(.a(gate58inter12), .b(gate58inter1), .O(N246));

  xor2  gate707(.a(N177), .b(N203), .O(gate59inter0));
  nand2 gate708(.a(gate59inter0), .b(s_78), .O(gate59inter1));
  and2  gate709(.a(N177), .b(N203), .O(gate59inter2));
  inv1  gate710(.a(s_78), .O(gate59inter3));
  inv1  gate711(.a(s_79), .O(gate59inter4));
  nand2 gate712(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate713(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate714(.a(N203), .O(gate59inter7));
  inv1  gate715(.a(N177), .O(gate59inter8));
  nand2 gate716(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate717(.a(s_79), .b(gate59inter3), .O(gate59inter10));
  nor2  gate718(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate719(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate720(.a(gate59inter12), .b(gate59inter1), .O(N247));
nand2 gate60( .a(N213), .b(N24), .O(N250) );
xor2 gate61( .a(N203), .b(N180), .O(N251) );

  xor2  gate231(.a(N37), .b(N213), .O(gate62inter0));
  nand2 gate232(.a(gate62inter0), .b(s_10), .O(gate62inter1));
  and2  gate233(.a(N37), .b(N213), .O(gate62inter2));
  inv1  gate234(.a(s_10), .O(gate62inter3));
  inv1  gate235(.a(s_11), .O(gate62inter4));
  nand2 gate236(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate237(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate238(.a(N213), .O(gate62inter7));
  inv1  gate239(.a(N37), .O(gate62inter8));
  nand2 gate240(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate241(.a(s_11), .b(gate62inter3), .O(gate62inter10));
  nor2  gate242(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate243(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate244(.a(gate62inter12), .b(gate62inter1), .O(N254));

  xor2  gate749(.a(N50), .b(N213), .O(gate63inter0));
  nand2 gate750(.a(gate63inter0), .b(s_84), .O(gate63inter1));
  and2  gate751(.a(N50), .b(N213), .O(gate63inter2));
  inv1  gate752(.a(s_84), .O(gate63inter3));
  inv1  gate753(.a(s_85), .O(gate63inter4));
  nand2 gate754(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate755(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate756(.a(N213), .O(gate63inter7));
  inv1  gate757(.a(N50), .O(gate63inter8));
  nand2 gate758(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate759(.a(s_85), .b(gate63inter3), .O(gate63inter10));
  nor2  gate760(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate761(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate762(.a(gate63inter12), .b(gate63inter1), .O(N255));

  xor2  gate679(.a(N63), .b(N213), .O(gate64inter0));
  nand2 gate680(.a(gate64inter0), .b(s_74), .O(gate64inter1));
  and2  gate681(.a(N63), .b(N213), .O(gate64inter2));
  inv1  gate682(.a(s_74), .O(gate64inter3));
  inv1  gate683(.a(s_75), .O(gate64inter4));
  nand2 gate684(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate685(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate686(.a(N213), .O(gate64inter7));
  inv1  gate687(.a(N63), .O(gate64inter8));
  nand2 gate688(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate689(.a(s_75), .b(gate64inter3), .O(gate64inter10));
  nor2  gate690(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate691(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate692(.a(gate64inter12), .b(gate64inter1), .O(N256));

  xor2  gate539(.a(N76), .b(N213), .O(gate65inter0));
  nand2 gate540(.a(gate65inter0), .b(s_54), .O(gate65inter1));
  and2  gate541(.a(N76), .b(N213), .O(gate65inter2));
  inv1  gate542(.a(s_54), .O(gate65inter3));
  inv1  gate543(.a(s_55), .O(gate65inter4));
  nand2 gate544(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate545(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate546(.a(N213), .O(gate65inter7));
  inv1  gate547(.a(N76), .O(gate65inter8));
  nand2 gate548(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate549(.a(s_55), .b(gate65inter3), .O(gate65inter10));
  nor2  gate550(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate551(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate552(.a(gate65inter12), .b(gate65inter1), .O(N257));

  xor2  gate903(.a(N89), .b(N213), .O(gate66inter0));
  nand2 gate904(.a(gate66inter0), .b(s_106), .O(gate66inter1));
  and2  gate905(.a(N89), .b(N213), .O(gate66inter2));
  inv1  gate906(.a(s_106), .O(gate66inter3));
  inv1  gate907(.a(s_107), .O(gate66inter4));
  nand2 gate908(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate909(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate910(.a(N213), .O(gate66inter7));
  inv1  gate911(.a(N89), .O(gate66inter8));
  nand2 gate912(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate913(.a(s_107), .b(gate66inter3), .O(gate66inter10));
  nor2  gate914(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate915(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate916(.a(gate66inter12), .b(gate66inter1), .O(N258));
nand2 gate67( .a(N213), .b(N102), .O(N259) );

  xor2  gate259(.a(N157), .b(N224), .O(gate68inter0));
  nand2 gate260(.a(gate68inter0), .b(s_14), .O(gate68inter1));
  and2  gate261(.a(N157), .b(N224), .O(gate68inter2));
  inv1  gate262(.a(s_14), .O(gate68inter3));
  inv1  gate263(.a(s_15), .O(gate68inter4));
  nand2 gate264(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate265(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate266(.a(N224), .O(gate68inter7));
  inv1  gate267(.a(N157), .O(gate68inter8));
  nand2 gate268(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate269(.a(s_15), .b(gate68inter3), .O(gate68inter10));
  nor2  gate270(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate271(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate272(.a(gate68inter12), .b(gate68inter1), .O(N260));

  xor2  gate623(.a(N158), .b(N224), .O(gate69inter0));
  nand2 gate624(.a(gate69inter0), .b(s_66), .O(gate69inter1));
  and2  gate625(.a(N158), .b(N224), .O(gate69inter2));
  inv1  gate626(.a(s_66), .O(gate69inter3));
  inv1  gate627(.a(s_67), .O(gate69inter4));
  nand2 gate628(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate629(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate630(.a(N224), .O(gate69inter7));
  inv1  gate631(.a(N158), .O(gate69inter8));
  nand2 gate632(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate633(.a(s_67), .b(gate69inter3), .O(gate69inter10));
  nor2  gate634(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate635(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate636(.a(gate69inter12), .b(gate69inter1), .O(N263));

  xor2  gate287(.a(N183), .b(N227), .O(gate70inter0));
  nand2 gate288(.a(gate70inter0), .b(s_18), .O(gate70inter1));
  and2  gate289(.a(N183), .b(N227), .O(gate70inter2));
  inv1  gate290(.a(s_18), .O(gate70inter3));
  inv1  gate291(.a(s_19), .O(gate70inter4));
  nand2 gate292(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate293(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate294(.a(N227), .O(gate70inter7));
  inv1  gate295(.a(N183), .O(gate70inter8));
  nand2 gate296(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate297(.a(s_19), .b(gate70inter3), .O(gate70inter10));
  nor2  gate298(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate299(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate300(.a(gate70inter12), .b(gate70inter1), .O(N264));
nand2 gate71( .a(N230), .b(N185), .O(N267) );

  xor2  gate861(.a(N187), .b(N233), .O(gate72inter0));
  nand2 gate862(.a(gate72inter0), .b(s_100), .O(gate72inter1));
  and2  gate863(.a(N187), .b(N233), .O(gate72inter2));
  inv1  gate864(.a(s_100), .O(gate72inter3));
  inv1  gate865(.a(s_101), .O(gate72inter4));
  nand2 gate866(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate867(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate868(.a(N233), .O(gate72inter7));
  inv1  gate869(.a(N187), .O(gate72inter8));
  nand2 gate870(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate871(.a(s_101), .b(gate72inter3), .O(gate72inter10));
  nor2  gate872(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate873(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate874(.a(gate72inter12), .b(gate72inter1), .O(N270));

  xor2  gate987(.a(N189), .b(N236), .O(gate73inter0));
  nand2 gate988(.a(gate73inter0), .b(s_118), .O(gate73inter1));
  and2  gate989(.a(N189), .b(N236), .O(gate73inter2));
  inv1  gate990(.a(s_118), .O(gate73inter3));
  inv1  gate991(.a(s_119), .O(gate73inter4));
  nand2 gate992(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate993(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate994(.a(N236), .O(gate73inter7));
  inv1  gate995(.a(N189), .O(gate73inter8));
  nand2 gate996(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate997(.a(s_119), .b(gate73inter3), .O(gate73inter10));
  nor2  gate998(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate999(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate1000(.a(gate73inter12), .b(gate73inter1), .O(N273));
nand2 gate74( .a(N239), .b(N191), .O(N276) );

  xor2  gate609(.a(N193), .b(N243), .O(gate75inter0));
  nand2 gate610(.a(gate75inter0), .b(s_64), .O(gate75inter1));
  and2  gate611(.a(N193), .b(N243), .O(gate75inter2));
  inv1  gate612(.a(s_64), .O(gate75inter3));
  inv1  gate613(.a(s_65), .O(gate75inter4));
  nand2 gate614(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate615(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate616(.a(N243), .O(gate75inter7));
  inv1  gate617(.a(N193), .O(gate75inter8));
  nand2 gate618(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate619(.a(s_65), .b(gate75inter3), .O(gate75inter10));
  nor2  gate620(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate621(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate622(.a(gate75inter12), .b(gate75inter1), .O(N279));
nand2 gate76( .a(N247), .b(N195), .O(N282) );
nand2 gate77( .a(N251), .b(N197), .O(N285) );

  xor2  gate567(.a(N184), .b(N227), .O(gate78inter0));
  nand2 gate568(.a(gate78inter0), .b(s_58), .O(gate78inter1));
  and2  gate569(.a(N184), .b(N227), .O(gate78inter2));
  inv1  gate570(.a(s_58), .O(gate78inter3));
  inv1  gate571(.a(s_59), .O(gate78inter4));
  nand2 gate572(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate573(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate574(.a(N227), .O(gate78inter7));
  inv1  gate575(.a(N184), .O(gate78inter8));
  nand2 gate576(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate577(.a(s_59), .b(gate78inter3), .O(gate78inter10));
  nor2  gate578(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate579(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate580(.a(gate78inter12), .b(gate78inter1), .O(N288));
nand2 gate79( .a(N230), .b(N186), .O(N289) );

  xor2  gate469(.a(N188), .b(N233), .O(gate80inter0));
  nand2 gate470(.a(gate80inter0), .b(s_44), .O(gate80inter1));
  and2  gate471(.a(N188), .b(N233), .O(gate80inter2));
  inv1  gate472(.a(s_44), .O(gate80inter3));
  inv1  gate473(.a(s_45), .O(gate80inter4));
  nand2 gate474(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate475(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate476(.a(N233), .O(gate80inter7));
  inv1  gate477(.a(N188), .O(gate80inter8));
  nand2 gate478(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate479(.a(s_45), .b(gate80inter3), .O(gate80inter10));
  nor2  gate480(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate481(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate482(.a(gate80inter12), .b(gate80inter1), .O(N290));
nand2 gate81( .a(N236), .b(N190), .O(N291) );

  xor2  gate497(.a(N192), .b(N239), .O(gate82inter0));
  nand2 gate498(.a(gate82inter0), .b(s_48), .O(gate82inter1));
  and2  gate499(.a(N192), .b(N239), .O(gate82inter2));
  inv1  gate500(.a(s_48), .O(gate82inter3));
  inv1  gate501(.a(s_49), .O(gate82inter4));
  nand2 gate502(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate503(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate504(.a(N239), .O(gate82inter7));
  inv1  gate505(.a(N192), .O(gate82inter8));
  nand2 gate506(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate507(.a(s_49), .b(gate82inter3), .O(gate82inter10));
  nor2  gate508(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate509(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate510(.a(gate82inter12), .b(gate82inter1), .O(N292));

  xor2  gate399(.a(N194), .b(N243), .O(gate83inter0));
  nand2 gate400(.a(gate83inter0), .b(s_34), .O(gate83inter1));
  and2  gate401(.a(N194), .b(N243), .O(gate83inter2));
  inv1  gate402(.a(s_34), .O(gate83inter3));
  inv1  gate403(.a(s_35), .O(gate83inter4));
  nand2 gate404(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate405(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate406(.a(N243), .O(gate83inter7));
  inv1  gate407(.a(N194), .O(gate83inter8));
  nand2 gate408(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate409(.a(s_35), .b(gate83inter3), .O(gate83inter10));
  nor2  gate410(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate411(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate412(.a(gate83inter12), .b(gate83inter1), .O(N293));

  xor2  gate483(.a(N196), .b(N247), .O(gate84inter0));
  nand2 gate484(.a(gate84inter0), .b(s_46), .O(gate84inter1));
  and2  gate485(.a(N196), .b(N247), .O(gate84inter2));
  inv1  gate486(.a(s_46), .O(gate84inter3));
  inv1  gate487(.a(s_47), .O(gate84inter4));
  nand2 gate488(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate489(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate490(.a(N247), .O(gate84inter7));
  inv1  gate491(.a(N196), .O(gate84inter8));
  nand2 gate492(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate493(.a(s_47), .b(gate84inter3), .O(gate84inter10));
  nor2  gate494(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate495(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate496(.a(gate84inter12), .b(gate84inter1), .O(N294));

  xor2  gate343(.a(N198), .b(N251), .O(gate85inter0));
  nand2 gate344(.a(gate85inter0), .b(s_26), .O(gate85inter1));
  and2  gate345(.a(N198), .b(N251), .O(gate85inter2));
  inv1  gate346(.a(s_26), .O(gate85inter3));
  inv1  gate347(.a(s_27), .O(gate85inter4));
  nand2 gate348(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate349(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate350(.a(N251), .O(gate85inter7));
  inv1  gate351(.a(N198), .O(gate85inter8));
  nand2 gate352(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate353(.a(s_27), .b(gate85inter3), .O(gate85inter10));
  nor2  gate354(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate355(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate356(.a(gate85inter12), .b(gate85inter1), .O(N295));
and9 gate86( .a(N260), .b(N264), .c(N267), .d(N270), .e(N273), .f(N276), .g(N279), .h(N282), .i(N285), .O(N296) );
inv1 gate87( .a(N263), .O(N300) );
inv1 gate88( .a(N288), .O(N301) );
inv1 gate89( .a(N289), .O(N302) );
inv1 gate90( .a(N290), .O(N303) );
inv1 gate91( .a(N291), .O(N304) );
inv1 gate92( .a(N292), .O(N305) );
inv1 gate93( .a(N293), .O(N306) );
inv1 gate94( .a(N294), .O(N307) );
inv1 gate95( .a(N295), .O(N308) );
inv1 gate96( .a(N296), .O(N309) );
inv1 gate97( .a(N296), .O(N319) );
inv1 gate98( .a(N296), .O(N329) );

  xor2  gate931(.a(N260), .b(N309), .O(gate99inter0));
  nand2 gate932(.a(gate99inter0), .b(s_110), .O(gate99inter1));
  and2  gate933(.a(N260), .b(N309), .O(gate99inter2));
  inv1  gate934(.a(s_110), .O(gate99inter3));
  inv1  gate935(.a(s_111), .O(gate99inter4));
  nand2 gate936(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate937(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate938(.a(N309), .O(gate99inter7));
  inv1  gate939(.a(N260), .O(gate99inter8));
  nand2 gate940(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate941(.a(s_111), .b(gate99inter3), .O(gate99inter10));
  nor2  gate942(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate943(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate944(.a(gate99inter12), .b(gate99inter1), .O(N330));

  xor2  gate1113(.a(N264), .b(N309), .O(gate100inter0));
  nand2 gate1114(.a(gate100inter0), .b(s_136), .O(gate100inter1));
  and2  gate1115(.a(N264), .b(N309), .O(gate100inter2));
  inv1  gate1116(.a(s_136), .O(gate100inter3));
  inv1  gate1117(.a(s_137), .O(gate100inter4));
  nand2 gate1118(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate1119(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate1120(.a(N309), .O(gate100inter7));
  inv1  gate1121(.a(N264), .O(gate100inter8));
  nand2 gate1122(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate1123(.a(s_137), .b(gate100inter3), .O(gate100inter10));
  nor2  gate1124(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate1125(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate1126(.a(gate100inter12), .b(gate100inter1), .O(N331));

  xor2  gate1029(.a(N267), .b(N309), .O(gate101inter0));
  nand2 gate1030(.a(gate101inter0), .b(s_124), .O(gate101inter1));
  and2  gate1031(.a(N267), .b(N309), .O(gate101inter2));
  inv1  gate1032(.a(s_124), .O(gate101inter3));
  inv1  gate1033(.a(s_125), .O(gate101inter4));
  nand2 gate1034(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate1035(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate1036(.a(N309), .O(gate101inter7));
  inv1  gate1037(.a(N267), .O(gate101inter8));
  nand2 gate1038(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate1039(.a(s_125), .b(gate101inter3), .O(gate101inter10));
  nor2  gate1040(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate1041(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate1042(.a(gate101inter12), .b(gate101inter1), .O(N332));

  xor2  gate875(.a(N270), .b(N309), .O(gate102inter0));
  nand2 gate876(.a(gate102inter0), .b(s_102), .O(gate102inter1));
  and2  gate877(.a(N270), .b(N309), .O(gate102inter2));
  inv1  gate878(.a(s_102), .O(gate102inter3));
  inv1  gate879(.a(s_103), .O(gate102inter4));
  nand2 gate880(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate881(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate882(.a(N309), .O(gate102inter7));
  inv1  gate883(.a(N270), .O(gate102inter8));
  nand2 gate884(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate885(.a(s_103), .b(gate102inter3), .O(gate102inter10));
  nor2  gate886(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate887(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate888(.a(gate102inter12), .b(gate102inter1), .O(N333));

  xor2  gate161(.a(N319), .b(N8), .O(gate103inter0));
  nand2 gate162(.a(gate103inter0), .b(s_0), .O(gate103inter1));
  and2  gate163(.a(N319), .b(N8), .O(gate103inter2));
  inv1  gate164(.a(s_0), .O(gate103inter3));
  inv1  gate165(.a(s_1), .O(gate103inter4));
  nand2 gate166(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate167(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate168(.a(N8), .O(gate103inter7));
  inv1  gate169(.a(N319), .O(gate103inter8));
  nand2 gate170(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate171(.a(s_1), .b(gate103inter3), .O(gate103inter10));
  nor2  gate172(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate173(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate174(.a(gate103inter12), .b(gate103inter1), .O(N334));

  xor2  gate693(.a(N273), .b(N309), .O(gate104inter0));
  nand2 gate694(.a(gate104inter0), .b(s_76), .O(gate104inter1));
  and2  gate695(.a(N273), .b(N309), .O(gate104inter2));
  inv1  gate696(.a(s_76), .O(gate104inter3));
  inv1  gate697(.a(s_77), .O(gate104inter4));
  nand2 gate698(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate699(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate700(.a(N309), .O(gate104inter7));
  inv1  gate701(.a(N273), .O(gate104inter8));
  nand2 gate702(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate703(.a(s_77), .b(gate104inter3), .O(gate104inter10));
  nor2  gate704(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate705(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate706(.a(gate104inter12), .b(gate104inter1), .O(N335));
nand2 gate105( .a(N319), .b(N21), .O(N336) );

  xor2  gate637(.a(N276), .b(N309), .O(gate106inter0));
  nand2 gate638(.a(gate106inter0), .b(s_68), .O(gate106inter1));
  and2  gate639(.a(N276), .b(N309), .O(gate106inter2));
  inv1  gate640(.a(s_68), .O(gate106inter3));
  inv1  gate641(.a(s_69), .O(gate106inter4));
  nand2 gate642(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate643(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate644(.a(N309), .O(gate106inter7));
  inv1  gate645(.a(N276), .O(gate106inter8));
  nand2 gate646(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate647(.a(s_69), .b(gate106inter3), .O(gate106inter10));
  nor2  gate648(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate649(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate650(.a(gate106inter12), .b(gate106inter1), .O(N337));

  xor2  gate1085(.a(N34), .b(N319), .O(gate107inter0));
  nand2 gate1086(.a(gate107inter0), .b(s_132), .O(gate107inter1));
  and2  gate1087(.a(N34), .b(N319), .O(gate107inter2));
  inv1  gate1088(.a(s_132), .O(gate107inter3));
  inv1  gate1089(.a(s_133), .O(gate107inter4));
  nand2 gate1090(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate1091(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate1092(.a(N319), .O(gate107inter7));
  inv1  gate1093(.a(N34), .O(gate107inter8));
  nand2 gate1094(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate1095(.a(s_133), .b(gate107inter3), .O(gate107inter10));
  nor2  gate1096(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate1097(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate1098(.a(gate107inter12), .b(gate107inter1), .O(N338));
xor2 gate108( .a(N309), .b(N279), .O(N339) );
nand2 gate109( .a(N319), .b(N47), .O(N340) );

  xor2  gate1043(.a(N282), .b(N309), .O(gate110inter0));
  nand2 gate1044(.a(gate110inter0), .b(s_126), .O(gate110inter1));
  and2  gate1045(.a(N282), .b(N309), .O(gate110inter2));
  inv1  gate1046(.a(s_126), .O(gate110inter3));
  inv1  gate1047(.a(s_127), .O(gate110inter4));
  nand2 gate1048(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1049(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1050(.a(N309), .O(gate110inter7));
  inv1  gate1051(.a(N282), .O(gate110inter8));
  nand2 gate1052(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1053(.a(s_127), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1054(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1055(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1056(.a(gate110inter12), .b(gate110inter1), .O(N341));

  xor2  gate189(.a(N60), .b(N319), .O(gate111inter0));
  nand2 gate190(.a(gate111inter0), .b(s_4), .O(gate111inter1));
  and2  gate191(.a(N60), .b(N319), .O(gate111inter2));
  inv1  gate192(.a(s_4), .O(gate111inter3));
  inv1  gate193(.a(s_5), .O(gate111inter4));
  nand2 gate194(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate195(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate196(.a(N319), .O(gate111inter7));
  inv1  gate197(.a(N60), .O(gate111inter8));
  nand2 gate198(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate199(.a(s_5), .b(gate111inter3), .O(gate111inter10));
  nor2  gate200(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate201(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate202(.a(gate111inter12), .b(gate111inter1), .O(N342));

  xor2  gate959(.a(N285), .b(N309), .O(gate112inter0));
  nand2 gate960(.a(gate112inter0), .b(s_114), .O(gate112inter1));
  and2  gate961(.a(N285), .b(N309), .O(gate112inter2));
  inv1  gate962(.a(s_114), .O(gate112inter3));
  inv1  gate963(.a(s_115), .O(gate112inter4));
  nand2 gate964(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate965(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate966(.a(N309), .O(gate112inter7));
  inv1  gate967(.a(N285), .O(gate112inter8));
  nand2 gate968(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate969(.a(s_115), .b(gate112inter3), .O(gate112inter10));
  nor2  gate970(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate971(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate972(.a(gate112inter12), .b(gate112inter1), .O(N343));

  xor2  gate511(.a(N73), .b(N319), .O(gate113inter0));
  nand2 gate512(.a(gate113inter0), .b(s_50), .O(gate113inter1));
  and2  gate513(.a(N73), .b(N319), .O(gate113inter2));
  inv1  gate514(.a(s_50), .O(gate113inter3));
  inv1  gate515(.a(s_51), .O(gate113inter4));
  nand2 gate516(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate517(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate518(.a(N319), .O(gate113inter7));
  inv1  gate519(.a(N73), .O(gate113inter8));
  nand2 gate520(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate521(.a(s_51), .b(gate113inter3), .O(gate113inter10));
  nor2  gate522(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate523(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate524(.a(gate113inter12), .b(gate113inter1), .O(N344));
nand2 gate114( .a(N319), .b(N86), .O(N345) );

  xor2  gate819(.a(N99), .b(N319), .O(gate115inter0));
  nand2 gate820(.a(gate115inter0), .b(s_94), .O(gate115inter1));
  and2  gate821(.a(N99), .b(N319), .O(gate115inter2));
  inv1  gate822(.a(s_94), .O(gate115inter3));
  inv1  gate823(.a(s_95), .O(gate115inter4));
  nand2 gate824(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate825(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate826(.a(N319), .O(gate115inter7));
  inv1  gate827(.a(N99), .O(gate115inter8));
  nand2 gate828(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate829(.a(s_95), .b(gate115inter3), .O(gate115inter10));
  nor2  gate830(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate831(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate832(.a(gate115inter12), .b(gate115inter1), .O(N346));

  xor2  gate833(.a(N112), .b(N319), .O(gate116inter0));
  nand2 gate834(.a(gate116inter0), .b(s_96), .O(gate116inter1));
  and2  gate835(.a(N112), .b(N319), .O(gate116inter2));
  inv1  gate836(.a(s_96), .O(gate116inter3));
  inv1  gate837(.a(s_97), .O(gate116inter4));
  nand2 gate838(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate839(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate840(.a(N319), .O(gate116inter7));
  inv1  gate841(.a(N112), .O(gate116inter8));
  nand2 gate842(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate843(.a(s_97), .b(gate116inter3), .O(gate116inter10));
  nor2  gate844(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate845(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate846(.a(gate116inter12), .b(gate116inter1), .O(N347));

  xor2  gate791(.a(N300), .b(N330), .O(gate117inter0));
  nand2 gate792(.a(gate117inter0), .b(s_90), .O(gate117inter1));
  and2  gate793(.a(N300), .b(N330), .O(gate117inter2));
  inv1  gate794(.a(s_90), .O(gate117inter3));
  inv1  gate795(.a(s_91), .O(gate117inter4));
  nand2 gate796(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate797(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate798(.a(N330), .O(gate117inter7));
  inv1  gate799(.a(N300), .O(gate117inter8));
  nand2 gate800(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate801(.a(s_91), .b(gate117inter3), .O(gate117inter10));
  nor2  gate802(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate803(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate804(.a(gate117inter12), .b(gate117inter1), .O(N348));

  xor2  gate1127(.a(N301), .b(N331), .O(gate118inter0));
  nand2 gate1128(.a(gate118inter0), .b(s_138), .O(gate118inter1));
  and2  gate1129(.a(N301), .b(N331), .O(gate118inter2));
  inv1  gate1130(.a(s_138), .O(gate118inter3));
  inv1  gate1131(.a(s_139), .O(gate118inter4));
  nand2 gate1132(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate1133(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate1134(.a(N331), .O(gate118inter7));
  inv1  gate1135(.a(N301), .O(gate118inter8));
  nand2 gate1136(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate1137(.a(s_139), .b(gate118inter3), .O(gate118inter10));
  nor2  gate1138(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate1139(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate1140(.a(gate118inter12), .b(gate118inter1), .O(N349));

  xor2  gate777(.a(N302), .b(N332), .O(gate119inter0));
  nand2 gate778(.a(gate119inter0), .b(s_88), .O(gate119inter1));
  and2  gate779(.a(N302), .b(N332), .O(gate119inter2));
  inv1  gate780(.a(s_88), .O(gate119inter3));
  inv1  gate781(.a(s_89), .O(gate119inter4));
  nand2 gate782(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate783(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate784(.a(N332), .O(gate119inter7));
  inv1  gate785(.a(N302), .O(gate119inter8));
  nand2 gate786(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate787(.a(s_89), .b(gate119inter3), .O(gate119inter10));
  nor2  gate788(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate789(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate790(.a(gate119inter12), .b(gate119inter1), .O(N350));

  xor2  gate665(.a(N303), .b(N333), .O(gate120inter0));
  nand2 gate666(.a(gate120inter0), .b(s_72), .O(gate120inter1));
  and2  gate667(.a(N303), .b(N333), .O(gate120inter2));
  inv1  gate668(.a(s_72), .O(gate120inter3));
  inv1  gate669(.a(s_73), .O(gate120inter4));
  nand2 gate670(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate671(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate672(.a(N333), .O(gate120inter7));
  inv1  gate673(.a(N303), .O(gate120inter8));
  nand2 gate674(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate675(.a(s_73), .b(gate120inter3), .O(gate120inter10));
  nor2  gate676(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate677(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate678(.a(gate120inter12), .b(gate120inter1), .O(N351));
nand2 gate121( .a(N335), .b(N304), .O(N352) );
nand2 gate122( .a(N337), .b(N305), .O(N353) );
nand2 gate123( .a(N339), .b(N306), .O(N354) );
nand2 gate124( .a(N341), .b(N307), .O(N355) );

  xor2  gate329(.a(N308), .b(N343), .O(gate125inter0));
  nand2 gate330(.a(gate125inter0), .b(s_24), .O(gate125inter1));
  and2  gate331(.a(N308), .b(N343), .O(gate125inter2));
  inv1  gate332(.a(s_24), .O(gate125inter3));
  inv1  gate333(.a(s_25), .O(gate125inter4));
  nand2 gate334(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate335(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate336(.a(N343), .O(gate125inter7));
  inv1  gate337(.a(N308), .O(gate125inter8));
  nand2 gate338(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate339(.a(s_25), .b(gate125inter3), .O(gate125inter10));
  nor2  gate340(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate341(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate342(.a(gate125inter12), .b(gate125inter1), .O(N356));
and9 gate126( .a(N348), .b(N349), .c(N350), .d(N351), .e(N352), .f(N353), .g(N354), .h(N355), .i(N356), .O(N357) );
inv1 gate127( .a(N357), .O(N360) );
inv1 gate128( .a(N357), .O(N370) );

  xor2  gate301(.a(N360), .b(N14), .O(gate129inter0));
  nand2 gate302(.a(gate129inter0), .b(s_20), .O(gate129inter1));
  and2  gate303(.a(N360), .b(N14), .O(gate129inter2));
  inv1  gate304(.a(s_20), .O(gate129inter3));
  inv1  gate305(.a(s_21), .O(gate129inter4));
  nand2 gate306(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate307(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate308(.a(N14), .O(gate129inter7));
  inv1  gate309(.a(N360), .O(gate129inter8));
  nand2 gate310(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate311(.a(s_21), .b(gate129inter3), .O(gate129inter10));
  nor2  gate312(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate313(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate314(.a(gate129inter12), .b(gate129inter1), .O(N371));
nand2 gate130( .a(N360), .b(N27), .O(N372) );

  xor2  gate245(.a(N40), .b(N360), .O(gate131inter0));
  nand2 gate246(.a(gate131inter0), .b(s_12), .O(gate131inter1));
  and2  gate247(.a(N40), .b(N360), .O(gate131inter2));
  inv1  gate248(.a(s_12), .O(gate131inter3));
  inv1  gate249(.a(s_13), .O(gate131inter4));
  nand2 gate250(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate251(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate252(.a(N360), .O(gate131inter7));
  inv1  gate253(.a(N40), .O(gate131inter8));
  nand2 gate254(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate255(.a(s_13), .b(gate131inter3), .O(gate131inter10));
  nor2  gate256(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate257(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate258(.a(gate131inter12), .b(gate131inter1), .O(N373));

  xor2  gate413(.a(N53), .b(N360), .O(gate132inter0));
  nand2 gate414(.a(gate132inter0), .b(s_36), .O(gate132inter1));
  and2  gate415(.a(N53), .b(N360), .O(gate132inter2));
  inv1  gate416(.a(s_36), .O(gate132inter3));
  inv1  gate417(.a(s_37), .O(gate132inter4));
  nand2 gate418(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate419(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate420(.a(N360), .O(gate132inter7));
  inv1  gate421(.a(N53), .O(gate132inter8));
  nand2 gate422(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate423(.a(s_37), .b(gate132inter3), .O(gate132inter10));
  nor2  gate424(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate425(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate426(.a(gate132inter12), .b(gate132inter1), .O(N374));
nand2 gate133( .a(N360), .b(N66), .O(N375) );
nand2 gate134( .a(N360), .b(N79), .O(N376) );

  xor2  gate525(.a(N92), .b(N360), .O(gate135inter0));
  nand2 gate526(.a(gate135inter0), .b(s_52), .O(gate135inter1));
  and2  gate527(.a(N92), .b(N360), .O(gate135inter2));
  inv1  gate528(.a(s_52), .O(gate135inter3));
  inv1  gate529(.a(s_53), .O(gate135inter4));
  nand2 gate530(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate531(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate532(.a(N360), .O(gate135inter7));
  inv1  gate533(.a(N92), .O(gate135inter8));
  nand2 gate534(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate535(.a(s_53), .b(gate135inter3), .O(gate135inter10));
  nor2  gate536(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate537(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate538(.a(gate135inter12), .b(gate135inter1), .O(N377));

  xor2  gate175(.a(N105), .b(N360), .O(gate136inter0));
  nand2 gate176(.a(gate136inter0), .b(s_2), .O(gate136inter1));
  and2  gate177(.a(N105), .b(N360), .O(gate136inter2));
  inv1  gate178(.a(s_2), .O(gate136inter3));
  inv1  gate179(.a(s_3), .O(gate136inter4));
  nand2 gate180(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate181(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate182(.a(N360), .O(gate136inter7));
  inv1  gate183(.a(N105), .O(gate136inter8));
  nand2 gate184(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate185(.a(s_3), .b(gate136inter3), .O(gate136inter10));
  nor2  gate186(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate187(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate188(.a(gate136inter12), .b(gate136inter1), .O(N378));

  xor2  gate273(.a(N115), .b(N360), .O(gate137inter0));
  nand2 gate274(.a(gate137inter0), .b(s_16), .O(gate137inter1));
  and2  gate275(.a(N115), .b(N360), .O(gate137inter2));
  inv1  gate276(.a(s_16), .O(gate137inter3));
  inv1  gate277(.a(s_17), .O(gate137inter4));
  nand2 gate278(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate279(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate280(.a(N360), .O(gate137inter7));
  inv1  gate281(.a(N115), .O(gate137inter8));
  nand2 gate282(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate283(.a(s_17), .b(gate137inter3), .O(gate137inter10));
  nor2  gate284(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate285(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate286(.a(gate137inter12), .b(gate137inter1), .O(N379));
nand4 gate138( .a(N4), .b(N242), .c(N334), .d(N371), .O(N380) );
nand4 gate139( .a(N246), .b(N336), .c(N372), .d(N17), .O(N381) );
nand4 gate140( .a(N250), .b(N338), .c(N373), .d(N30), .O(N386) );
nand4 gate141( .a(N254), .b(N340), .c(N374), .d(N43), .O(N393) );
nand4 gate142( .a(N255), .b(N342), .c(N375), .d(N56), .O(N399) );
nand4 gate143( .a(N256), .b(N344), .c(N376), .d(N69), .O(N404) );
nand4 gate144( .a(N257), .b(N345), .c(N377), .d(N82), .O(N407) );
nand4 gate145( .a(N258), .b(N346), .c(N378), .d(N95), .O(N411) );
nand4 gate146( .a(N259), .b(N347), .c(N379), .d(N108), .O(N414) );
inv1 gate147( .a(N380), .O(N415) );
and8 gate148( .a(N381), .b(N386), .c(N393), .d(N399), .e(N404), .f(N407), .g(N411), .h(N414), .O(N416) );
inv1 gate149( .a(N393), .O(N417) );
inv1 gate150( .a(N404), .O(N418) );
inv1 gate151( .a(N407), .O(N419) );
inv1 gate152( .a(N411), .O(N420) );
nor2 gate153( .a(N415), .b(N416), .O(N421) );

  xor2  gate1071(.a(N417), .b(N386), .O(gate154inter0));
  nand2 gate1072(.a(gate154inter0), .b(s_130), .O(gate154inter1));
  and2  gate1073(.a(N417), .b(N386), .O(gate154inter2));
  inv1  gate1074(.a(s_130), .O(gate154inter3));
  inv1  gate1075(.a(s_131), .O(gate154inter4));
  nand2 gate1076(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate1077(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate1078(.a(N386), .O(gate154inter7));
  inv1  gate1079(.a(N417), .O(gate154inter8));
  nand2 gate1080(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate1081(.a(s_131), .b(gate154inter3), .O(gate154inter10));
  nor2  gate1082(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate1083(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate1084(.a(gate154inter12), .b(gate154inter1), .O(N422));
nand4 gate155( .a(N386), .b(N393), .c(N418), .d(N399), .O(N425) );
nand3 gate156( .a(N399), .b(N393), .c(N419), .O(N428) );
nand4 gate157( .a(N386), .b(N393), .c(N407), .d(N420), .O(N429) );
nand4 gate158( .a(N381), .b(N386), .c(N422), .d(N399), .O(N430) );
nand4 gate159( .a(N381), .b(N386), .c(N425), .d(N428), .O(N431) );
nand4 gate160( .a(N381), .b(N422), .c(N425), .d(N429), .O(N432) );

endmodule