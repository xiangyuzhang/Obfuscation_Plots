module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate217inter0, gate217inter1, gate217inter2, gate217inter3, gate217inter4, gate217inter5, gate217inter6, gate217inter7, gate217inter8, gate217inter9, gate217inter10, gate217inter11, gate217inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate1989(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate1990(.a(gate11inter0), .b(s_206), .O(gate11inter1));
  and2  gate1991(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate1992(.a(s_206), .O(gate11inter3));
  inv1  gate1993(.a(s_207), .O(gate11inter4));
  nand2 gate1994(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate1995(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate1996(.a(G5), .O(gate11inter7));
  inv1  gate1997(.a(G6), .O(gate11inter8));
  nand2 gate1998(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate1999(.a(s_207), .b(gate11inter3), .O(gate11inter10));
  nor2  gate2000(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate2001(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate2002(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate827(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate828(.a(gate13inter0), .b(s_40), .O(gate13inter1));
  and2  gate829(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate830(.a(s_40), .O(gate13inter3));
  inv1  gate831(.a(s_41), .O(gate13inter4));
  nand2 gate832(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate833(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate834(.a(G9), .O(gate13inter7));
  inv1  gate835(.a(G10), .O(gate13inter8));
  nand2 gate836(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate837(.a(s_41), .b(gate13inter3), .O(gate13inter10));
  nor2  gate838(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate839(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate840(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate1891(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate1892(.a(gate15inter0), .b(s_192), .O(gate15inter1));
  and2  gate1893(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate1894(.a(s_192), .O(gate15inter3));
  inv1  gate1895(.a(s_193), .O(gate15inter4));
  nand2 gate1896(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate1897(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate1898(.a(G13), .O(gate15inter7));
  inv1  gate1899(.a(G14), .O(gate15inter8));
  nand2 gate1900(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate1901(.a(s_193), .b(gate15inter3), .O(gate15inter10));
  nor2  gate1902(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate1903(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate1904(.a(gate15inter12), .b(gate15inter1), .O(G284));

  xor2  gate1737(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate1738(.a(gate16inter0), .b(s_170), .O(gate16inter1));
  and2  gate1739(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate1740(.a(s_170), .O(gate16inter3));
  inv1  gate1741(.a(s_171), .O(gate16inter4));
  nand2 gate1742(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate1743(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate1744(.a(G15), .O(gate16inter7));
  inv1  gate1745(.a(G16), .O(gate16inter8));
  nand2 gate1746(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate1747(.a(s_171), .b(gate16inter3), .O(gate16inter10));
  nor2  gate1748(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate1749(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate1750(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate547(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate548(.a(gate19inter0), .b(s_0), .O(gate19inter1));
  and2  gate549(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate550(.a(s_0), .O(gate19inter3));
  inv1  gate551(.a(s_1), .O(gate19inter4));
  nand2 gate552(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate553(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate554(.a(G21), .O(gate19inter7));
  inv1  gate555(.a(G22), .O(gate19inter8));
  nand2 gate556(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate557(.a(s_1), .b(gate19inter3), .O(gate19inter10));
  nor2  gate558(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate559(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate560(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate2087(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate2088(.a(gate22inter0), .b(s_220), .O(gate22inter1));
  and2  gate2089(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate2090(.a(s_220), .O(gate22inter3));
  inv1  gate2091(.a(s_221), .O(gate22inter4));
  nand2 gate2092(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate2093(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate2094(.a(G27), .O(gate22inter7));
  inv1  gate2095(.a(G28), .O(gate22inter8));
  nand2 gate2096(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate2097(.a(s_221), .b(gate22inter3), .O(gate22inter10));
  nor2  gate2098(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate2099(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate2100(.a(gate22inter12), .b(gate22inter1), .O(G305));

  xor2  gate1373(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate1374(.a(gate23inter0), .b(s_118), .O(gate23inter1));
  and2  gate1375(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate1376(.a(s_118), .O(gate23inter3));
  inv1  gate1377(.a(s_119), .O(gate23inter4));
  nand2 gate1378(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate1379(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate1380(.a(G29), .O(gate23inter7));
  inv1  gate1381(.a(G30), .O(gate23inter8));
  nand2 gate1382(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate1383(.a(s_119), .b(gate23inter3), .O(gate23inter10));
  nor2  gate1384(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate1385(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate1386(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate897(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate898(.a(gate29inter0), .b(s_50), .O(gate29inter1));
  and2  gate899(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate900(.a(s_50), .O(gate29inter3));
  inv1  gate901(.a(s_51), .O(gate29inter4));
  nand2 gate902(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate903(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate904(.a(G3), .O(gate29inter7));
  inv1  gate905(.a(G7), .O(gate29inter8));
  nand2 gate906(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate907(.a(s_51), .b(gate29inter3), .O(gate29inter10));
  nor2  gate908(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate909(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate910(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );

  xor2  gate757(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate758(.a(gate42inter0), .b(s_30), .O(gate42inter1));
  and2  gate759(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate760(.a(s_30), .O(gate42inter3));
  inv1  gate761(.a(s_31), .O(gate42inter4));
  nand2 gate762(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate763(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate764(.a(G2), .O(gate42inter7));
  inv1  gate765(.a(G266), .O(gate42inter8));
  nand2 gate766(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate767(.a(s_31), .b(gate42inter3), .O(gate42inter10));
  nor2  gate768(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate769(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate770(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );

  xor2  gate1387(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate1388(.a(gate45inter0), .b(s_120), .O(gate45inter1));
  and2  gate1389(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate1390(.a(s_120), .O(gate45inter3));
  inv1  gate1391(.a(s_121), .O(gate45inter4));
  nand2 gate1392(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate1393(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate1394(.a(G5), .O(gate45inter7));
  inv1  gate1395(.a(G272), .O(gate45inter8));
  nand2 gate1396(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate1397(.a(s_121), .b(gate45inter3), .O(gate45inter10));
  nor2  gate1398(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate1399(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate1400(.a(gate45inter12), .b(gate45inter1), .O(G366));
nand2 gate46( .a(G6), .b(G272), .O(G367) );

  xor2  gate995(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate996(.a(gate47inter0), .b(s_64), .O(gate47inter1));
  and2  gate997(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate998(.a(s_64), .O(gate47inter3));
  inv1  gate999(.a(s_65), .O(gate47inter4));
  nand2 gate1000(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate1001(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate1002(.a(G7), .O(gate47inter7));
  inv1  gate1003(.a(G275), .O(gate47inter8));
  nand2 gate1004(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate1005(.a(s_65), .b(gate47inter3), .O(gate47inter10));
  nor2  gate1006(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate1007(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate1008(.a(gate47inter12), .b(gate47inter1), .O(G368));
nand2 gate48( .a(G8), .b(G275), .O(G369) );

  xor2  gate603(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate604(.a(gate49inter0), .b(s_8), .O(gate49inter1));
  and2  gate605(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate606(.a(s_8), .O(gate49inter3));
  inv1  gate607(.a(s_9), .O(gate49inter4));
  nand2 gate608(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate609(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate610(.a(G9), .O(gate49inter7));
  inv1  gate611(.a(G278), .O(gate49inter8));
  nand2 gate612(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate613(.a(s_9), .b(gate49inter3), .O(gate49inter10));
  nor2  gate614(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate615(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate616(.a(gate49inter12), .b(gate49inter1), .O(G370));
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate1317(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate1318(.a(gate51inter0), .b(s_110), .O(gate51inter1));
  and2  gate1319(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate1320(.a(s_110), .O(gate51inter3));
  inv1  gate1321(.a(s_111), .O(gate51inter4));
  nand2 gate1322(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate1323(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate1324(.a(G11), .O(gate51inter7));
  inv1  gate1325(.a(G281), .O(gate51inter8));
  nand2 gate1326(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate1327(.a(s_111), .b(gate51inter3), .O(gate51inter10));
  nor2  gate1328(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate1329(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate1330(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate883(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate884(.a(gate55inter0), .b(s_48), .O(gate55inter1));
  and2  gate885(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate886(.a(s_48), .O(gate55inter3));
  inv1  gate887(.a(s_49), .O(gate55inter4));
  nand2 gate888(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate889(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate890(.a(G15), .O(gate55inter7));
  inv1  gate891(.a(G287), .O(gate55inter8));
  nand2 gate892(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate893(.a(s_49), .b(gate55inter3), .O(gate55inter10));
  nor2  gate894(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate895(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate896(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate1835(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate1836(.a(gate60inter0), .b(s_184), .O(gate60inter1));
  and2  gate1837(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate1838(.a(s_184), .O(gate60inter3));
  inv1  gate1839(.a(s_185), .O(gate60inter4));
  nand2 gate1840(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate1841(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate1842(.a(G20), .O(gate60inter7));
  inv1  gate1843(.a(G293), .O(gate60inter8));
  nand2 gate1844(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate1845(.a(s_185), .b(gate60inter3), .O(gate60inter10));
  nor2  gate1846(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate1847(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate1848(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );

  xor2  gate2269(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate2270(.a(gate64inter0), .b(s_246), .O(gate64inter1));
  and2  gate2271(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate2272(.a(s_246), .O(gate64inter3));
  inv1  gate2273(.a(s_247), .O(gate64inter4));
  nand2 gate2274(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate2275(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate2276(.a(G24), .O(gate64inter7));
  inv1  gate2277(.a(G299), .O(gate64inter8));
  nand2 gate2278(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate2279(.a(s_247), .b(gate64inter3), .O(gate64inter10));
  nor2  gate2280(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate2281(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate2282(.a(gate64inter12), .b(gate64inter1), .O(G385));

  xor2  gate2059(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate2060(.a(gate65inter0), .b(s_216), .O(gate65inter1));
  and2  gate2061(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate2062(.a(s_216), .O(gate65inter3));
  inv1  gate2063(.a(s_217), .O(gate65inter4));
  nand2 gate2064(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate2065(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate2066(.a(G25), .O(gate65inter7));
  inv1  gate2067(.a(G302), .O(gate65inter8));
  nand2 gate2068(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate2069(.a(s_217), .b(gate65inter3), .O(gate65inter10));
  nor2  gate2070(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate2071(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate2072(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate743(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate744(.a(gate69inter0), .b(s_28), .O(gate69inter1));
  and2  gate745(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate746(.a(s_28), .O(gate69inter3));
  inv1  gate747(.a(s_29), .O(gate69inter4));
  nand2 gate748(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate749(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate750(.a(G29), .O(gate69inter7));
  inv1  gate751(.a(G308), .O(gate69inter8));
  nand2 gate752(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate753(.a(s_29), .b(gate69inter3), .O(gate69inter10));
  nor2  gate754(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate755(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate756(.a(gate69inter12), .b(gate69inter1), .O(G390));

  xor2  gate1751(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate1752(.a(gate70inter0), .b(s_172), .O(gate70inter1));
  and2  gate1753(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate1754(.a(s_172), .O(gate70inter3));
  inv1  gate1755(.a(s_173), .O(gate70inter4));
  nand2 gate1756(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate1757(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate1758(.a(G30), .O(gate70inter7));
  inv1  gate1759(.a(G308), .O(gate70inter8));
  nand2 gate1760(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate1761(.a(s_173), .b(gate70inter3), .O(gate70inter10));
  nor2  gate1762(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate1763(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate1764(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );

  xor2  gate2255(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate2256(.a(gate72inter0), .b(s_244), .O(gate72inter1));
  and2  gate2257(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate2258(.a(s_244), .O(gate72inter3));
  inv1  gate2259(.a(s_245), .O(gate72inter4));
  nand2 gate2260(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate2261(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate2262(.a(G32), .O(gate72inter7));
  inv1  gate2263(.a(G311), .O(gate72inter8));
  nand2 gate2264(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate2265(.a(s_245), .b(gate72inter3), .O(gate72inter10));
  nor2  gate2266(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate2267(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate2268(.a(gate72inter12), .b(gate72inter1), .O(G393));
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate1065(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate1066(.a(gate75inter0), .b(s_74), .O(gate75inter1));
  and2  gate1067(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate1068(.a(s_74), .O(gate75inter3));
  inv1  gate1069(.a(s_75), .O(gate75inter4));
  nand2 gate1070(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate1071(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate1072(.a(G9), .O(gate75inter7));
  inv1  gate1073(.a(G317), .O(gate75inter8));
  nand2 gate1074(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate1075(.a(s_75), .b(gate75inter3), .O(gate75inter10));
  nor2  gate1076(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate1077(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate1078(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate869(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate870(.a(gate82inter0), .b(s_46), .O(gate82inter1));
  and2  gate871(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate872(.a(s_46), .O(gate82inter3));
  inv1  gate873(.a(s_47), .O(gate82inter4));
  nand2 gate874(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate875(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate876(.a(G7), .O(gate82inter7));
  inv1  gate877(.a(G326), .O(gate82inter8));
  nand2 gate878(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate879(.a(s_47), .b(gate82inter3), .O(gate82inter10));
  nor2  gate880(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate881(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate882(.a(gate82inter12), .b(gate82inter1), .O(G403));

  xor2  gate2213(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate2214(.a(gate83inter0), .b(s_238), .O(gate83inter1));
  and2  gate2215(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate2216(.a(s_238), .O(gate83inter3));
  inv1  gate2217(.a(s_239), .O(gate83inter4));
  nand2 gate2218(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate2219(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate2220(.a(G11), .O(gate83inter7));
  inv1  gate2221(.a(G329), .O(gate83inter8));
  nand2 gate2222(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate2223(.a(s_239), .b(gate83inter3), .O(gate83inter10));
  nor2  gate2224(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate2225(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate2226(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );

  xor2  gate1877(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate1878(.a(gate87inter0), .b(s_190), .O(gate87inter1));
  and2  gate1879(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate1880(.a(s_190), .O(gate87inter3));
  inv1  gate1881(.a(s_191), .O(gate87inter4));
  nand2 gate1882(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate1883(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate1884(.a(G12), .O(gate87inter7));
  inv1  gate1885(.a(G335), .O(gate87inter8));
  nand2 gate1886(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate1887(.a(s_191), .b(gate87inter3), .O(gate87inter10));
  nor2  gate1888(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate1889(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate1890(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );

  xor2  gate1709(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate1710(.a(gate89inter0), .b(s_166), .O(gate89inter1));
  and2  gate1711(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate1712(.a(s_166), .O(gate89inter3));
  inv1  gate1713(.a(s_167), .O(gate89inter4));
  nand2 gate1714(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate1715(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate1716(.a(G17), .O(gate89inter7));
  inv1  gate1717(.a(G338), .O(gate89inter8));
  nand2 gate1718(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate1719(.a(s_167), .b(gate89inter3), .O(gate89inter10));
  nor2  gate1720(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate1721(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate1722(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate1569(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate1570(.a(gate91inter0), .b(s_146), .O(gate91inter1));
  and2  gate1571(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate1572(.a(s_146), .O(gate91inter3));
  inv1  gate1573(.a(s_147), .O(gate91inter4));
  nand2 gate1574(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate1575(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate1576(.a(G25), .O(gate91inter7));
  inv1  gate1577(.a(G341), .O(gate91inter8));
  nand2 gate1578(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate1579(.a(s_147), .b(gate91inter3), .O(gate91inter10));
  nor2  gate1580(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate1581(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate1582(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );

  xor2  gate673(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate674(.a(gate93inter0), .b(s_18), .O(gate93inter1));
  and2  gate675(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate676(.a(s_18), .O(gate93inter3));
  inv1  gate677(.a(s_19), .O(gate93inter4));
  nand2 gate678(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate679(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate680(.a(G18), .O(gate93inter7));
  inv1  gate681(.a(G344), .O(gate93inter8));
  nand2 gate682(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate683(.a(s_19), .b(gate93inter3), .O(gate93inter10));
  nor2  gate684(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate685(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate686(.a(gate93inter12), .b(gate93inter1), .O(G414));

  xor2  gate785(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate786(.a(gate94inter0), .b(s_34), .O(gate94inter1));
  and2  gate787(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate788(.a(s_34), .O(gate94inter3));
  inv1  gate789(.a(s_35), .O(gate94inter4));
  nand2 gate790(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate791(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate792(.a(G22), .O(gate94inter7));
  inv1  gate793(.a(G344), .O(gate94inter8));
  nand2 gate794(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate795(.a(s_35), .b(gate94inter3), .O(gate94inter10));
  nor2  gate796(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate797(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate798(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );

  xor2  gate715(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate716(.a(gate97inter0), .b(s_24), .O(gate97inter1));
  and2  gate717(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate718(.a(s_24), .O(gate97inter3));
  inv1  gate719(.a(s_25), .O(gate97inter4));
  nand2 gate720(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate721(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate722(.a(G19), .O(gate97inter7));
  inv1  gate723(.a(G350), .O(gate97inter8));
  nand2 gate724(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate725(.a(s_25), .b(gate97inter3), .O(gate97inter10));
  nor2  gate726(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate727(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate728(.a(gate97inter12), .b(gate97inter1), .O(G418));

  xor2  gate589(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate590(.a(gate98inter0), .b(s_6), .O(gate98inter1));
  and2  gate591(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate592(.a(s_6), .O(gate98inter3));
  inv1  gate593(.a(s_7), .O(gate98inter4));
  nand2 gate594(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate595(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate596(.a(G23), .O(gate98inter7));
  inv1  gate597(.a(G350), .O(gate98inter8));
  nand2 gate598(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate599(.a(s_7), .b(gate98inter3), .O(gate98inter10));
  nor2  gate600(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate601(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate602(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate855(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate856(.a(gate100inter0), .b(s_44), .O(gate100inter1));
  and2  gate857(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate858(.a(s_44), .O(gate100inter3));
  inv1  gate859(.a(s_45), .O(gate100inter4));
  nand2 gate860(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate861(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate862(.a(G31), .O(gate100inter7));
  inv1  gate863(.a(G353), .O(gate100inter8));
  nand2 gate864(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate865(.a(s_45), .b(gate100inter3), .O(gate100inter10));
  nor2  gate866(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate867(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate868(.a(gate100inter12), .b(gate100inter1), .O(G421));

  xor2  gate1653(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate1654(.a(gate101inter0), .b(s_158), .O(gate101inter1));
  and2  gate1655(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate1656(.a(s_158), .O(gate101inter3));
  inv1  gate1657(.a(s_159), .O(gate101inter4));
  nand2 gate1658(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate1659(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate1660(.a(G20), .O(gate101inter7));
  inv1  gate1661(.a(G356), .O(gate101inter8));
  nand2 gate1662(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate1663(.a(s_159), .b(gate101inter3), .O(gate101inter10));
  nor2  gate1664(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate1665(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate1666(.a(gate101inter12), .b(gate101inter1), .O(G422));
nand2 gate102( .a(G24), .b(G356), .O(G423) );

  xor2  gate1135(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate1136(.a(gate103inter0), .b(s_84), .O(gate103inter1));
  and2  gate1137(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate1138(.a(s_84), .O(gate103inter3));
  inv1  gate1139(.a(s_85), .O(gate103inter4));
  nand2 gate1140(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate1141(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate1142(.a(G28), .O(gate103inter7));
  inv1  gate1143(.a(G359), .O(gate103inter8));
  nand2 gate1144(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate1145(.a(s_85), .b(gate103inter3), .O(gate103inter10));
  nor2  gate1146(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate1147(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate1148(.a(gate103inter12), .b(gate103inter1), .O(G424));
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate2241(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate2242(.a(gate108inter0), .b(s_242), .O(gate108inter1));
  and2  gate2243(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate2244(.a(s_242), .O(gate108inter3));
  inv1  gate2245(.a(s_243), .O(gate108inter4));
  nand2 gate2246(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate2247(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate2248(.a(G368), .O(gate108inter7));
  inv1  gate2249(.a(G369), .O(gate108inter8));
  nand2 gate2250(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate2251(.a(s_243), .b(gate108inter3), .O(gate108inter10));
  nor2  gate2252(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate2253(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate2254(.a(gate108inter12), .b(gate108inter1), .O(G435));

  xor2  gate1037(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate1038(.a(gate109inter0), .b(s_70), .O(gate109inter1));
  and2  gate1039(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate1040(.a(s_70), .O(gate109inter3));
  inv1  gate1041(.a(s_71), .O(gate109inter4));
  nand2 gate1042(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate1043(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate1044(.a(G370), .O(gate109inter7));
  inv1  gate1045(.a(G371), .O(gate109inter8));
  nand2 gate1046(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate1047(.a(s_71), .b(gate109inter3), .O(gate109inter10));
  nor2  gate1048(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate1049(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate1050(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );

  xor2  gate1401(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate1402(.a(gate111inter0), .b(s_122), .O(gate111inter1));
  and2  gate1403(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate1404(.a(s_122), .O(gate111inter3));
  inv1  gate1405(.a(s_123), .O(gate111inter4));
  nand2 gate1406(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate1407(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate1408(.a(G374), .O(gate111inter7));
  inv1  gate1409(.a(G375), .O(gate111inter8));
  nand2 gate1410(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate1411(.a(s_123), .b(gate111inter3), .O(gate111inter10));
  nor2  gate1412(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate1413(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate1414(.a(gate111inter12), .b(gate111inter1), .O(G444));
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate939(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate940(.a(gate124inter0), .b(s_56), .O(gate124inter1));
  and2  gate941(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate942(.a(s_56), .O(gate124inter3));
  inv1  gate943(.a(s_57), .O(gate124inter4));
  nand2 gate944(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate945(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate946(.a(G400), .O(gate124inter7));
  inv1  gate947(.a(G401), .O(gate124inter8));
  nand2 gate948(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate949(.a(s_57), .b(gate124inter3), .O(gate124inter10));
  nor2  gate950(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate951(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate952(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate687(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate688(.a(gate126inter0), .b(s_20), .O(gate126inter1));
  and2  gate689(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate690(.a(s_20), .O(gate126inter3));
  inv1  gate691(.a(s_21), .O(gate126inter4));
  nand2 gate692(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate693(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate694(.a(G404), .O(gate126inter7));
  inv1  gate695(.a(G405), .O(gate126inter8));
  nand2 gate696(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate697(.a(s_21), .b(gate126inter3), .O(gate126inter10));
  nor2  gate698(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate699(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate700(.a(gate126inter12), .b(gate126inter1), .O(G489));

  xor2  gate925(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate926(.a(gate127inter0), .b(s_54), .O(gate127inter1));
  and2  gate927(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate928(.a(s_54), .O(gate127inter3));
  inv1  gate929(.a(s_55), .O(gate127inter4));
  nand2 gate930(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate931(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate932(.a(G406), .O(gate127inter7));
  inv1  gate933(.a(G407), .O(gate127inter8));
  nand2 gate934(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate935(.a(s_55), .b(gate127inter3), .O(gate127inter10));
  nor2  gate936(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate937(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate938(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );

  xor2  gate1191(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate1192(.a(gate130inter0), .b(s_92), .O(gate130inter1));
  and2  gate1193(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate1194(.a(s_92), .O(gate130inter3));
  inv1  gate1195(.a(s_93), .O(gate130inter4));
  nand2 gate1196(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate1197(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate1198(.a(G412), .O(gate130inter7));
  inv1  gate1199(.a(G413), .O(gate130inter8));
  nand2 gate1200(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate1201(.a(s_93), .b(gate130inter3), .O(gate130inter10));
  nor2  gate1202(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate1203(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate1204(.a(gate130inter12), .b(gate130inter1), .O(G501));
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );

  xor2  gate1597(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate1598(.a(gate133inter0), .b(s_150), .O(gate133inter1));
  and2  gate1599(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate1600(.a(s_150), .O(gate133inter3));
  inv1  gate1601(.a(s_151), .O(gate133inter4));
  nand2 gate1602(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate1603(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate1604(.a(G418), .O(gate133inter7));
  inv1  gate1605(.a(G419), .O(gate133inter8));
  nand2 gate1606(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate1607(.a(s_151), .b(gate133inter3), .O(gate133inter10));
  nor2  gate1608(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate1609(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate1610(.a(gate133inter12), .b(gate133inter1), .O(G510));
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate1765(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate1766(.a(gate136inter0), .b(s_174), .O(gate136inter1));
  and2  gate1767(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate1768(.a(s_174), .O(gate136inter3));
  inv1  gate1769(.a(s_175), .O(gate136inter4));
  nand2 gate1770(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate1771(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate1772(.a(G424), .O(gate136inter7));
  inv1  gate1773(.a(G425), .O(gate136inter8));
  nand2 gate1774(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate1775(.a(s_175), .b(gate136inter3), .O(gate136inter10));
  nor2  gate1776(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate1777(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate1778(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate1121(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate1122(.a(gate138inter0), .b(s_82), .O(gate138inter1));
  and2  gate1123(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate1124(.a(s_82), .O(gate138inter3));
  inv1  gate1125(.a(s_83), .O(gate138inter4));
  nand2 gate1126(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate1127(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate1128(.a(G432), .O(gate138inter7));
  inv1  gate1129(.a(G435), .O(gate138inter8));
  nand2 gate1130(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate1131(.a(s_83), .b(gate138inter3), .O(gate138inter10));
  nor2  gate1132(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate1133(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate1134(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );

  xor2  gate953(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate954(.a(gate140inter0), .b(s_58), .O(gate140inter1));
  and2  gate955(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate956(.a(s_58), .O(gate140inter3));
  inv1  gate957(.a(s_59), .O(gate140inter4));
  nand2 gate958(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate959(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate960(.a(G444), .O(gate140inter7));
  inv1  gate961(.a(G447), .O(gate140inter8));
  nand2 gate962(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate963(.a(s_59), .b(gate140inter3), .O(gate140inter10));
  nor2  gate964(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate965(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate966(.a(gate140inter12), .b(gate140inter1), .O(G531));
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate2157(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate2158(.a(gate143inter0), .b(s_230), .O(gate143inter1));
  and2  gate2159(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate2160(.a(s_230), .O(gate143inter3));
  inv1  gate2161(.a(s_231), .O(gate143inter4));
  nand2 gate2162(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate2163(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate2164(.a(G462), .O(gate143inter7));
  inv1  gate2165(.a(G465), .O(gate143inter8));
  nand2 gate2166(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate2167(.a(s_231), .b(gate143inter3), .O(gate143inter10));
  nor2  gate2168(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate2169(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate2170(.a(gate143inter12), .b(gate143inter1), .O(G540));

  xor2  gate1625(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate1626(.a(gate144inter0), .b(s_154), .O(gate144inter1));
  and2  gate1627(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate1628(.a(s_154), .O(gate144inter3));
  inv1  gate1629(.a(s_155), .O(gate144inter4));
  nand2 gate1630(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate1631(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate1632(.a(G468), .O(gate144inter7));
  inv1  gate1633(.a(G471), .O(gate144inter8));
  nand2 gate1634(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate1635(.a(s_155), .b(gate144inter3), .O(gate144inter10));
  nor2  gate1636(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate1637(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate1638(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );

  xor2  gate1849(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate1850(.a(gate146inter0), .b(s_186), .O(gate146inter1));
  and2  gate1851(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate1852(.a(s_186), .O(gate146inter3));
  inv1  gate1853(.a(s_187), .O(gate146inter4));
  nand2 gate1854(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate1855(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate1856(.a(G480), .O(gate146inter7));
  inv1  gate1857(.a(G483), .O(gate146inter8));
  nand2 gate1858(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate1859(.a(s_187), .b(gate146inter3), .O(gate146inter10));
  nor2  gate1860(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate1861(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate1862(.a(gate146inter12), .b(gate146inter1), .O(G549));
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate1443(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate1444(.a(gate161inter0), .b(s_128), .O(gate161inter1));
  and2  gate1445(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate1446(.a(s_128), .O(gate161inter3));
  inv1  gate1447(.a(s_129), .O(gate161inter4));
  nand2 gate1448(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate1449(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate1450(.a(G450), .O(gate161inter7));
  inv1  gate1451(.a(G534), .O(gate161inter8));
  nand2 gate1452(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate1453(.a(s_129), .b(gate161inter3), .O(gate161inter10));
  nor2  gate1454(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate1455(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate1456(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );

  xor2  gate771(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate772(.a(gate163inter0), .b(s_32), .O(gate163inter1));
  and2  gate773(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate774(.a(s_32), .O(gate163inter3));
  inv1  gate775(.a(s_33), .O(gate163inter4));
  nand2 gate776(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate777(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate778(.a(G456), .O(gate163inter7));
  inv1  gate779(.a(G537), .O(gate163inter8));
  nand2 gate780(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate781(.a(s_33), .b(gate163inter3), .O(gate163inter10));
  nor2  gate782(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate783(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate784(.a(gate163inter12), .b(gate163inter1), .O(G580));

  xor2  gate659(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate660(.a(gate164inter0), .b(s_16), .O(gate164inter1));
  and2  gate661(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate662(.a(s_16), .O(gate164inter3));
  inv1  gate663(.a(s_17), .O(gate164inter4));
  nand2 gate664(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate665(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate666(.a(G459), .O(gate164inter7));
  inv1  gate667(.a(G537), .O(gate164inter8));
  nand2 gate668(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate669(.a(s_17), .b(gate164inter3), .O(gate164inter10));
  nor2  gate670(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate671(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate672(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );

  xor2  gate2171(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate2172(.a(gate166inter0), .b(s_232), .O(gate166inter1));
  and2  gate2173(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate2174(.a(s_232), .O(gate166inter3));
  inv1  gate2175(.a(s_233), .O(gate166inter4));
  nand2 gate2176(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate2177(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate2178(.a(G465), .O(gate166inter7));
  inv1  gate2179(.a(G540), .O(gate166inter8));
  nand2 gate2180(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate2181(.a(s_233), .b(gate166inter3), .O(gate166inter10));
  nor2  gate2182(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate2183(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate2184(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate1947(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate1948(.a(gate170inter0), .b(s_200), .O(gate170inter1));
  and2  gate1949(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate1950(.a(s_200), .O(gate170inter3));
  inv1  gate1951(.a(s_201), .O(gate170inter4));
  nand2 gate1952(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate1953(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate1954(.a(G477), .O(gate170inter7));
  inv1  gate1955(.a(G546), .O(gate170inter8));
  nand2 gate1956(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate1957(.a(s_201), .b(gate170inter3), .O(gate170inter10));
  nor2  gate1958(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate1959(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate1960(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate1359(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate1360(.a(gate178inter0), .b(s_116), .O(gate178inter1));
  and2  gate1361(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate1362(.a(s_116), .O(gate178inter3));
  inv1  gate1363(.a(s_117), .O(gate178inter4));
  nand2 gate1364(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate1365(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate1366(.a(G501), .O(gate178inter7));
  inv1  gate1367(.a(G558), .O(gate178inter8));
  nand2 gate1368(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate1369(.a(s_117), .b(gate178inter3), .O(gate178inter10));
  nor2  gate1370(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate1371(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate1372(.a(gate178inter12), .b(gate178inter1), .O(G595));
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate1779(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate1780(.a(gate187inter0), .b(s_176), .O(gate187inter1));
  and2  gate1781(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate1782(.a(s_176), .O(gate187inter3));
  inv1  gate1783(.a(s_177), .O(gate187inter4));
  nand2 gate1784(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate1785(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate1786(.a(G574), .O(gate187inter7));
  inv1  gate1787(.a(G575), .O(gate187inter8));
  nand2 gate1788(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate1789(.a(s_177), .b(gate187inter3), .O(gate187inter10));
  nor2  gate1790(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate1791(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate1792(.a(gate187inter12), .b(gate187inter1), .O(G612));

  xor2  gate1919(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate1920(.a(gate188inter0), .b(s_196), .O(gate188inter1));
  and2  gate1921(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate1922(.a(s_196), .O(gate188inter3));
  inv1  gate1923(.a(s_197), .O(gate188inter4));
  nand2 gate1924(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate1925(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate1926(.a(G576), .O(gate188inter7));
  inv1  gate1927(.a(G577), .O(gate188inter8));
  nand2 gate1928(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate1929(.a(s_197), .b(gate188inter3), .O(gate188inter10));
  nor2  gate1930(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate1931(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate1932(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate2101(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate2102(.a(gate193inter0), .b(s_222), .O(gate193inter1));
  and2  gate2103(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate2104(.a(s_222), .O(gate193inter3));
  inv1  gate2105(.a(s_223), .O(gate193inter4));
  nand2 gate2106(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate2107(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate2108(.a(G586), .O(gate193inter7));
  inv1  gate2109(.a(G587), .O(gate193inter8));
  nand2 gate2110(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate2111(.a(s_223), .b(gate193inter3), .O(gate193inter10));
  nor2  gate2112(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate2113(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate2114(.a(gate193inter12), .b(gate193inter1), .O(G642));

  xor2  gate2367(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate2368(.a(gate194inter0), .b(s_260), .O(gate194inter1));
  and2  gate2369(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate2370(.a(s_260), .O(gate194inter3));
  inv1  gate2371(.a(s_261), .O(gate194inter4));
  nand2 gate2372(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate2373(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate2374(.a(G588), .O(gate194inter7));
  inv1  gate2375(.a(G589), .O(gate194inter8));
  nand2 gate2376(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate2377(.a(s_261), .b(gate194inter3), .O(gate194inter10));
  nor2  gate2378(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate2379(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate2380(.a(gate194inter12), .b(gate194inter1), .O(G645));

  xor2  gate1205(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate1206(.a(gate195inter0), .b(s_94), .O(gate195inter1));
  and2  gate1207(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate1208(.a(s_94), .O(gate195inter3));
  inv1  gate1209(.a(s_95), .O(gate195inter4));
  nand2 gate1210(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate1211(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate1212(.a(G590), .O(gate195inter7));
  inv1  gate1213(.a(G591), .O(gate195inter8));
  nand2 gate1214(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate1215(.a(s_95), .b(gate195inter3), .O(gate195inter10));
  nor2  gate1216(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate1217(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate1218(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate1009(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate1010(.a(gate201inter0), .b(s_66), .O(gate201inter1));
  and2  gate1011(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate1012(.a(s_66), .O(gate201inter3));
  inv1  gate1013(.a(s_67), .O(gate201inter4));
  nand2 gate1014(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate1015(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate1016(.a(G602), .O(gate201inter7));
  inv1  gate1017(.a(G607), .O(gate201inter8));
  nand2 gate1018(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate1019(.a(s_67), .b(gate201inter3), .O(gate201inter10));
  nor2  gate1020(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate1021(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate1022(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate1471(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate1472(.a(gate205inter0), .b(s_132), .O(gate205inter1));
  and2  gate1473(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate1474(.a(s_132), .O(gate205inter3));
  inv1  gate1475(.a(s_133), .O(gate205inter4));
  nand2 gate1476(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate1477(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate1478(.a(G622), .O(gate205inter7));
  inv1  gate1479(.a(G627), .O(gate205inter8));
  nand2 gate1480(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate1481(.a(s_133), .b(gate205inter3), .O(gate205inter10));
  nor2  gate1482(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate1483(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate1484(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate1821(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate1822(.a(gate211inter0), .b(s_182), .O(gate211inter1));
  and2  gate1823(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate1824(.a(s_182), .O(gate211inter3));
  inv1  gate1825(.a(s_183), .O(gate211inter4));
  nand2 gate1826(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate1827(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate1828(.a(G612), .O(gate211inter7));
  inv1  gate1829(.a(G669), .O(gate211inter8));
  nand2 gate1830(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate1831(.a(s_183), .b(gate211inter3), .O(gate211inter10));
  nor2  gate1832(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate1833(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate1834(.a(gate211inter12), .b(gate211inter1), .O(G692));
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate1275(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate1276(.a(gate214inter0), .b(s_104), .O(gate214inter1));
  and2  gate1277(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate1278(.a(s_104), .O(gate214inter3));
  inv1  gate1279(.a(s_105), .O(gate214inter4));
  nand2 gate1280(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate1281(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate1282(.a(G612), .O(gate214inter7));
  inv1  gate1283(.a(G672), .O(gate214inter8));
  nand2 gate1284(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate1285(.a(s_105), .b(gate214inter3), .O(gate214inter10));
  nor2  gate1286(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate1287(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate1288(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate1429(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate1430(.a(gate216inter0), .b(s_126), .O(gate216inter1));
  and2  gate1431(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate1432(.a(s_126), .O(gate216inter3));
  inv1  gate1433(.a(s_127), .O(gate216inter4));
  nand2 gate1434(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate1435(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate1436(.a(G617), .O(gate216inter7));
  inv1  gate1437(.a(G675), .O(gate216inter8));
  nand2 gate1438(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate1439(.a(s_127), .b(gate216inter3), .O(gate216inter10));
  nor2  gate1440(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate1441(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate1442(.a(gate216inter12), .b(gate216inter1), .O(G697));

  xor2  gate1457(.a(G678), .b(G622), .O(gate217inter0));
  nand2 gate1458(.a(gate217inter0), .b(s_130), .O(gate217inter1));
  and2  gate1459(.a(G678), .b(G622), .O(gate217inter2));
  inv1  gate1460(.a(s_130), .O(gate217inter3));
  inv1  gate1461(.a(s_131), .O(gate217inter4));
  nand2 gate1462(.a(gate217inter4), .b(gate217inter3), .O(gate217inter5));
  nor2  gate1463(.a(gate217inter5), .b(gate217inter2), .O(gate217inter6));
  inv1  gate1464(.a(G622), .O(gate217inter7));
  inv1  gate1465(.a(G678), .O(gate217inter8));
  nand2 gate1466(.a(gate217inter8), .b(gate217inter7), .O(gate217inter9));
  nand2 gate1467(.a(s_131), .b(gate217inter3), .O(gate217inter10));
  nor2  gate1468(.a(gate217inter10), .b(gate217inter9), .O(gate217inter11));
  nor2  gate1469(.a(gate217inter11), .b(gate217inter6), .O(gate217inter12));
  nand2 gate1470(.a(gate217inter12), .b(gate217inter1), .O(G698));
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate1051(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate1052(.a(gate219inter0), .b(s_72), .O(gate219inter1));
  and2  gate1053(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate1054(.a(s_72), .O(gate219inter3));
  inv1  gate1055(.a(s_73), .O(gate219inter4));
  nand2 gate1056(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate1057(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate1058(.a(G632), .O(gate219inter7));
  inv1  gate1059(.a(G681), .O(gate219inter8));
  nand2 gate1060(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate1061(.a(s_73), .b(gate219inter3), .O(gate219inter10));
  nor2  gate1062(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate1063(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate1064(.a(gate219inter12), .b(gate219inter1), .O(G700));

  xor2  gate1639(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate1640(.a(gate220inter0), .b(s_156), .O(gate220inter1));
  and2  gate1641(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate1642(.a(s_156), .O(gate220inter3));
  inv1  gate1643(.a(s_157), .O(gate220inter4));
  nand2 gate1644(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate1645(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate1646(.a(G637), .O(gate220inter7));
  inv1  gate1647(.a(G681), .O(gate220inter8));
  nand2 gate1648(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate1649(.a(s_157), .b(gate220inter3), .O(gate220inter10));
  nor2  gate1650(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate1651(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate1652(.a(gate220inter12), .b(gate220inter1), .O(G701));
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate841(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate842(.a(gate228inter0), .b(s_42), .O(gate228inter1));
  and2  gate843(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate844(.a(s_42), .O(gate228inter3));
  inv1  gate845(.a(s_43), .O(gate228inter4));
  nand2 gate846(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate847(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate848(.a(G696), .O(gate228inter7));
  inv1  gate849(.a(G697), .O(gate228inter8));
  nand2 gate850(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate851(.a(s_43), .b(gate228inter3), .O(gate228inter10));
  nor2  gate852(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate853(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate854(.a(gate228inter12), .b(gate228inter1), .O(G715));

  xor2  gate2199(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate2200(.a(gate229inter0), .b(s_236), .O(gate229inter1));
  and2  gate2201(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate2202(.a(s_236), .O(gate229inter3));
  inv1  gate2203(.a(s_237), .O(gate229inter4));
  nand2 gate2204(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate2205(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate2206(.a(G698), .O(gate229inter7));
  inv1  gate2207(.a(G699), .O(gate229inter8));
  nand2 gate2208(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate2209(.a(s_237), .b(gate229inter3), .O(gate229inter10));
  nor2  gate2210(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate2211(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate2212(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate2129(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate2130(.a(gate231inter0), .b(s_226), .O(gate231inter1));
  and2  gate2131(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate2132(.a(s_226), .O(gate231inter3));
  inv1  gate2133(.a(s_227), .O(gate231inter4));
  nand2 gate2134(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate2135(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate2136(.a(G702), .O(gate231inter7));
  inv1  gate2137(.a(G703), .O(gate231inter8));
  nand2 gate2138(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate2139(.a(s_227), .b(gate231inter3), .O(gate231inter10));
  nor2  gate2140(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate2141(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate2142(.a(gate231inter12), .b(gate231inter1), .O(G724));

  xor2  gate1233(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate1234(.a(gate232inter0), .b(s_98), .O(gate232inter1));
  and2  gate1235(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate1236(.a(s_98), .O(gate232inter3));
  inv1  gate1237(.a(s_99), .O(gate232inter4));
  nand2 gate1238(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate1239(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate1240(.a(G704), .O(gate232inter7));
  inv1  gate1241(.a(G705), .O(gate232inter8));
  nand2 gate1242(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate1243(.a(s_99), .b(gate232inter3), .O(gate232inter10));
  nor2  gate1244(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate1245(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate1246(.a(gate232inter12), .b(gate232inter1), .O(G727));
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate1163(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate1164(.a(gate236inter0), .b(s_88), .O(gate236inter1));
  and2  gate1165(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate1166(.a(s_88), .O(gate236inter3));
  inv1  gate1167(.a(s_89), .O(gate236inter4));
  nand2 gate1168(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate1169(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate1170(.a(G251), .O(gate236inter7));
  inv1  gate1171(.a(G727), .O(gate236inter8));
  nand2 gate1172(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate1173(.a(s_89), .b(gate236inter3), .O(gate236inter10));
  nor2  gate1174(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate1175(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate1176(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate1219(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate1220(.a(gate245inter0), .b(s_96), .O(gate245inter1));
  and2  gate1221(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate1222(.a(s_96), .O(gate245inter3));
  inv1  gate1223(.a(s_97), .O(gate245inter4));
  nand2 gate1224(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate1225(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate1226(.a(G248), .O(gate245inter7));
  inv1  gate1227(.a(G736), .O(gate245inter8));
  nand2 gate1228(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate1229(.a(s_97), .b(gate245inter3), .O(gate245inter10));
  nor2  gate1230(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate1231(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate1232(.a(gate245inter12), .b(gate245inter1), .O(G758));

  xor2  gate2003(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate2004(.a(gate246inter0), .b(s_208), .O(gate246inter1));
  and2  gate2005(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate2006(.a(s_208), .O(gate246inter3));
  inv1  gate2007(.a(s_209), .O(gate246inter4));
  nand2 gate2008(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate2009(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate2010(.a(G724), .O(gate246inter7));
  inv1  gate2011(.a(G736), .O(gate246inter8));
  nand2 gate2012(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate2013(.a(s_209), .b(gate246inter3), .O(gate246inter10));
  nor2  gate2014(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate2015(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate2016(.a(gate246inter12), .b(gate246inter1), .O(G759));
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate2017(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate2018(.a(gate248inter0), .b(s_210), .O(gate248inter1));
  and2  gate2019(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate2020(.a(s_210), .O(gate248inter3));
  inv1  gate2021(.a(s_211), .O(gate248inter4));
  nand2 gate2022(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate2023(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate2024(.a(G727), .O(gate248inter7));
  inv1  gate2025(.a(G739), .O(gate248inter8));
  nand2 gate2026(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate2027(.a(s_211), .b(gate248inter3), .O(gate248inter10));
  nor2  gate2028(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate2029(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate2030(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate1905(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate1906(.a(gate250inter0), .b(s_194), .O(gate250inter1));
  and2  gate1907(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate1908(.a(s_194), .O(gate250inter3));
  inv1  gate1909(.a(s_195), .O(gate250inter4));
  nand2 gate1910(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate1911(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate1912(.a(G706), .O(gate250inter7));
  inv1  gate1913(.a(G742), .O(gate250inter8));
  nand2 gate1914(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate1915(.a(s_195), .b(gate250inter3), .O(gate250inter10));
  nor2  gate1916(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate1917(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate1918(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate2143(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate2144(.a(gate253inter0), .b(s_228), .O(gate253inter1));
  and2  gate2145(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate2146(.a(s_228), .O(gate253inter3));
  inv1  gate2147(.a(s_229), .O(gate253inter4));
  nand2 gate2148(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate2149(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate2150(.a(G260), .O(gate253inter7));
  inv1  gate2151(.a(G748), .O(gate253inter8));
  nand2 gate2152(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate2153(.a(s_229), .b(gate253inter3), .O(gate253inter10));
  nor2  gate2154(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate2155(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate2156(.a(gate253inter12), .b(gate253inter1), .O(G766));

  xor2  gate1807(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate1808(.a(gate254inter0), .b(s_180), .O(gate254inter1));
  and2  gate1809(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate1810(.a(s_180), .O(gate254inter3));
  inv1  gate1811(.a(s_181), .O(gate254inter4));
  nand2 gate1812(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate1813(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate1814(.a(G712), .O(gate254inter7));
  inv1  gate1815(.a(G748), .O(gate254inter8));
  nand2 gate1816(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate1817(.a(s_181), .b(gate254inter3), .O(gate254inter10));
  nor2  gate1818(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate1819(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate1820(.a(gate254inter12), .b(gate254inter1), .O(G767));

  xor2  gate1303(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate1304(.a(gate255inter0), .b(s_108), .O(gate255inter1));
  and2  gate1305(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate1306(.a(s_108), .O(gate255inter3));
  inv1  gate1307(.a(s_109), .O(gate255inter4));
  nand2 gate1308(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate1309(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate1310(.a(G263), .O(gate255inter7));
  inv1  gate1311(.a(G751), .O(gate255inter8));
  nand2 gate1312(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate1313(.a(s_109), .b(gate255inter3), .O(gate255inter10));
  nor2  gate1314(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate1315(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate1316(.a(gate255inter12), .b(gate255inter1), .O(G768));
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate2031(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate2032(.a(gate262inter0), .b(s_212), .O(gate262inter1));
  and2  gate2033(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate2034(.a(s_212), .O(gate262inter3));
  inv1  gate2035(.a(s_213), .O(gate262inter4));
  nand2 gate2036(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate2037(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate2038(.a(G764), .O(gate262inter7));
  inv1  gate2039(.a(G765), .O(gate262inter8));
  nand2 gate2040(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate2041(.a(s_213), .b(gate262inter3), .O(gate262inter10));
  nor2  gate2042(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate2043(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate2044(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate1793(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate1794(.a(gate265inter0), .b(s_178), .O(gate265inter1));
  and2  gate1795(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate1796(.a(s_178), .O(gate265inter3));
  inv1  gate1797(.a(s_179), .O(gate265inter4));
  nand2 gate1798(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate1799(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate1800(.a(G642), .O(gate265inter7));
  inv1  gate1801(.a(G770), .O(gate265inter8));
  nand2 gate1802(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate1803(.a(s_179), .b(gate265inter3), .O(gate265inter10));
  nor2  gate1804(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate1805(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate1806(.a(gate265inter12), .b(gate265inter1), .O(G794));

  xor2  gate981(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate982(.a(gate266inter0), .b(s_62), .O(gate266inter1));
  and2  gate983(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate984(.a(s_62), .O(gate266inter3));
  inv1  gate985(.a(s_63), .O(gate266inter4));
  nand2 gate986(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate987(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate988(.a(G645), .O(gate266inter7));
  inv1  gate989(.a(G773), .O(gate266inter8));
  nand2 gate990(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate991(.a(s_63), .b(gate266inter3), .O(gate266inter10));
  nor2  gate992(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate993(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate994(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate1695(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate1696(.a(gate268inter0), .b(s_164), .O(gate268inter1));
  and2  gate1697(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate1698(.a(s_164), .O(gate268inter3));
  inv1  gate1699(.a(s_165), .O(gate268inter4));
  nand2 gate1700(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1701(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1702(.a(G651), .O(gate268inter7));
  inv1  gate1703(.a(G779), .O(gate268inter8));
  nand2 gate1704(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1705(.a(s_165), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1706(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1707(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1708(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate1415(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate1416(.a(gate270inter0), .b(s_124), .O(gate270inter1));
  and2  gate1417(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate1418(.a(s_124), .O(gate270inter3));
  inv1  gate1419(.a(s_125), .O(gate270inter4));
  nand2 gate1420(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate1421(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate1422(.a(G657), .O(gate270inter7));
  inv1  gate1423(.a(G785), .O(gate270inter8));
  nand2 gate1424(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate1425(.a(s_125), .b(gate270inter3), .O(gate270inter10));
  nor2  gate1426(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate1427(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate1428(.a(gate270inter12), .b(gate270inter1), .O(G809));

  xor2  gate1541(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate1542(.a(gate271inter0), .b(s_142), .O(gate271inter1));
  and2  gate1543(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate1544(.a(s_142), .O(gate271inter3));
  inv1  gate1545(.a(s_143), .O(gate271inter4));
  nand2 gate1546(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate1547(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate1548(.a(G660), .O(gate271inter7));
  inv1  gate1549(.a(G788), .O(gate271inter8));
  nand2 gate1550(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate1551(.a(s_143), .b(gate271inter3), .O(gate271inter10));
  nor2  gate1552(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate1553(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate1554(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate1345(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate1346(.a(gate276inter0), .b(s_114), .O(gate276inter1));
  and2  gate1347(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate1348(.a(s_114), .O(gate276inter3));
  inv1  gate1349(.a(s_115), .O(gate276inter4));
  nand2 gate1350(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate1351(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate1352(.a(G773), .O(gate276inter7));
  inv1  gate1353(.a(G797), .O(gate276inter8));
  nand2 gate1354(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate1355(.a(s_115), .b(gate276inter3), .O(gate276inter10));
  nor2  gate1356(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate1357(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate1358(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate575(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate576(.a(gate279inter0), .b(s_4), .O(gate279inter1));
  and2  gate577(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate578(.a(s_4), .O(gate279inter3));
  inv1  gate579(.a(s_5), .O(gate279inter4));
  nand2 gate580(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate581(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate582(.a(G651), .O(gate279inter7));
  inv1  gate583(.a(G803), .O(gate279inter8));
  nand2 gate584(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate585(.a(s_5), .b(gate279inter3), .O(gate279inter10));
  nor2  gate586(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate587(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate588(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );

  xor2  gate1177(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate1178(.a(gate281inter0), .b(s_90), .O(gate281inter1));
  and2  gate1179(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate1180(.a(s_90), .O(gate281inter3));
  inv1  gate1181(.a(s_91), .O(gate281inter4));
  nand2 gate1182(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate1183(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate1184(.a(G654), .O(gate281inter7));
  inv1  gate1185(.a(G806), .O(gate281inter8));
  nand2 gate1186(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate1187(.a(s_91), .b(gate281inter3), .O(gate281inter10));
  nor2  gate1188(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate1189(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate1190(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate1023(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate1024(.a(gate287inter0), .b(s_68), .O(gate287inter1));
  and2  gate1025(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate1026(.a(s_68), .O(gate287inter3));
  inv1  gate1027(.a(s_69), .O(gate287inter4));
  nand2 gate1028(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate1029(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate1030(.a(G663), .O(gate287inter7));
  inv1  gate1031(.a(G815), .O(gate287inter8));
  nand2 gate1032(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate1033(.a(s_69), .b(gate287inter3), .O(gate287inter10));
  nor2  gate1034(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate1035(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate1036(.a(gate287inter12), .b(gate287inter1), .O(G832));

  xor2  gate1611(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate1612(.a(gate288inter0), .b(s_152), .O(gate288inter1));
  and2  gate1613(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate1614(.a(s_152), .O(gate288inter3));
  inv1  gate1615(.a(s_153), .O(gate288inter4));
  nand2 gate1616(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate1617(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate1618(.a(G791), .O(gate288inter7));
  inv1  gate1619(.a(G815), .O(gate288inter8));
  nand2 gate1620(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate1621(.a(s_153), .b(gate288inter3), .O(gate288inter10));
  nor2  gate1622(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate1623(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate1624(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate813(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate814(.a(gate290inter0), .b(s_38), .O(gate290inter1));
  and2  gate815(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate816(.a(s_38), .O(gate290inter3));
  inv1  gate817(.a(s_39), .O(gate290inter4));
  nand2 gate818(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate819(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate820(.a(G820), .O(gate290inter7));
  inv1  gate821(.a(G821), .O(gate290inter8));
  nand2 gate822(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate823(.a(s_39), .b(gate290inter3), .O(gate290inter10));
  nor2  gate824(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate825(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate826(.a(gate290inter12), .b(gate290inter1), .O(G847));

  xor2  gate645(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate646(.a(gate291inter0), .b(s_14), .O(gate291inter1));
  and2  gate647(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate648(.a(s_14), .O(gate291inter3));
  inv1  gate649(.a(s_15), .O(gate291inter4));
  nand2 gate650(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate651(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate652(.a(G822), .O(gate291inter7));
  inv1  gate653(.a(G823), .O(gate291inter8));
  nand2 gate654(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate655(.a(s_15), .b(gate291inter3), .O(gate291inter10));
  nor2  gate656(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate657(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate658(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate1247(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate1248(.a(gate296inter0), .b(s_100), .O(gate296inter1));
  and2  gate1249(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate1250(.a(s_100), .O(gate296inter3));
  inv1  gate1251(.a(s_101), .O(gate296inter4));
  nand2 gate1252(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate1253(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate1254(.a(G826), .O(gate296inter7));
  inv1  gate1255(.a(G827), .O(gate296inter8));
  nand2 gate1256(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate1257(.a(s_101), .b(gate296inter3), .O(gate296inter10));
  nor2  gate1258(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate1259(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate1260(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate2045(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate2046(.a(gate388inter0), .b(s_214), .O(gate388inter1));
  and2  gate2047(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate2048(.a(s_214), .O(gate388inter3));
  inv1  gate2049(.a(s_215), .O(gate388inter4));
  nand2 gate2050(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate2051(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate2052(.a(G2), .O(gate388inter7));
  inv1  gate2053(.a(G1039), .O(gate388inter8));
  nand2 gate2054(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate2055(.a(s_215), .b(gate388inter3), .O(gate388inter10));
  nor2  gate2056(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate2057(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate2058(.a(gate388inter12), .b(gate388inter1), .O(G1135));

  xor2  gate729(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate730(.a(gate389inter0), .b(s_26), .O(gate389inter1));
  and2  gate731(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate732(.a(s_26), .O(gate389inter3));
  inv1  gate733(.a(s_27), .O(gate389inter4));
  nand2 gate734(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate735(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate736(.a(G3), .O(gate389inter7));
  inv1  gate737(.a(G1042), .O(gate389inter8));
  nand2 gate738(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate739(.a(s_27), .b(gate389inter3), .O(gate389inter10));
  nor2  gate740(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate741(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate742(.a(gate389inter12), .b(gate389inter1), .O(G1138));

  xor2  gate1079(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate1080(.a(gate390inter0), .b(s_76), .O(gate390inter1));
  and2  gate1081(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate1082(.a(s_76), .O(gate390inter3));
  inv1  gate1083(.a(s_77), .O(gate390inter4));
  nand2 gate1084(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate1085(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate1086(.a(G4), .O(gate390inter7));
  inv1  gate1087(.a(G1045), .O(gate390inter8));
  nand2 gate1088(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate1089(.a(s_77), .b(gate390inter3), .O(gate390inter10));
  nor2  gate1090(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate1091(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate1092(.a(gate390inter12), .b(gate390inter1), .O(G1141));

  xor2  gate1513(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate1514(.a(gate391inter0), .b(s_138), .O(gate391inter1));
  and2  gate1515(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate1516(.a(s_138), .O(gate391inter3));
  inv1  gate1517(.a(s_139), .O(gate391inter4));
  nand2 gate1518(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate1519(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate1520(.a(G5), .O(gate391inter7));
  inv1  gate1521(.a(G1048), .O(gate391inter8));
  nand2 gate1522(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate1523(.a(s_139), .b(gate391inter3), .O(gate391inter10));
  nor2  gate1524(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate1525(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate1526(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate1961(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate1962(.a(gate394inter0), .b(s_202), .O(gate394inter1));
  and2  gate1963(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate1964(.a(s_202), .O(gate394inter3));
  inv1  gate1965(.a(s_203), .O(gate394inter4));
  nand2 gate1966(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate1967(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate1968(.a(G8), .O(gate394inter7));
  inv1  gate1969(.a(G1057), .O(gate394inter8));
  nand2 gate1970(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate1971(.a(s_203), .b(gate394inter3), .O(gate394inter10));
  nor2  gate1972(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate1973(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate1974(.a(gate394inter12), .b(gate394inter1), .O(G1153));

  xor2  gate1093(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1094(.a(gate395inter0), .b(s_78), .O(gate395inter1));
  and2  gate1095(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1096(.a(s_78), .O(gate395inter3));
  inv1  gate1097(.a(s_79), .O(gate395inter4));
  nand2 gate1098(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1099(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1100(.a(G9), .O(gate395inter7));
  inv1  gate1101(.a(G1060), .O(gate395inter8));
  nand2 gate1102(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1103(.a(s_79), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1104(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1105(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1106(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate911(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate912(.a(gate400inter0), .b(s_52), .O(gate400inter1));
  and2  gate913(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate914(.a(s_52), .O(gate400inter3));
  inv1  gate915(.a(s_53), .O(gate400inter4));
  nand2 gate916(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate917(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate918(.a(G14), .O(gate400inter7));
  inv1  gate919(.a(G1075), .O(gate400inter8));
  nand2 gate920(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate921(.a(s_53), .b(gate400inter3), .O(gate400inter10));
  nor2  gate922(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate923(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate924(.a(gate400inter12), .b(gate400inter1), .O(G1171));

  xor2  gate2311(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate2312(.a(gate401inter0), .b(s_252), .O(gate401inter1));
  and2  gate2313(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate2314(.a(s_252), .O(gate401inter3));
  inv1  gate2315(.a(s_253), .O(gate401inter4));
  nand2 gate2316(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate2317(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate2318(.a(G15), .O(gate401inter7));
  inv1  gate2319(.a(G1078), .O(gate401inter8));
  nand2 gate2320(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate2321(.a(s_253), .b(gate401inter3), .O(gate401inter10));
  nor2  gate2322(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate2323(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate2324(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate1863(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate1864(.a(gate410inter0), .b(s_188), .O(gate410inter1));
  and2  gate1865(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate1866(.a(s_188), .O(gate410inter3));
  inv1  gate1867(.a(s_189), .O(gate410inter4));
  nand2 gate1868(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate1869(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate1870(.a(G24), .O(gate410inter7));
  inv1  gate1871(.a(G1105), .O(gate410inter8));
  nand2 gate1872(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate1873(.a(s_189), .b(gate410inter3), .O(gate410inter10));
  nor2  gate1874(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate1875(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate1876(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate2339(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate2340(.a(gate413inter0), .b(s_256), .O(gate413inter1));
  and2  gate2341(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate2342(.a(s_256), .O(gate413inter3));
  inv1  gate2343(.a(s_257), .O(gate413inter4));
  nand2 gate2344(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate2345(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate2346(.a(G27), .O(gate413inter7));
  inv1  gate2347(.a(G1114), .O(gate413inter8));
  nand2 gate2348(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate2349(.a(s_257), .b(gate413inter3), .O(gate413inter10));
  nor2  gate2350(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate2351(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate2352(.a(gate413inter12), .b(gate413inter1), .O(G1210));

  xor2  gate2325(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate2326(.a(gate414inter0), .b(s_254), .O(gate414inter1));
  and2  gate2327(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate2328(.a(s_254), .O(gate414inter3));
  inv1  gate2329(.a(s_255), .O(gate414inter4));
  nand2 gate2330(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate2331(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate2332(.a(G28), .O(gate414inter7));
  inv1  gate2333(.a(G1117), .O(gate414inter8));
  nand2 gate2334(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate2335(.a(s_255), .b(gate414inter3), .O(gate414inter10));
  nor2  gate2336(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate2337(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate2338(.a(gate414inter12), .b(gate414inter1), .O(G1213));

  xor2  gate1555(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate1556(.a(gate415inter0), .b(s_144), .O(gate415inter1));
  and2  gate1557(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate1558(.a(s_144), .O(gate415inter3));
  inv1  gate1559(.a(s_145), .O(gate415inter4));
  nand2 gate1560(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate1561(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate1562(.a(G29), .O(gate415inter7));
  inv1  gate1563(.a(G1120), .O(gate415inter8));
  nand2 gate1564(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate1565(.a(s_145), .b(gate415inter3), .O(gate415inter10));
  nor2  gate1566(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate1567(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate1568(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate1527(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1528(.a(gate420inter0), .b(s_140), .O(gate420inter1));
  and2  gate1529(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1530(.a(s_140), .O(gate420inter3));
  inv1  gate1531(.a(s_141), .O(gate420inter4));
  nand2 gate1532(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1533(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1534(.a(G1036), .O(gate420inter7));
  inv1  gate1535(.a(G1132), .O(gate420inter8));
  nand2 gate1536(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1537(.a(s_141), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1538(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1539(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1540(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate1933(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate1934(.a(gate422inter0), .b(s_198), .O(gate422inter1));
  and2  gate1935(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate1936(.a(s_198), .O(gate422inter3));
  inv1  gate1937(.a(s_199), .O(gate422inter4));
  nand2 gate1938(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate1939(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate1940(.a(G1039), .O(gate422inter7));
  inv1  gate1941(.a(G1135), .O(gate422inter8));
  nand2 gate1942(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate1943(.a(s_199), .b(gate422inter3), .O(gate422inter10));
  nor2  gate1944(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate1945(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate1946(.a(gate422inter12), .b(gate422inter1), .O(G1231));

  xor2  gate967(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate968(.a(gate423inter0), .b(s_60), .O(gate423inter1));
  and2  gate969(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate970(.a(s_60), .O(gate423inter3));
  inv1  gate971(.a(s_61), .O(gate423inter4));
  nand2 gate972(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate973(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate974(.a(G3), .O(gate423inter7));
  inv1  gate975(.a(G1138), .O(gate423inter8));
  nand2 gate976(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate977(.a(s_61), .b(gate423inter3), .O(gate423inter10));
  nor2  gate978(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate979(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate980(.a(gate423inter12), .b(gate423inter1), .O(G1232));

  xor2  gate1485(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate1486(.a(gate424inter0), .b(s_134), .O(gate424inter1));
  and2  gate1487(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate1488(.a(s_134), .O(gate424inter3));
  inv1  gate1489(.a(s_135), .O(gate424inter4));
  nand2 gate1490(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate1491(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate1492(.a(G1042), .O(gate424inter7));
  inv1  gate1493(.a(G1138), .O(gate424inter8));
  nand2 gate1494(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate1495(.a(s_135), .b(gate424inter3), .O(gate424inter10));
  nor2  gate1496(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate1497(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate1498(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );

  xor2  gate2283(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate2284(.a(gate426inter0), .b(s_248), .O(gate426inter1));
  and2  gate2285(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate2286(.a(s_248), .O(gate426inter3));
  inv1  gate2287(.a(s_249), .O(gate426inter4));
  nand2 gate2288(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate2289(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate2290(.a(G1045), .O(gate426inter7));
  inv1  gate2291(.a(G1141), .O(gate426inter8));
  nand2 gate2292(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate2293(.a(s_249), .b(gate426inter3), .O(gate426inter10));
  nor2  gate2294(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate2295(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate2296(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate1499(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate1500(.a(gate434inter0), .b(s_136), .O(gate434inter1));
  and2  gate1501(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate1502(.a(s_136), .O(gate434inter3));
  inv1  gate1503(.a(s_137), .O(gate434inter4));
  nand2 gate1504(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate1505(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate1506(.a(G1057), .O(gate434inter7));
  inv1  gate1507(.a(G1153), .O(gate434inter8));
  nand2 gate1508(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate1509(.a(s_137), .b(gate434inter3), .O(gate434inter10));
  nor2  gate1510(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate1511(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate1512(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate1289(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate1290(.a(gate438inter0), .b(s_106), .O(gate438inter1));
  and2  gate1291(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate1292(.a(s_106), .O(gate438inter3));
  inv1  gate1293(.a(s_107), .O(gate438inter4));
  nand2 gate1294(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate1295(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate1296(.a(G1063), .O(gate438inter7));
  inv1  gate1297(.a(G1159), .O(gate438inter8));
  nand2 gate1298(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate1299(.a(s_107), .b(gate438inter3), .O(gate438inter10));
  nor2  gate1300(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate1301(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate1302(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate1681(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate1682(.a(gate443inter0), .b(s_162), .O(gate443inter1));
  and2  gate1683(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate1684(.a(s_162), .O(gate443inter3));
  inv1  gate1685(.a(s_163), .O(gate443inter4));
  nand2 gate1686(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate1687(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate1688(.a(G13), .O(gate443inter7));
  inv1  gate1689(.a(G1168), .O(gate443inter8));
  nand2 gate1690(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate1691(.a(s_163), .b(gate443inter3), .O(gate443inter10));
  nor2  gate1692(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate1693(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate1694(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );

  xor2  gate1331(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate1332(.a(gate447inter0), .b(s_112), .O(gate447inter1));
  and2  gate1333(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate1334(.a(s_112), .O(gate447inter3));
  inv1  gate1335(.a(s_113), .O(gate447inter4));
  nand2 gate1336(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate1337(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate1338(.a(G15), .O(gate447inter7));
  inv1  gate1339(.a(G1174), .O(gate447inter8));
  nand2 gate1340(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate1341(.a(s_113), .b(gate447inter3), .O(gate447inter10));
  nor2  gate1342(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate1343(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate1344(.a(gate447inter12), .b(gate447inter1), .O(G1256));
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );

  xor2  gate1261(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate1262(.a(gate450inter0), .b(s_102), .O(gate450inter1));
  and2  gate1263(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate1264(.a(s_102), .O(gate450inter3));
  inv1  gate1265(.a(s_103), .O(gate450inter4));
  nand2 gate1266(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate1267(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate1268(.a(G1081), .O(gate450inter7));
  inv1  gate1269(.a(G1177), .O(gate450inter8));
  nand2 gate1270(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate1271(.a(s_103), .b(gate450inter3), .O(gate450inter10));
  nor2  gate1272(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate1273(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate1274(.a(gate450inter12), .b(gate450inter1), .O(G1259));

  xor2  gate617(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate618(.a(gate451inter0), .b(s_10), .O(gate451inter1));
  and2  gate619(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate620(.a(s_10), .O(gate451inter3));
  inv1  gate621(.a(s_11), .O(gate451inter4));
  nand2 gate622(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate623(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate624(.a(G17), .O(gate451inter7));
  inv1  gate625(.a(G1180), .O(gate451inter8));
  nand2 gate626(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate627(.a(s_11), .b(gate451inter3), .O(gate451inter10));
  nor2  gate628(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate629(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate630(.a(gate451inter12), .b(gate451inter1), .O(G1260));

  xor2  gate1149(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate1150(.a(gate452inter0), .b(s_86), .O(gate452inter1));
  and2  gate1151(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate1152(.a(s_86), .O(gate452inter3));
  inv1  gate1153(.a(s_87), .O(gate452inter4));
  nand2 gate1154(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate1155(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate1156(.a(G1084), .O(gate452inter7));
  inv1  gate1157(.a(G1180), .O(gate452inter8));
  nand2 gate1158(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate1159(.a(s_87), .b(gate452inter3), .O(gate452inter10));
  nor2  gate1160(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate1161(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate1162(.a(gate452inter12), .b(gate452inter1), .O(G1261));

  xor2  gate631(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate632(.a(gate453inter0), .b(s_12), .O(gate453inter1));
  and2  gate633(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate634(.a(s_12), .O(gate453inter3));
  inv1  gate635(.a(s_13), .O(gate453inter4));
  nand2 gate636(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate637(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate638(.a(G18), .O(gate453inter7));
  inv1  gate639(.a(G1183), .O(gate453inter8));
  nand2 gate640(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate641(.a(s_13), .b(gate453inter3), .O(gate453inter10));
  nor2  gate642(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate643(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate644(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate561(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate562(.a(gate457inter0), .b(s_2), .O(gate457inter1));
  and2  gate563(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate564(.a(s_2), .O(gate457inter3));
  inv1  gate565(.a(s_3), .O(gate457inter4));
  nand2 gate566(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate567(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate568(.a(G20), .O(gate457inter7));
  inv1  gate569(.a(G1189), .O(gate457inter8));
  nand2 gate570(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate571(.a(s_3), .b(gate457inter3), .O(gate457inter10));
  nor2  gate572(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate573(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate574(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate1107(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate1108(.a(gate463inter0), .b(s_80), .O(gate463inter1));
  and2  gate1109(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate1110(.a(s_80), .O(gate463inter3));
  inv1  gate1111(.a(s_81), .O(gate463inter4));
  nand2 gate1112(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate1113(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate1114(.a(G23), .O(gate463inter7));
  inv1  gate1115(.a(G1198), .O(gate463inter8));
  nand2 gate1116(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate1117(.a(s_81), .b(gate463inter3), .O(gate463inter10));
  nor2  gate1118(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate1119(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate1120(.a(gate463inter12), .b(gate463inter1), .O(G1272));

  xor2  gate2185(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate2186(.a(gate464inter0), .b(s_234), .O(gate464inter1));
  and2  gate2187(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate2188(.a(s_234), .O(gate464inter3));
  inv1  gate2189(.a(s_235), .O(gate464inter4));
  nand2 gate2190(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate2191(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate2192(.a(G1102), .O(gate464inter7));
  inv1  gate2193(.a(G1198), .O(gate464inter8));
  nand2 gate2194(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate2195(.a(s_235), .b(gate464inter3), .O(gate464inter10));
  nor2  gate2196(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate2197(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate2198(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );

  xor2  gate1667(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate1668(.a(gate468inter0), .b(s_160), .O(gate468inter1));
  and2  gate1669(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate1670(.a(s_160), .O(gate468inter3));
  inv1  gate1671(.a(s_161), .O(gate468inter4));
  nand2 gate1672(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate1673(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate1674(.a(G1108), .O(gate468inter7));
  inv1  gate1675(.a(G1204), .O(gate468inter8));
  nand2 gate1676(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate1677(.a(s_161), .b(gate468inter3), .O(gate468inter10));
  nor2  gate1678(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate1679(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate1680(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate2353(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate2354(.a(gate474inter0), .b(s_258), .O(gate474inter1));
  and2  gate2355(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate2356(.a(s_258), .O(gate474inter3));
  inv1  gate2357(.a(s_259), .O(gate474inter4));
  nand2 gate2358(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate2359(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate2360(.a(G1117), .O(gate474inter7));
  inv1  gate2361(.a(G1213), .O(gate474inter8));
  nand2 gate2362(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate2363(.a(s_259), .b(gate474inter3), .O(gate474inter10));
  nor2  gate2364(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate2365(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate2366(.a(gate474inter12), .b(gate474inter1), .O(G1283));

  xor2  gate2297(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate2298(.a(gate475inter0), .b(s_250), .O(gate475inter1));
  and2  gate2299(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate2300(.a(s_250), .O(gate475inter3));
  inv1  gate2301(.a(s_251), .O(gate475inter4));
  nand2 gate2302(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate2303(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate2304(.a(G29), .O(gate475inter7));
  inv1  gate2305(.a(G1216), .O(gate475inter8));
  nand2 gate2306(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate2307(.a(s_251), .b(gate475inter3), .O(gate475inter10));
  nor2  gate2308(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate2309(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate2310(.a(gate475inter12), .b(gate475inter1), .O(G1284));
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );

  xor2  gate2227(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate2228(.a(gate478inter0), .b(s_240), .O(gate478inter1));
  and2  gate2229(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate2230(.a(s_240), .O(gate478inter3));
  inv1  gate2231(.a(s_241), .O(gate478inter4));
  nand2 gate2232(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate2233(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate2234(.a(G1123), .O(gate478inter7));
  inv1  gate2235(.a(G1219), .O(gate478inter8));
  nand2 gate2236(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate2237(.a(s_241), .b(gate478inter3), .O(gate478inter10));
  nor2  gate2238(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate2239(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate2240(.a(gate478inter12), .b(gate478inter1), .O(G1287));

  xor2  gate1723(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate1724(.a(gate479inter0), .b(s_168), .O(gate479inter1));
  and2  gate1725(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate1726(.a(s_168), .O(gate479inter3));
  inv1  gate1727(.a(s_169), .O(gate479inter4));
  nand2 gate1728(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate1729(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate1730(.a(G31), .O(gate479inter7));
  inv1  gate1731(.a(G1222), .O(gate479inter8));
  nand2 gate1732(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate1733(.a(s_169), .b(gate479inter3), .O(gate479inter10));
  nor2  gate1734(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate1735(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate1736(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate2115(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate2116(.a(gate488inter0), .b(s_224), .O(gate488inter1));
  and2  gate2117(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate2118(.a(s_224), .O(gate488inter3));
  inv1  gate2119(.a(s_225), .O(gate488inter4));
  nand2 gate2120(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate2121(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate2122(.a(G1238), .O(gate488inter7));
  inv1  gate2123(.a(G1239), .O(gate488inter8));
  nand2 gate2124(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate2125(.a(s_225), .b(gate488inter3), .O(gate488inter10));
  nor2  gate2126(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate2127(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate2128(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate799(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate800(.a(gate492inter0), .b(s_36), .O(gate492inter1));
  and2  gate801(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate802(.a(s_36), .O(gate492inter3));
  inv1  gate803(.a(s_37), .O(gate492inter4));
  nand2 gate804(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate805(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate806(.a(G1246), .O(gate492inter7));
  inv1  gate807(.a(G1247), .O(gate492inter8));
  nand2 gate808(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate809(.a(s_37), .b(gate492inter3), .O(gate492inter10));
  nor2  gate810(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate811(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate812(.a(gate492inter12), .b(gate492inter1), .O(G1301));
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate701(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate702(.a(gate497inter0), .b(s_22), .O(gate497inter1));
  and2  gate703(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate704(.a(s_22), .O(gate497inter3));
  inv1  gate705(.a(s_23), .O(gate497inter4));
  nand2 gate706(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate707(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate708(.a(G1256), .O(gate497inter7));
  inv1  gate709(.a(G1257), .O(gate497inter8));
  nand2 gate710(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate711(.a(s_23), .b(gate497inter3), .O(gate497inter10));
  nor2  gate712(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate713(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate714(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate1583(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate1584(.a(gate500inter0), .b(s_148), .O(gate500inter1));
  and2  gate1585(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate1586(.a(s_148), .O(gate500inter3));
  inv1  gate1587(.a(s_149), .O(gate500inter4));
  nand2 gate1588(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate1589(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate1590(.a(G1262), .O(gate500inter7));
  inv1  gate1591(.a(G1263), .O(gate500inter8));
  nand2 gate1592(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate1593(.a(s_149), .b(gate500inter3), .O(gate500inter10));
  nor2  gate1594(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate1595(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate1596(.a(gate500inter12), .b(gate500inter1), .O(G1309));
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate1975(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate1976(.a(gate504inter0), .b(s_204), .O(gate504inter1));
  and2  gate1977(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate1978(.a(s_204), .O(gate504inter3));
  inv1  gate1979(.a(s_205), .O(gate504inter4));
  nand2 gate1980(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate1981(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate1982(.a(G1270), .O(gate504inter7));
  inv1  gate1983(.a(G1271), .O(gate504inter8));
  nand2 gate1984(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate1985(.a(s_205), .b(gate504inter3), .O(gate504inter10));
  nor2  gate1986(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate1987(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate1988(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate2073(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate2074(.a(gate511inter0), .b(s_218), .O(gate511inter1));
  and2  gate2075(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate2076(.a(s_218), .O(gate511inter3));
  inv1  gate2077(.a(s_219), .O(gate511inter4));
  nand2 gate2078(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate2079(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate2080(.a(G1284), .O(gate511inter7));
  inv1  gate2081(.a(G1285), .O(gate511inter8));
  nand2 gate2082(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate2083(.a(s_219), .b(gate511inter3), .O(gate511inter10));
  nor2  gate2084(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate2085(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate2086(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule