module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate1079(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate1080(.a(gate11inter0), .b(s_76), .O(gate11inter1));
  and2  gate1081(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate1082(.a(s_76), .O(gate11inter3));
  inv1  gate1083(.a(s_77), .O(gate11inter4));
  nand2 gate1084(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate1085(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate1086(.a(G5), .O(gate11inter7));
  inv1  gate1087(.a(G6), .O(gate11inter8));
  nand2 gate1088(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate1089(.a(s_77), .b(gate11inter3), .O(gate11inter10));
  nor2  gate1090(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate1091(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate1092(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate617(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate618(.a(gate18inter0), .b(s_10), .O(gate18inter1));
  and2  gate619(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate620(.a(s_10), .O(gate18inter3));
  inv1  gate621(.a(s_11), .O(gate18inter4));
  nand2 gate622(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate623(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate624(.a(G19), .O(gate18inter7));
  inv1  gate625(.a(G20), .O(gate18inter8));
  nand2 gate626(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate627(.a(s_11), .b(gate18inter3), .O(gate18inter10));
  nor2  gate628(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate629(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate630(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate967(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate968(.a(gate21inter0), .b(s_60), .O(gate21inter1));
  and2  gate969(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate970(.a(s_60), .O(gate21inter3));
  inv1  gate971(.a(s_61), .O(gate21inter4));
  nand2 gate972(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate973(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate974(.a(G25), .O(gate21inter7));
  inv1  gate975(.a(G26), .O(gate21inter8));
  nand2 gate976(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate977(.a(s_61), .b(gate21inter3), .O(gate21inter10));
  nor2  gate978(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate979(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate980(.a(gate21inter12), .b(gate21inter1), .O(G302));
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate687(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate688(.a(gate23inter0), .b(s_20), .O(gate23inter1));
  and2  gate689(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate690(.a(s_20), .O(gate23inter3));
  inv1  gate691(.a(s_21), .O(gate23inter4));
  nand2 gate692(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate693(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate694(.a(G29), .O(gate23inter7));
  inv1  gate695(.a(G30), .O(gate23inter8));
  nand2 gate696(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate697(.a(s_21), .b(gate23inter3), .O(gate23inter10));
  nor2  gate698(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate699(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate700(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate575(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate576(.a(gate29inter0), .b(s_4), .O(gate29inter1));
  and2  gate577(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate578(.a(s_4), .O(gate29inter3));
  inv1  gate579(.a(s_5), .O(gate29inter4));
  nand2 gate580(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate581(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate582(.a(G3), .O(gate29inter7));
  inv1  gate583(.a(G7), .O(gate29inter8));
  nand2 gate584(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate585(.a(s_5), .b(gate29inter3), .O(gate29inter10));
  nor2  gate586(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate587(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate588(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate715(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate716(.a(gate33inter0), .b(s_24), .O(gate33inter1));
  and2  gate717(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate718(.a(s_24), .O(gate33inter3));
  inv1  gate719(.a(s_25), .O(gate33inter4));
  nand2 gate720(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate721(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate722(.a(G17), .O(gate33inter7));
  inv1  gate723(.a(G21), .O(gate33inter8));
  nand2 gate724(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate725(.a(s_25), .b(gate33inter3), .O(gate33inter10));
  nor2  gate726(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate727(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate728(.a(gate33inter12), .b(gate33inter1), .O(G338));
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate673(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate674(.a(gate51inter0), .b(s_18), .O(gate51inter1));
  and2  gate675(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate676(.a(s_18), .O(gate51inter3));
  inv1  gate677(.a(s_19), .O(gate51inter4));
  nand2 gate678(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate679(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate680(.a(G11), .O(gate51inter7));
  inv1  gate681(.a(G281), .O(gate51inter8));
  nand2 gate682(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate683(.a(s_19), .b(gate51inter3), .O(gate51inter10));
  nor2  gate684(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate685(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate686(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate1135(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate1136(.a(gate75inter0), .b(s_84), .O(gate75inter1));
  and2  gate1137(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate1138(.a(s_84), .O(gate75inter3));
  inv1  gate1139(.a(s_85), .O(gate75inter4));
  nand2 gate1140(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate1141(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate1142(.a(G9), .O(gate75inter7));
  inv1  gate1143(.a(G317), .O(gate75inter8));
  nand2 gate1144(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate1145(.a(s_85), .b(gate75inter3), .O(gate75inter10));
  nor2  gate1146(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate1147(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate1148(.a(gate75inter12), .b(gate75inter1), .O(G396));

  xor2  gate1205(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate1206(.a(gate76inter0), .b(s_94), .O(gate76inter1));
  and2  gate1207(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate1208(.a(s_94), .O(gate76inter3));
  inv1  gate1209(.a(s_95), .O(gate76inter4));
  nand2 gate1210(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate1211(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate1212(.a(G13), .O(gate76inter7));
  inv1  gate1213(.a(G317), .O(gate76inter8));
  nand2 gate1214(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate1215(.a(s_95), .b(gate76inter3), .O(gate76inter10));
  nor2  gate1216(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate1217(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate1218(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );

  xor2  gate547(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate548(.a(gate78inter0), .b(s_0), .O(gate78inter1));
  and2  gate549(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate550(.a(s_0), .O(gate78inter3));
  inv1  gate551(.a(s_1), .O(gate78inter4));
  nand2 gate552(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate553(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate554(.a(G6), .O(gate78inter7));
  inv1  gate555(.a(G320), .O(gate78inter8));
  nand2 gate556(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate557(.a(s_1), .b(gate78inter3), .O(gate78inter10));
  nor2  gate558(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate559(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate560(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate939(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate940(.a(gate80inter0), .b(s_56), .O(gate80inter1));
  and2  gate941(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate942(.a(s_56), .O(gate80inter3));
  inv1  gate943(.a(s_57), .O(gate80inter4));
  nand2 gate944(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate945(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate946(.a(G14), .O(gate80inter7));
  inv1  gate947(.a(G323), .O(gate80inter8));
  nand2 gate948(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate949(.a(s_57), .b(gate80inter3), .O(gate80inter10));
  nor2  gate950(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate951(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate952(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate799(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate800(.a(gate86inter0), .b(s_36), .O(gate86inter1));
  and2  gate801(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate802(.a(s_36), .O(gate86inter3));
  inv1  gate803(.a(s_37), .O(gate86inter4));
  nand2 gate804(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate805(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate806(.a(G8), .O(gate86inter7));
  inv1  gate807(.a(G332), .O(gate86inter8));
  nand2 gate808(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate809(.a(s_37), .b(gate86inter3), .O(gate86inter10));
  nor2  gate810(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate811(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate812(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );

  xor2  gate1037(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate1038(.a(gate92inter0), .b(s_70), .O(gate92inter1));
  and2  gate1039(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate1040(.a(s_70), .O(gate92inter3));
  inv1  gate1041(.a(s_71), .O(gate92inter4));
  nand2 gate1042(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate1043(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate1044(.a(G29), .O(gate92inter7));
  inv1  gate1045(.a(G341), .O(gate92inter8));
  nand2 gate1046(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate1047(.a(s_71), .b(gate92inter3), .O(gate92inter10));
  nor2  gate1048(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate1049(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate1050(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate855(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate856(.a(gate104inter0), .b(s_44), .O(gate104inter1));
  and2  gate857(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate858(.a(s_44), .O(gate104inter3));
  inv1  gate859(.a(s_45), .O(gate104inter4));
  nand2 gate860(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate861(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate862(.a(G32), .O(gate104inter7));
  inv1  gate863(.a(G359), .O(gate104inter8));
  nand2 gate864(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate865(.a(s_45), .b(gate104inter3), .O(gate104inter10));
  nor2  gate866(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate867(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate868(.a(gate104inter12), .b(gate104inter1), .O(G425));

  xor2  gate561(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate562(.a(gate105inter0), .b(s_2), .O(gate105inter1));
  and2  gate563(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate564(.a(s_2), .O(gate105inter3));
  inv1  gate565(.a(s_3), .O(gate105inter4));
  nand2 gate566(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate567(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate568(.a(G362), .O(gate105inter7));
  inv1  gate569(.a(G363), .O(gate105inter8));
  nand2 gate570(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate571(.a(s_3), .b(gate105inter3), .O(gate105inter10));
  nor2  gate572(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate573(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate574(.a(gate105inter12), .b(gate105inter1), .O(G426));
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate813(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate814(.a(gate117inter0), .b(s_38), .O(gate117inter1));
  and2  gate815(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate816(.a(s_38), .O(gate117inter3));
  inv1  gate817(.a(s_39), .O(gate117inter4));
  nand2 gate818(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate819(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate820(.a(G386), .O(gate117inter7));
  inv1  gate821(.a(G387), .O(gate117inter8));
  nand2 gate822(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate823(.a(s_39), .b(gate117inter3), .O(gate117inter10));
  nor2  gate824(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate825(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate826(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );

  xor2  gate603(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate604(.a(gate139inter0), .b(s_8), .O(gate139inter1));
  and2  gate605(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate606(.a(s_8), .O(gate139inter3));
  inv1  gate607(.a(s_9), .O(gate139inter4));
  nand2 gate608(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate609(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate610(.a(G438), .O(gate139inter7));
  inv1  gate611(.a(G441), .O(gate139inter8));
  nand2 gate612(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate613(.a(s_9), .b(gate139inter3), .O(gate139inter10));
  nor2  gate614(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate615(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate616(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate645(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate646(.a(gate147inter0), .b(s_14), .O(gate147inter1));
  and2  gate647(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate648(.a(s_14), .O(gate147inter3));
  inv1  gate649(.a(s_15), .O(gate147inter4));
  nand2 gate650(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate651(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate652(.a(G486), .O(gate147inter7));
  inv1  gate653(.a(G489), .O(gate147inter8));
  nand2 gate654(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate655(.a(s_15), .b(gate147inter3), .O(gate147inter10));
  nor2  gate656(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate657(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate658(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate701(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate702(.a(gate157inter0), .b(s_22), .O(gate157inter1));
  and2  gate703(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate704(.a(s_22), .O(gate157inter3));
  inv1  gate705(.a(s_23), .O(gate157inter4));
  nand2 gate706(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate707(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate708(.a(G438), .O(gate157inter7));
  inv1  gate709(.a(G528), .O(gate157inter8));
  nand2 gate710(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate711(.a(s_23), .b(gate157inter3), .O(gate157inter10));
  nor2  gate712(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate713(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate714(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate1149(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate1150(.a(gate160inter0), .b(s_86), .O(gate160inter1));
  and2  gate1151(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate1152(.a(s_86), .O(gate160inter3));
  inv1  gate1153(.a(s_87), .O(gate160inter4));
  nand2 gate1154(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate1155(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate1156(.a(G447), .O(gate160inter7));
  inv1  gate1157(.a(G531), .O(gate160inter8));
  nand2 gate1158(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate1159(.a(s_87), .b(gate160inter3), .O(gate160inter10));
  nor2  gate1160(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate1161(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate1162(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );

  xor2  gate1233(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate1234(.a(gate163inter0), .b(s_98), .O(gate163inter1));
  and2  gate1235(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate1236(.a(s_98), .O(gate163inter3));
  inv1  gate1237(.a(s_99), .O(gate163inter4));
  nand2 gate1238(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate1239(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate1240(.a(G456), .O(gate163inter7));
  inv1  gate1241(.a(G537), .O(gate163inter8));
  nand2 gate1242(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate1243(.a(s_99), .b(gate163inter3), .O(gate163inter10));
  nor2  gate1244(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate1245(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate1246(.a(gate163inter12), .b(gate163inter1), .O(G580));
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate897(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate898(.a(gate165inter0), .b(s_50), .O(gate165inter1));
  and2  gate899(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate900(.a(s_50), .O(gate165inter3));
  inv1  gate901(.a(s_51), .O(gate165inter4));
  nand2 gate902(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate903(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate904(.a(G462), .O(gate165inter7));
  inv1  gate905(.a(G540), .O(gate165inter8));
  nand2 gate906(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate907(.a(s_51), .b(gate165inter3), .O(gate165inter10));
  nor2  gate908(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate909(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate910(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );

  xor2  gate883(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate884(.a(gate167inter0), .b(s_48), .O(gate167inter1));
  and2  gate885(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate886(.a(s_48), .O(gate167inter3));
  inv1  gate887(.a(s_49), .O(gate167inter4));
  nand2 gate888(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate889(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate890(.a(G468), .O(gate167inter7));
  inv1  gate891(.a(G543), .O(gate167inter8));
  nand2 gate892(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate893(.a(s_49), .b(gate167inter3), .O(gate167inter10));
  nor2  gate894(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate895(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate896(.a(gate167inter12), .b(gate167inter1), .O(G584));
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate953(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate954(.a(gate187inter0), .b(s_58), .O(gate187inter1));
  and2  gate955(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate956(.a(s_58), .O(gate187inter3));
  inv1  gate957(.a(s_59), .O(gate187inter4));
  nand2 gate958(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate959(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate960(.a(G574), .O(gate187inter7));
  inv1  gate961(.a(G575), .O(gate187inter8));
  nand2 gate962(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate963(.a(s_59), .b(gate187inter3), .O(gate187inter10));
  nor2  gate964(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate965(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate966(.a(gate187inter12), .b(gate187inter1), .O(G612));
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate659(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate660(.a(gate191inter0), .b(s_16), .O(gate191inter1));
  and2  gate661(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate662(.a(s_16), .O(gate191inter3));
  inv1  gate663(.a(s_17), .O(gate191inter4));
  nand2 gate664(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate665(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate666(.a(G582), .O(gate191inter7));
  inv1  gate667(.a(G583), .O(gate191inter8));
  nand2 gate668(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate669(.a(s_17), .b(gate191inter3), .O(gate191inter10));
  nor2  gate670(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate671(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate672(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );

  xor2  gate981(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate982(.a(gate199inter0), .b(s_62), .O(gate199inter1));
  and2  gate983(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate984(.a(s_62), .O(gate199inter3));
  inv1  gate985(.a(s_63), .O(gate199inter4));
  nand2 gate986(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate987(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate988(.a(G598), .O(gate199inter7));
  inv1  gate989(.a(G599), .O(gate199inter8));
  nand2 gate990(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate991(.a(s_63), .b(gate199inter3), .O(gate199inter10));
  nor2  gate992(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate993(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate994(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );

  xor2  gate743(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate744(.a(gate212inter0), .b(s_28), .O(gate212inter1));
  and2  gate745(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate746(.a(s_28), .O(gate212inter3));
  inv1  gate747(.a(s_29), .O(gate212inter4));
  nand2 gate748(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate749(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate750(.a(G617), .O(gate212inter7));
  inv1  gate751(.a(G669), .O(gate212inter8));
  nand2 gate752(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate753(.a(s_29), .b(gate212inter3), .O(gate212inter10));
  nor2  gate754(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate755(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate756(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate911(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate912(.a(gate214inter0), .b(s_52), .O(gate214inter1));
  and2  gate913(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate914(.a(s_52), .O(gate214inter3));
  inv1  gate915(.a(s_53), .O(gate214inter4));
  nand2 gate916(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate917(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate918(.a(G612), .O(gate214inter7));
  inv1  gate919(.a(G672), .O(gate214inter8));
  nand2 gate920(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate921(.a(s_53), .b(gate214inter3), .O(gate214inter10));
  nor2  gate922(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate923(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate924(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate1051(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate1052(.a(gate233inter0), .b(s_72), .O(gate233inter1));
  and2  gate1053(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate1054(.a(s_72), .O(gate233inter3));
  inv1  gate1055(.a(s_73), .O(gate233inter4));
  nand2 gate1056(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1057(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1058(.a(G242), .O(gate233inter7));
  inv1  gate1059(.a(G718), .O(gate233inter8));
  nand2 gate1060(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1061(.a(s_73), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1062(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1063(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1064(.a(gate233inter12), .b(gate233inter1), .O(G730));

  xor2  gate1107(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate1108(.a(gate234inter0), .b(s_80), .O(gate234inter1));
  and2  gate1109(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate1110(.a(s_80), .O(gate234inter3));
  inv1  gate1111(.a(s_81), .O(gate234inter4));
  nand2 gate1112(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1113(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1114(.a(G245), .O(gate234inter7));
  inv1  gate1115(.a(G721), .O(gate234inter8));
  nand2 gate1116(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1117(.a(s_81), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1118(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1119(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1120(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );

  xor2  gate1009(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate1010(.a(gate242inter0), .b(s_66), .O(gate242inter1));
  and2  gate1011(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate1012(.a(s_66), .O(gate242inter3));
  inv1  gate1013(.a(s_67), .O(gate242inter4));
  nand2 gate1014(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate1015(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate1016(.a(G718), .O(gate242inter7));
  inv1  gate1017(.a(G730), .O(gate242inter8));
  nand2 gate1018(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate1019(.a(s_67), .b(gate242inter3), .O(gate242inter10));
  nor2  gate1020(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate1021(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate1022(.a(gate242inter12), .b(gate242inter1), .O(G755));

  xor2  gate1023(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1024(.a(gate243inter0), .b(s_68), .O(gate243inter1));
  and2  gate1025(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1026(.a(s_68), .O(gate243inter3));
  inv1  gate1027(.a(s_69), .O(gate243inter4));
  nand2 gate1028(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1029(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1030(.a(G245), .O(gate243inter7));
  inv1  gate1031(.a(G733), .O(gate243inter8));
  nand2 gate1032(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1033(.a(s_69), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1034(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1035(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1036(.a(gate243inter12), .b(gate243inter1), .O(G756));

  xor2  gate785(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate786(.a(gate244inter0), .b(s_34), .O(gate244inter1));
  and2  gate787(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate788(.a(s_34), .O(gate244inter3));
  inv1  gate789(.a(s_35), .O(gate244inter4));
  nand2 gate790(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate791(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate792(.a(G721), .O(gate244inter7));
  inv1  gate793(.a(G733), .O(gate244inter8));
  nand2 gate794(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate795(.a(s_35), .b(gate244inter3), .O(gate244inter10));
  nor2  gate796(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate797(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate798(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );

  xor2  gate995(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate996(.a(gate246inter0), .b(s_64), .O(gate246inter1));
  and2  gate997(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate998(.a(s_64), .O(gate246inter3));
  inv1  gate999(.a(s_65), .O(gate246inter4));
  nand2 gate1000(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate1001(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate1002(.a(G724), .O(gate246inter7));
  inv1  gate1003(.a(G736), .O(gate246inter8));
  nand2 gate1004(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate1005(.a(s_65), .b(gate246inter3), .O(gate246inter10));
  nor2  gate1006(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate1007(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate1008(.a(gate246inter12), .b(gate246inter1), .O(G759));
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate1177(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate1178(.a(gate262inter0), .b(s_90), .O(gate262inter1));
  and2  gate1179(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate1180(.a(s_90), .O(gate262inter3));
  inv1  gate1181(.a(s_91), .O(gate262inter4));
  nand2 gate1182(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate1183(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate1184(.a(G764), .O(gate262inter7));
  inv1  gate1185(.a(G765), .O(gate262inter8));
  nand2 gate1186(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate1187(.a(s_91), .b(gate262inter3), .O(gate262inter10));
  nor2  gate1188(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate1189(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate1190(.a(gate262inter12), .b(gate262inter1), .O(G785));

  xor2  gate631(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate632(.a(gate263inter0), .b(s_12), .O(gate263inter1));
  and2  gate633(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate634(.a(s_12), .O(gate263inter3));
  inv1  gate635(.a(s_13), .O(gate263inter4));
  nand2 gate636(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate637(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate638(.a(G766), .O(gate263inter7));
  inv1  gate639(.a(G767), .O(gate263inter8));
  nand2 gate640(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate641(.a(s_13), .b(gate263inter3), .O(gate263inter10));
  nor2  gate642(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate643(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate644(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate729(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate730(.a(gate267inter0), .b(s_26), .O(gate267inter1));
  and2  gate731(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate732(.a(s_26), .O(gate267inter3));
  inv1  gate733(.a(s_27), .O(gate267inter4));
  nand2 gate734(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate735(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate736(.a(G648), .O(gate267inter7));
  inv1  gate737(.a(G776), .O(gate267inter8));
  nand2 gate738(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate739(.a(s_27), .b(gate267inter3), .O(gate267inter10));
  nor2  gate740(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate741(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate742(.a(gate267inter12), .b(gate267inter1), .O(G800));

  xor2  gate757(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate758(.a(gate268inter0), .b(s_30), .O(gate268inter1));
  and2  gate759(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate760(.a(s_30), .O(gate268inter3));
  inv1  gate761(.a(s_31), .O(gate268inter4));
  nand2 gate762(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate763(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate764(.a(G651), .O(gate268inter7));
  inv1  gate765(.a(G779), .O(gate268inter8));
  nand2 gate766(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate767(.a(s_31), .b(gate268inter3), .O(gate268inter10));
  nor2  gate768(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate769(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate770(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate589(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate590(.a(gate270inter0), .b(s_6), .O(gate270inter1));
  and2  gate591(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate592(.a(s_6), .O(gate270inter3));
  inv1  gate593(.a(s_7), .O(gate270inter4));
  nand2 gate594(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate595(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate596(.a(G657), .O(gate270inter7));
  inv1  gate597(.a(G785), .O(gate270inter8));
  nand2 gate598(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate599(.a(s_7), .b(gate270inter3), .O(gate270inter10));
  nor2  gate600(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate601(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate602(.a(gate270inter12), .b(gate270inter1), .O(G809));

  xor2  gate1163(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate1164(.a(gate271inter0), .b(s_88), .O(gate271inter1));
  and2  gate1165(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate1166(.a(s_88), .O(gate271inter3));
  inv1  gate1167(.a(s_89), .O(gate271inter4));
  nand2 gate1168(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate1169(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate1170(.a(G660), .O(gate271inter7));
  inv1  gate1171(.a(G788), .O(gate271inter8));
  nand2 gate1172(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate1173(.a(s_89), .b(gate271inter3), .O(gate271inter10));
  nor2  gate1174(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate1175(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate1176(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate1121(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate1122(.a(gate290inter0), .b(s_82), .O(gate290inter1));
  and2  gate1123(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate1124(.a(s_82), .O(gate290inter3));
  inv1  gate1125(.a(s_83), .O(gate290inter4));
  nand2 gate1126(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate1127(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate1128(.a(G820), .O(gate290inter7));
  inv1  gate1129(.a(G821), .O(gate290inter8));
  nand2 gate1130(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate1131(.a(s_83), .b(gate290inter3), .O(gate290inter10));
  nor2  gate1132(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate1133(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate1134(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate1093(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate1094(.a(gate389inter0), .b(s_78), .O(gate389inter1));
  and2  gate1095(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate1096(.a(s_78), .O(gate389inter3));
  inv1  gate1097(.a(s_79), .O(gate389inter4));
  nand2 gate1098(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate1099(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate1100(.a(G3), .O(gate389inter7));
  inv1  gate1101(.a(G1042), .O(gate389inter8));
  nand2 gate1102(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate1103(.a(s_79), .b(gate389inter3), .O(gate389inter10));
  nor2  gate1104(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate1105(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate1106(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate1191(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate1192(.a(gate417inter0), .b(s_92), .O(gate417inter1));
  and2  gate1193(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate1194(.a(s_92), .O(gate417inter3));
  inv1  gate1195(.a(s_93), .O(gate417inter4));
  nand2 gate1196(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate1197(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate1198(.a(G31), .O(gate417inter7));
  inv1  gate1199(.a(G1126), .O(gate417inter8));
  nand2 gate1200(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate1201(.a(s_93), .b(gate417inter3), .O(gate417inter10));
  nor2  gate1202(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate1203(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate1204(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate1065(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate1066(.a(gate434inter0), .b(s_74), .O(gate434inter1));
  and2  gate1067(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate1068(.a(s_74), .O(gate434inter3));
  inv1  gate1069(.a(s_75), .O(gate434inter4));
  nand2 gate1070(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate1071(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate1072(.a(G1057), .O(gate434inter7));
  inv1  gate1073(.a(G1153), .O(gate434inter8));
  nand2 gate1074(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate1075(.a(s_75), .b(gate434inter3), .O(gate434inter10));
  nor2  gate1076(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate1077(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate1078(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate771(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate772(.a(gate438inter0), .b(s_32), .O(gate438inter1));
  and2  gate773(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate774(.a(s_32), .O(gate438inter3));
  inv1  gate775(.a(s_33), .O(gate438inter4));
  nand2 gate776(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate777(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate778(.a(G1063), .O(gate438inter7));
  inv1  gate779(.a(G1159), .O(gate438inter8));
  nand2 gate780(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate781(.a(s_33), .b(gate438inter3), .O(gate438inter10));
  nor2  gate782(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate783(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate784(.a(gate438inter12), .b(gate438inter1), .O(G1247));

  xor2  gate869(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate870(.a(gate439inter0), .b(s_46), .O(gate439inter1));
  and2  gate871(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate872(.a(s_46), .O(gate439inter3));
  inv1  gate873(.a(s_47), .O(gate439inter4));
  nand2 gate874(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate875(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate876(.a(G11), .O(gate439inter7));
  inv1  gate877(.a(G1162), .O(gate439inter8));
  nand2 gate878(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate879(.a(s_47), .b(gate439inter3), .O(gate439inter10));
  nor2  gate880(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate881(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate882(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate841(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate842(.a(gate459inter0), .b(s_42), .O(gate459inter1));
  and2  gate843(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate844(.a(s_42), .O(gate459inter3));
  inv1  gate845(.a(s_43), .O(gate459inter4));
  nand2 gate846(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate847(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate848(.a(G21), .O(gate459inter7));
  inv1  gate849(.a(G1192), .O(gate459inter8));
  nand2 gate850(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate851(.a(s_43), .b(gate459inter3), .O(gate459inter10));
  nor2  gate852(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate853(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate854(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate1247(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate1248(.a(gate492inter0), .b(s_100), .O(gate492inter1));
  and2  gate1249(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate1250(.a(s_100), .O(gate492inter3));
  inv1  gate1251(.a(s_101), .O(gate492inter4));
  nand2 gate1252(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate1253(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate1254(.a(G1246), .O(gate492inter7));
  inv1  gate1255(.a(G1247), .O(gate492inter8));
  nand2 gate1256(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate1257(.a(s_101), .b(gate492inter3), .O(gate492inter10));
  nor2  gate1258(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate1259(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate1260(.a(gate492inter12), .b(gate492inter1), .O(G1301));
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );

  xor2  gate1219(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate1220(.a(gate507inter0), .b(s_96), .O(gate507inter1));
  and2  gate1221(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate1222(.a(s_96), .O(gate507inter3));
  inv1  gate1223(.a(s_97), .O(gate507inter4));
  nand2 gate1224(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate1225(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate1226(.a(G1276), .O(gate507inter7));
  inv1  gate1227(.a(G1277), .O(gate507inter8));
  nand2 gate1228(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate1229(.a(s_97), .b(gate507inter3), .O(gate507inter10));
  nor2  gate1230(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate1231(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate1232(.a(gate507inter12), .b(gate507inter1), .O(G1316));

  xor2  gate925(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate926(.a(gate508inter0), .b(s_54), .O(gate508inter1));
  and2  gate927(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate928(.a(s_54), .O(gate508inter3));
  inv1  gate929(.a(s_55), .O(gate508inter4));
  nand2 gate930(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate931(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate932(.a(G1278), .O(gate508inter7));
  inv1  gate933(.a(G1279), .O(gate508inter8));
  nand2 gate934(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate935(.a(s_55), .b(gate508inter3), .O(gate508inter10));
  nor2  gate936(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate937(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate938(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate827(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate828(.a(gate510inter0), .b(s_40), .O(gate510inter1));
  and2  gate829(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate830(.a(s_40), .O(gate510inter3));
  inv1  gate831(.a(s_41), .O(gate510inter4));
  nand2 gate832(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate833(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate834(.a(G1282), .O(gate510inter7));
  inv1  gate835(.a(G1283), .O(gate510inter8));
  nand2 gate836(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate837(.a(s_41), .b(gate510inter3), .O(gate510inter10));
  nor2  gate838(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate839(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate840(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule