module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate502inter0, gate502inter1, gate502inter2, gate502inter3, gate502inter4, gate502inter5, gate502inter6, gate502inter7, gate502inter8, gate502inter9, gate502inter10, gate502inter11, gate502inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate2283(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate2284(.a(gate11inter0), .b(s_248), .O(gate11inter1));
  and2  gate2285(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate2286(.a(s_248), .O(gate11inter3));
  inv1  gate2287(.a(s_249), .O(gate11inter4));
  nand2 gate2288(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate2289(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate2290(.a(G5), .O(gate11inter7));
  inv1  gate2291(.a(G6), .O(gate11inter8));
  nand2 gate2292(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate2293(.a(s_249), .b(gate11inter3), .O(gate11inter10));
  nor2  gate2294(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate2295(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate2296(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate2241(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate2242(.a(gate15inter0), .b(s_242), .O(gate15inter1));
  and2  gate2243(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate2244(.a(s_242), .O(gate15inter3));
  inv1  gate2245(.a(s_243), .O(gate15inter4));
  nand2 gate2246(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate2247(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate2248(.a(G13), .O(gate15inter7));
  inv1  gate2249(.a(G14), .O(gate15inter8));
  nand2 gate2250(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate2251(.a(s_243), .b(gate15inter3), .O(gate15inter10));
  nor2  gate2252(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate2253(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate2254(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );

  xor2  gate1681(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate1682(.a(gate18inter0), .b(s_162), .O(gate18inter1));
  and2  gate1683(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate1684(.a(s_162), .O(gate18inter3));
  inv1  gate1685(.a(s_163), .O(gate18inter4));
  nand2 gate1686(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate1687(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate1688(.a(G19), .O(gate18inter7));
  inv1  gate1689(.a(G20), .O(gate18inter8));
  nand2 gate1690(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate1691(.a(s_163), .b(gate18inter3), .O(gate18inter10));
  nor2  gate1692(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate1693(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate1694(.a(gate18inter12), .b(gate18inter1), .O(G293));

  xor2  gate1751(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate1752(.a(gate19inter0), .b(s_172), .O(gate19inter1));
  and2  gate1753(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate1754(.a(s_172), .O(gate19inter3));
  inv1  gate1755(.a(s_173), .O(gate19inter4));
  nand2 gate1756(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate1757(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate1758(.a(G21), .O(gate19inter7));
  inv1  gate1759(.a(G22), .O(gate19inter8));
  nand2 gate1760(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate1761(.a(s_173), .b(gate19inter3), .O(gate19inter10));
  nor2  gate1762(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate1763(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate1764(.a(gate19inter12), .b(gate19inter1), .O(G296));

  xor2  gate1583(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate1584(.a(gate20inter0), .b(s_148), .O(gate20inter1));
  and2  gate1585(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate1586(.a(s_148), .O(gate20inter3));
  inv1  gate1587(.a(s_149), .O(gate20inter4));
  nand2 gate1588(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate1589(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate1590(.a(G23), .O(gate20inter7));
  inv1  gate1591(.a(G24), .O(gate20inter8));
  nand2 gate1592(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate1593(.a(s_149), .b(gate20inter3), .O(gate20inter10));
  nor2  gate1594(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate1595(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate1596(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate2171(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate2172(.a(gate25inter0), .b(s_232), .O(gate25inter1));
  and2  gate2173(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate2174(.a(s_232), .O(gate25inter3));
  inv1  gate2175(.a(s_233), .O(gate25inter4));
  nand2 gate2176(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate2177(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate2178(.a(G1), .O(gate25inter7));
  inv1  gate2179(.a(G5), .O(gate25inter8));
  nand2 gate2180(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate2181(.a(s_233), .b(gate25inter3), .O(gate25inter10));
  nor2  gate2182(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate2183(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate2184(.a(gate25inter12), .b(gate25inter1), .O(G314));

  xor2  gate2423(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate2424(.a(gate26inter0), .b(s_268), .O(gate26inter1));
  and2  gate2425(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate2426(.a(s_268), .O(gate26inter3));
  inv1  gate2427(.a(s_269), .O(gate26inter4));
  nand2 gate2428(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate2429(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate2430(.a(G9), .O(gate26inter7));
  inv1  gate2431(.a(G13), .O(gate26inter8));
  nand2 gate2432(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate2433(.a(s_269), .b(gate26inter3), .O(gate26inter10));
  nor2  gate2434(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate2435(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate2436(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate2353(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate2354(.a(gate31inter0), .b(s_258), .O(gate31inter1));
  and2  gate2355(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate2356(.a(s_258), .O(gate31inter3));
  inv1  gate2357(.a(s_259), .O(gate31inter4));
  nand2 gate2358(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate2359(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate2360(.a(G4), .O(gate31inter7));
  inv1  gate2361(.a(G8), .O(gate31inter8));
  nand2 gate2362(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate2363(.a(s_259), .b(gate31inter3), .O(gate31inter10));
  nor2  gate2364(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate2365(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate2366(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate2409(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate2410(.a(gate33inter0), .b(s_266), .O(gate33inter1));
  and2  gate2411(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate2412(.a(s_266), .O(gate33inter3));
  inv1  gate2413(.a(s_267), .O(gate33inter4));
  nand2 gate2414(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate2415(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate2416(.a(G17), .O(gate33inter7));
  inv1  gate2417(.a(G21), .O(gate33inter8));
  nand2 gate2418(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate2419(.a(s_267), .b(gate33inter3), .O(gate33inter10));
  nor2  gate2420(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate2421(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate2422(.a(gate33inter12), .b(gate33inter1), .O(G338));

  xor2  gate603(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate604(.a(gate34inter0), .b(s_8), .O(gate34inter1));
  and2  gate605(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate606(.a(s_8), .O(gate34inter3));
  inv1  gate607(.a(s_9), .O(gate34inter4));
  nand2 gate608(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate609(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate610(.a(G25), .O(gate34inter7));
  inv1  gate611(.a(G29), .O(gate34inter8));
  nand2 gate612(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate613(.a(s_9), .b(gate34inter3), .O(gate34inter10));
  nor2  gate614(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate615(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate616(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate1387(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1388(.a(gate36inter0), .b(s_120), .O(gate36inter1));
  and2  gate1389(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1390(.a(s_120), .O(gate36inter3));
  inv1  gate1391(.a(s_121), .O(gate36inter4));
  nand2 gate1392(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1393(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1394(.a(G26), .O(gate36inter7));
  inv1  gate1395(.a(G30), .O(gate36inter8));
  nand2 gate1396(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1397(.a(s_121), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1398(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1399(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1400(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate869(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate870(.a(gate43inter0), .b(s_46), .O(gate43inter1));
  and2  gate871(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate872(.a(s_46), .O(gate43inter3));
  inv1  gate873(.a(s_47), .O(gate43inter4));
  nand2 gate874(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate875(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate876(.a(G3), .O(gate43inter7));
  inv1  gate877(.a(G269), .O(gate43inter8));
  nand2 gate878(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate879(.a(s_47), .b(gate43inter3), .O(gate43inter10));
  nor2  gate880(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate881(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate882(.a(gate43inter12), .b(gate43inter1), .O(G364));
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate1219(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate1220(.a(gate46inter0), .b(s_96), .O(gate46inter1));
  and2  gate1221(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate1222(.a(s_96), .O(gate46inter3));
  inv1  gate1223(.a(s_97), .O(gate46inter4));
  nand2 gate1224(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate1225(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate1226(.a(G6), .O(gate46inter7));
  inv1  gate1227(.a(G272), .O(gate46inter8));
  nand2 gate1228(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate1229(.a(s_97), .b(gate46inter3), .O(gate46inter10));
  nor2  gate1230(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate1231(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate1232(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );

  xor2  gate743(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate744(.a(gate53inter0), .b(s_28), .O(gate53inter1));
  and2  gate745(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate746(.a(s_28), .O(gate53inter3));
  inv1  gate747(.a(s_29), .O(gate53inter4));
  nand2 gate748(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate749(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate750(.a(G13), .O(gate53inter7));
  inv1  gate751(.a(G284), .O(gate53inter8));
  nand2 gate752(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate753(.a(s_29), .b(gate53inter3), .O(gate53inter10));
  nor2  gate754(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate755(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate756(.a(gate53inter12), .b(gate53inter1), .O(G374));
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate1821(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate1822(.a(gate60inter0), .b(s_182), .O(gate60inter1));
  and2  gate1823(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate1824(.a(s_182), .O(gate60inter3));
  inv1  gate1825(.a(s_183), .O(gate60inter4));
  nand2 gate1826(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate1827(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate1828(.a(G20), .O(gate60inter7));
  inv1  gate1829(.a(G293), .O(gate60inter8));
  nand2 gate1830(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate1831(.a(s_183), .b(gate60inter3), .O(gate60inter10));
  nor2  gate1832(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate1833(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate1834(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate2017(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate2018(.a(gate62inter0), .b(s_210), .O(gate62inter1));
  and2  gate2019(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate2020(.a(s_210), .O(gate62inter3));
  inv1  gate2021(.a(s_211), .O(gate62inter4));
  nand2 gate2022(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate2023(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate2024(.a(G22), .O(gate62inter7));
  inv1  gate2025(.a(G296), .O(gate62inter8));
  nand2 gate2026(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate2027(.a(s_211), .b(gate62inter3), .O(gate62inter10));
  nor2  gate2028(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate2029(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate2030(.a(gate62inter12), .b(gate62inter1), .O(G383));

  xor2  gate2073(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate2074(.a(gate63inter0), .b(s_218), .O(gate63inter1));
  and2  gate2075(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate2076(.a(s_218), .O(gate63inter3));
  inv1  gate2077(.a(s_219), .O(gate63inter4));
  nand2 gate2078(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate2079(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate2080(.a(G23), .O(gate63inter7));
  inv1  gate2081(.a(G299), .O(gate63inter8));
  nand2 gate2082(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate2083(.a(s_219), .b(gate63inter3), .O(gate63inter10));
  nor2  gate2084(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate2085(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate2086(.a(gate63inter12), .b(gate63inter1), .O(G384));

  xor2  gate1177(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate1178(.a(gate64inter0), .b(s_90), .O(gate64inter1));
  and2  gate1179(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate1180(.a(s_90), .O(gate64inter3));
  inv1  gate1181(.a(s_91), .O(gate64inter4));
  nand2 gate1182(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate1183(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate1184(.a(G24), .O(gate64inter7));
  inv1  gate1185(.a(G299), .O(gate64inter8));
  nand2 gate1186(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate1187(.a(s_91), .b(gate64inter3), .O(gate64inter10));
  nor2  gate1188(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate1189(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate1190(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate1723(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate1724(.a(gate66inter0), .b(s_168), .O(gate66inter1));
  and2  gate1725(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate1726(.a(s_168), .O(gate66inter3));
  inv1  gate1727(.a(s_169), .O(gate66inter4));
  nand2 gate1728(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate1729(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate1730(.a(G26), .O(gate66inter7));
  inv1  gate1731(.a(G302), .O(gate66inter8));
  nand2 gate1732(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate1733(.a(s_169), .b(gate66inter3), .O(gate66inter10));
  nor2  gate1734(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate1735(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate1736(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );

  xor2  gate1569(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate1570(.a(gate68inter0), .b(s_146), .O(gate68inter1));
  and2  gate1571(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate1572(.a(s_146), .O(gate68inter3));
  inv1  gate1573(.a(s_147), .O(gate68inter4));
  nand2 gate1574(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate1575(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate1576(.a(G28), .O(gate68inter7));
  inv1  gate1577(.a(G305), .O(gate68inter8));
  nand2 gate1578(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate1579(.a(s_147), .b(gate68inter3), .O(gate68inter10));
  nor2  gate1580(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate1581(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate1582(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate547(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate548(.a(gate70inter0), .b(s_0), .O(gate70inter1));
  and2  gate549(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate550(.a(s_0), .O(gate70inter3));
  inv1  gate551(.a(s_1), .O(gate70inter4));
  nand2 gate552(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate553(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate554(.a(G30), .O(gate70inter7));
  inv1  gate555(.a(G308), .O(gate70inter8));
  nand2 gate556(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate557(.a(s_1), .b(gate70inter3), .O(gate70inter10));
  nor2  gate558(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate559(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate560(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );

  xor2  gate827(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate828(.a(gate73inter0), .b(s_40), .O(gate73inter1));
  and2  gate829(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate830(.a(s_40), .O(gate73inter3));
  inv1  gate831(.a(s_41), .O(gate73inter4));
  nand2 gate832(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate833(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate834(.a(G1), .O(gate73inter7));
  inv1  gate835(.a(G314), .O(gate73inter8));
  nand2 gate836(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate837(.a(s_41), .b(gate73inter3), .O(gate73inter10));
  nor2  gate838(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate839(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate840(.a(gate73inter12), .b(gate73inter1), .O(G394));

  xor2  gate897(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate898(.a(gate74inter0), .b(s_50), .O(gate74inter1));
  and2  gate899(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate900(.a(s_50), .O(gate74inter3));
  inv1  gate901(.a(s_51), .O(gate74inter4));
  nand2 gate902(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate903(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate904(.a(G5), .O(gate74inter7));
  inv1  gate905(.a(G314), .O(gate74inter8));
  nand2 gate906(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate907(.a(s_51), .b(gate74inter3), .O(gate74inter10));
  nor2  gate908(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate909(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate910(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate1149(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate1150(.a(gate77inter0), .b(s_86), .O(gate77inter1));
  and2  gate1151(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate1152(.a(s_86), .O(gate77inter3));
  inv1  gate1153(.a(s_87), .O(gate77inter4));
  nand2 gate1154(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate1155(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate1156(.a(G2), .O(gate77inter7));
  inv1  gate1157(.a(G320), .O(gate77inter8));
  nand2 gate1158(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate1159(.a(s_87), .b(gate77inter3), .O(gate77inter10));
  nor2  gate1160(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate1161(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate1162(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate1835(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate1836(.a(gate81inter0), .b(s_184), .O(gate81inter1));
  and2  gate1837(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate1838(.a(s_184), .O(gate81inter3));
  inv1  gate1839(.a(s_185), .O(gate81inter4));
  nand2 gate1840(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate1841(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate1842(.a(G3), .O(gate81inter7));
  inv1  gate1843(.a(G326), .O(gate81inter8));
  nand2 gate1844(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate1845(.a(s_185), .b(gate81inter3), .O(gate81inter10));
  nor2  gate1846(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate1847(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate1848(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate1527(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate1528(.a(gate85inter0), .b(s_140), .O(gate85inter1));
  and2  gate1529(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate1530(.a(s_140), .O(gate85inter3));
  inv1  gate1531(.a(s_141), .O(gate85inter4));
  nand2 gate1532(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate1533(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate1534(.a(G4), .O(gate85inter7));
  inv1  gate1535(.a(G332), .O(gate85inter8));
  nand2 gate1536(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate1537(.a(s_141), .b(gate85inter3), .O(gate85inter10));
  nor2  gate1538(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate1539(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate1540(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate2199(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate2200(.a(gate91inter0), .b(s_236), .O(gate91inter1));
  and2  gate2201(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate2202(.a(s_236), .O(gate91inter3));
  inv1  gate2203(.a(s_237), .O(gate91inter4));
  nand2 gate2204(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate2205(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate2206(.a(G25), .O(gate91inter7));
  inv1  gate2207(.a(G341), .O(gate91inter8));
  nand2 gate2208(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate2209(.a(s_237), .b(gate91inter3), .O(gate91inter10));
  nor2  gate2210(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate2211(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate2212(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate1625(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate1626(.a(gate96inter0), .b(s_154), .O(gate96inter1));
  and2  gate1627(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate1628(.a(s_154), .O(gate96inter3));
  inv1  gate1629(.a(s_155), .O(gate96inter4));
  nand2 gate1630(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate1631(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate1632(.a(G30), .O(gate96inter7));
  inv1  gate1633(.a(G347), .O(gate96inter8));
  nand2 gate1634(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate1635(.a(s_155), .b(gate96inter3), .O(gate96inter10));
  nor2  gate1636(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate1637(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate1638(.a(gate96inter12), .b(gate96inter1), .O(G417));
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate687(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate688(.a(gate99inter0), .b(s_20), .O(gate99inter1));
  and2  gate689(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate690(.a(s_20), .O(gate99inter3));
  inv1  gate691(.a(s_21), .O(gate99inter4));
  nand2 gate692(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate693(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate694(.a(G27), .O(gate99inter7));
  inv1  gate695(.a(G353), .O(gate99inter8));
  nand2 gate696(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate697(.a(s_21), .b(gate99inter3), .O(gate99inter10));
  nor2  gate698(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate699(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate700(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate673(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate674(.a(gate106inter0), .b(s_18), .O(gate106inter1));
  and2  gate675(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate676(.a(s_18), .O(gate106inter3));
  inv1  gate677(.a(s_19), .O(gate106inter4));
  nand2 gate678(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate679(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate680(.a(G364), .O(gate106inter7));
  inv1  gate681(.a(G365), .O(gate106inter8));
  nand2 gate682(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate683(.a(s_19), .b(gate106inter3), .O(gate106inter10));
  nor2  gate684(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate685(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate686(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate1289(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate1290(.a(gate109inter0), .b(s_106), .O(gate109inter1));
  and2  gate1291(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate1292(.a(s_106), .O(gate109inter3));
  inv1  gate1293(.a(s_107), .O(gate109inter4));
  nand2 gate1294(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate1295(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate1296(.a(G370), .O(gate109inter7));
  inv1  gate1297(.a(G371), .O(gate109inter8));
  nand2 gate1298(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate1299(.a(s_107), .b(gate109inter3), .O(gate109inter10));
  nor2  gate1300(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate1301(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate1302(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );

  xor2  gate1121(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate1122(.a(gate111inter0), .b(s_82), .O(gate111inter1));
  and2  gate1123(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate1124(.a(s_82), .O(gate111inter3));
  inv1  gate1125(.a(s_83), .O(gate111inter4));
  nand2 gate1126(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate1127(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate1128(.a(G374), .O(gate111inter7));
  inv1  gate1129(.a(G375), .O(gate111inter8));
  nand2 gate1130(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate1131(.a(s_83), .b(gate111inter3), .O(gate111inter10));
  nor2  gate1132(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate1133(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate1134(.a(gate111inter12), .b(gate111inter1), .O(G444));
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate561(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate562(.a(gate118inter0), .b(s_2), .O(gate118inter1));
  and2  gate563(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate564(.a(s_2), .O(gate118inter3));
  inv1  gate565(.a(s_3), .O(gate118inter4));
  nand2 gate566(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate567(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate568(.a(G388), .O(gate118inter7));
  inv1  gate569(.a(G389), .O(gate118inter8));
  nand2 gate570(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate571(.a(s_3), .b(gate118inter3), .O(gate118inter10));
  nor2  gate572(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate573(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate574(.a(gate118inter12), .b(gate118inter1), .O(G465));

  xor2  gate1191(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate1192(.a(gate119inter0), .b(s_92), .O(gate119inter1));
  and2  gate1193(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate1194(.a(s_92), .O(gate119inter3));
  inv1  gate1195(.a(s_93), .O(gate119inter4));
  nand2 gate1196(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate1197(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate1198(.a(G390), .O(gate119inter7));
  inv1  gate1199(.a(G391), .O(gate119inter8));
  nand2 gate1200(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate1201(.a(s_93), .b(gate119inter3), .O(gate119inter10));
  nor2  gate1202(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate1203(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate1204(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );

  xor2  gate1345(.a(G399), .b(G398), .O(gate123inter0));
  nand2 gate1346(.a(gate123inter0), .b(s_114), .O(gate123inter1));
  and2  gate1347(.a(G399), .b(G398), .O(gate123inter2));
  inv1  gate1348(.a(s_114), .O(gate123inter3));
  inv1  gate1349(.a(s_115), .O(gate123inter4));
  nand2 gate1350(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate1351(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate1352(.a(G398), .O(gate123inter7));
  inv1  gate1353(.a(G399), .O(gate123inter8));
  nand2 gate1354(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate1355(.a(s_115), .b(gate123inter3), .O(gate123inter10));
  nor2  gate1356(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate1357(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate1358(.a(gate123inter12), .b(gate123inter1), .O(G480));
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );

  xor2  gate883(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate884(.a(gate133inter0), .b(s_48), .O(gate133inter1));
  and2  gate885(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate886(.a(s_48), .O(gate133inter3));
  inv1  gate887(.a(s_49), .O(gate133inter4));
  nand2 gate888(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate889(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate890(.a(G418), .O(gate133inter7));
  inv1  gate891(.a(G419), .O(gate133inter8));
  nand2 gate892(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate893(.a(s_49), .b(gate133inter3), .O(gate133inter10));
  nor2  gate894(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate895(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate896(.a(gate133inter12), .b(gate133inter1), .O(G510));
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate1135(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate1136(.a(gate135inter0), .b(s_84), .O(gate135inter1));
  and2  gate1137(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate1138(.a(s_84), .O(gate135inter3));
  inv1  gate1139(.a(s_85), .O(gate135inter4));
  nand2 gate1140(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate1141(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate1142(.a(G422), .O(gate135inter7));
  inv1  gate1143(.a(G423), .O(gate135inter8));
  nand2 gate1144(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate1145(.a(s_85), .b(gate135inter3), .O(gate135inter10));
  nor2  gate1146(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate1147(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate1148(.a(gate135inter12), .b(gate135inter1), .O(G516));
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate2255(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate2256(.a(gate137inter0), .b(s_244), .O(gate137inter1));
  and2  gate2257(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate2258(.a(s_244), .O(gate137inter3));
  inv1  gate2259(.a(s_245), .O(gate137inter4));
  nand2 gate2260(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate2261(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate2262(.a(G426), .O(gate137inter7));
  inv1  gate2263(.a(G429), .O(gate137inter8));
  nand2 gate2264(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate2265(.a(s_245), .b(gate137inter3), .O(gate137inter10));
  nor2  gate2266(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate2267(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate2268(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate1863(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate1864(.a(gate142inter0), .b(s_188), .O(gate142inter1));
  and2  gate1865(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate1866(.a(s_188), .O(gate142inter3));
  inv1  gate1867(.a(s_189), .O(gate142inter4));
  nand2 gate1868(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate1869(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate1870(.a(G456), .O(gate142inter7));
  inv1  gate1871(.a(G459), .O(gate142inter8));
  nand2 gate1872(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate1873(.a(s_189), .b(gate142inter3), .O(gate142inter10));
  nor2  gate1874(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate1875(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate1876(.a(gate142inter12), .b(gate142inter1), .O(G537));

  xor2  gate1163(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate1164(.a(gate143inter0), .b(s_88), .O(gate143inter1));
  and2  gate1165(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate1166(.a(s_88), .O(gate143inter3));
  inv1  gate1167(.a(s_89), .O(gate143inter4));
  nand2 gate1168(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate1169(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate1170(.a(G462), .O(gate143inter7));
  inv1  gate1171(.a(G465), .O(gate143inter8));
  nand2 gate1172(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate1173(.a(s_89), .b(gate143inter3), .O(gate143inter10));
  nor2  gate1174(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate1175(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate1176(.a(gate143inter12), .b(gate143inter1), .O(G540));
nand2 gate144( .a(G468), .b(G471), .O(G543) );

  xor2  gate1779(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate1780(.a(gate145inter0), .b(s_176), .O(gate145inter1));
  and2  gate1781(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate1782(.a(s_176), .O(gate145inter3));
  inv1  gate1783(.a(s_177), .O(gate145inter4));
  nand2 gate1784(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate1785(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate1786(.a(G474), .O(gate145inter7));
  inv1  gate1787(.a(G477), .O(gate145inter8));
  nand2 gate1788(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate1789(.a(s_177), .b(gate145inter3), .O(gate145inter10));
  nor2  gate1790(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate1791(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate1792(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate1695(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1696(.a(gate148inter0), .b(s_164), .O(gate148inter1));
  and2  gate1697(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1698(.a(s_164), .O(gate148inter3));
  inv1  gate1699(.a(s_165), .O(gate148inter4));
  nand2 gate1700(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1701(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1702(.a(G492), .O(gate148inter7));
  inv1  gate1703(.a(G495), .O(gate148inter8));
  nand2 gate1704(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1705(.a(s_165), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1706(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1707(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1708(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate1877(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate1878(.a(gate155inter0), .b(s_190), .O(gate155inter1));
  and2  gate1879(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate1880(.a(s_190), .O(gate155inter3));
  inv1  gate1881(.a(s_191), .O(gate155inter4));
  nand2 gate1882(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1883(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1884(.a(G432), .O(gate155inter7));
  inv1  gate1885(.a(G525), .O(gate155inter8));
  nand2 gate1886(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1887(.a(s_191), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1888(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1889(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1890(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate1205(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate1206(.a(gate157inter0), .b(s_94), .O(gate157inter1));
  and2  gate1207(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate1208(.a(s_94), .O(gate157inter3));
  inv1  gate1209(.a(s_95), .O(gate157inter4));
  nand2 gate1210(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate1211(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate1212(.a(G438), .O(gate157inter7));
  inv1  gate1213(.a(G528), .O(gate157inter8));
  nand2 gate1214(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate1215(.a(s_95), .b(gate157inter3), .O(gate157inter10));
  nor2  gate1216(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate1217(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate1218(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate1023(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate1024(.a(gate160inter0), .b(s_68), .O(gate160inter1));
  and2  gate1025(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate1026(.a(s_68), .O(gate160inter3));
  inv1  gate1027(.a(s_69), .O(gate160inter4));
  nand2 gate1028(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate1029(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate1030(.a(G447), .O(gate160inter7));
  inv1  gate1031(.a(G531), .O(gate160inter8));
  nand2 gate1032(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate1033(.a(s_69), .b(gate160inter3), .O(gate160inter10));
  nor2  gate1034(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate1035(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate1036(.a(gate160inter12), .b(gate160inter1), .O(G577));

  xor2  gate631(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate632(.a(gate161inter0), .b(s_12), .O(gate161inter1));
  and2  gate633(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate634(.a(s_12), .O(gate161inter3));
  inv1  gate635(.a(s_13), .O(gate161inter4));
  nand2 gate636(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate637(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate638(.a(G450), .O(gate161inter7));
  inv1  gate639(.a(G534), .O(gate161inter8));
  nand2 gate640(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate641(.a(s_13), .b(gate161inter3), .O(gate161inter10));
  nor2  gate642(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate643(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate644(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate953(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate954(.a(gate165inter0), .b(s_58), .O(gate165inter1));
  and2  gate955(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate956(.a(s_58), .O(gate165inter3));
  inv1  gate957(.a(s_59), .O(gate165inter4));
  nand2 gate958(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate959(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate960(.a(G462), .O(gate165inter7));
  inv1  gate961(.a(G540), .O(gate165inter8));
  nand2 gate962(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate963(.a(s_59), .b(gate165inter3), .O(gate165inter10));
  nor2  gate964(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate965(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate966(.a(gate165inter12), .b(gate165inter1), .O(G582));

  xor2  gate1443(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate1444(.a(gate166inter0), .b(s_128), .O(gate166inter1));
  and2  gate1445(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate1446(.a(s_128), .O(gate166inter3));
  inv1  gate1447(.a(s_129), .O(gate166inter4));
  nand2 gate1448(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate1449(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate1450(.a(G465), .O(gate166inter7));
  inv1  gate1451(.a(G540), .O(gate166inter8));
  nand2 gate1452(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate1453(.a(s_129), .b(gate166inter3), .O(gate166inter10));
  nor2  gate1454(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate1455(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate1456(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate2367(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate2368(.a(gate172inter0), .b(s_260), .O(gate172inter1));
  and2  gate2369(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate2370(.a(s_260), .O(gate172inter3));
  inv1  gate2371(.a(s_261), .O(gate172inter4));
  nand2 gate2372(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate2373(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate2374(.a(G483), .O(gate172inter7));
  inv1  gate2375(.a(G549), .O(gate172inter8));
  nand2 gate2376(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate2377(.a(s_261), .b(gate172inter3), .O(gate172inter10));
  nor2  gate2378(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate2379(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate2380(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );

  xor2  gate1317(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate1318(.a(gate182inter0), .b(s_110), .O(gate182inter1));
  and2  gate1319(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate1320(.a(s_110), .O(gate182inter3));
  inv1  gate1321(.a(s_111), .O(gate182inter4));
  nand2 gate1322(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate1323(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate1324(.a(G513), .O(gate182inter7));
  inv1  gate1325(.a(G564), .O(gate182inter8));
  nand2 gate1326(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate1327(.a(s_111), .b(gate182inter3), .O(gate182inter10));
  nor2  gate1328(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate1329(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate1330(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate939(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate940(.a(gate184inter0), .b(s_56), .O(gate184inter1));
  and2  gate941(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate942(.a(s_56), .O(gate184inter3));
  inv1  gate943(.a(s_57), .O(gate184inter4));
  nand2 gate944(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate945(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate946(.a(G519), .O(gate184inter7));
  inv1  gate947(.a(G567), .O(gate184inter8));
  nand2 gate948(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate949(.a(s_57), .b(gate184inter3), .O(gate184inter10));
  nor2  gate950(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate951(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate952(.a(gate184inter12), .b(gate184inter1), .O(G601));
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate1485(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1486(.a(gate186inter0), .b(s_134), .O(gate186inter1));
  and2  gate1487(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1488(.a(s_134), .O(gate186inter3));
  inv1  gate1489(.a(s_135), .O(gate186inter4));
  nand2 gate1490(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1491(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1492(.a(G572), .O(gate186inter7));
  inv1  gate1493(.a(G573), .O(gate186inter8));
  nand2 gate1494(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1495(.a(s_135), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1496(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1497(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1498(.a(gate186inter12), .b(gate186inter1), .O(G607));

  xor2  gate841(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate842(.a(gate187inter0), .b(s_42), .O(gate187inter1));
  and2  gate843(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate844(.a(s_42), .O(gate187inter3));
  inv1  gate845(.a(s_43), .O(gate187inter4));
  nand2 gate846(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate847(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate848(.a(G574), .O(gate187inter7));
  inv1  gate849(.a(G575), .O(gate187inter8));
  nand2 gate850(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate851(.a(s_43), .b(gate187inter3), .O(gate187inter10));
  nor2  gate852(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate853(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate854(.a(gate187inter12), .b(gate187inter1), .O(G612));

  xor2  gate1639(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate1640(.a(gate188inter0), .b(s_156), .O(gate188inter1));
  and2  gate1641(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate1642(.a(s_156), .O(gate188inter3));
  inv1  gate1643(.a(s_157), .O(gate188inter4));
  nand2 gate1644(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate1645(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate1646(.a(G576), .O(gate188inter7));
  inv1  gate1647(.a(G577), .O(gate188inter8));
  nand2 gate1648(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate1649(.a(s_157), .b(gate188inter3), .O(gate188inter10));
  nor2  gate1650(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate1651(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate1652(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate2143(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate2144(.a(gate195inter0), .b(s_228), .O(gate195inter1));
  and2  gate2145(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate2146(.a(s_228), .O(gate195inter3));
  inv1  gate2147(.a(s_229), .O(gate195inter4));
  nand2 gate2148(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate2149(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate2150(.a(G590), .O(gate195inter7));
  inv1  gate2151(.a(G591), .O(gate195inter8));
  nand2 gate2152(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate2153(.a(s_229), .b(gate195inter3), .O(gate195inter10));
  nor2  gate2154(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate2155(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate2156(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate729(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate730(.a(gate197inter0), .b(s_26), .O(gate197inter1));
  and2  gate731(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate732(.a(s_26), .O(gate197inter3));
  inv1  gate733(.a(s_27), .O(gate197inter4));
  nand2 gate734(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate735(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate736(.a(G594), .O(gate197inter7));
  inv1  gate737(.a(G595), .O(gate197inter8));
  nand2 gate738(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate739(.a(s_27), .b(gate197inter3), .O(gate197inter10));
  nor2  gate740(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate741(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate742(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate2115(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate2116(.a(gate200inter0), .b(s_224), .O(gate200inter1));
  and2  gate2117(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate2118(.a(s_224), .O(gate200inter3));
  inv1  gate2119(.a(s_225), .O(gate200inter4));
  nand2 gate2120(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate2121(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate2122(.a(G600), .O(gate200inter7));
  inv1  gate2123(.a(G601), .O(gate200inter8));
  nand2 gate2124(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate2125(.a(s_225), .b(gate200inter3), .O(gate200inter10));
  nor2  gate2126(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate2127(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate2128(.a(gate200inter12), .b(gate200inter1), .O(G663));
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );

  xor2  gate813(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate814(.a(gate204inter0), .b(s_38), .O(gate204inter1));
  and2  gate815(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate816(.a(s_38), .O(gate204inter3));
  inv1  gate817(.a(s_39), .O(gate204inter4));
  nand2 gate818(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate819(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate820(.a(G607), .O(gate204inter7));
  inv1  gate821(.a(G617), .O(gate204inter8));
  nand2 gate822(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate823(.a(s_39), .b(gate204inter3), .O(gate204inter10));
  nor2  gate824(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate825(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate826(.a(gate204inter12), .b(gate204inter1), .O(G675));

  xor2  gate2297(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate2298(.a(gate205inter0), .b(s_250), .O(gate205inter1));
  and2  gate2299(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate2300(.a(s_250), .O(gate205inter3));
  inv1  gate2301(.a(s_251), .O(gate205inter4));
  nand2 gate2302(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate2303(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate2304(.a(G622), .O(gate205inter7));
  inv1  gate2305(.a(G627), .O(gate205inter8));
  nand2 gate2306(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate2307(.a(s_251), .b(gate205inter3), .O(gate205inter10));
  nor2  gate2308(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate2309(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate2310(.a(gate205inter12), .b(gate205inter1), .O(G678));

  xor2  gate785(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate786(.a(gate206inter0), .b(s_34), .O(gate206inter1));
  and2  gate787(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate788(.a(s_34), .O(gate206inter3));
  inv1  gate789(.a(s_35), .O(gate206inter4));
  nand2 gate790(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate791(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate792(.a(G632), .O(gate206inter7));
  inv1  gate793(.a(G637), .O(gate206inter8));
  nand2 gate794(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate795(.a(s_35), .b(gate206inter3), .O(gate206inter10));
  nor2  gate796(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate797(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate798(.a(gate206inter12), .b(gate206inter1), .O(G681));

  xor2  gate981(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate982(.a(gate207inter0), .b(s_62), .O(gate207inter1));
  and2  gate983(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate984(.a(s_62), .O(gate207inter3));
  inv1  gate985(.a(s_63), .O(gate207inter4));
  nand2 gate986(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate987(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate988(.a(G622), .O(gate207inter7));
  inv1  gate989(.a(G632), .O(gate207inter8));
  nand2 gate990(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate991(.a(s_63), .b(gate207inter3), .O(gate207inter10));
  nor2  gate992(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate993(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate994(.a(gate207inter12), .b(gate207inter1), .O(G684));

  xor2  gate1107(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate1108(.a(gate208inter0), .b(s_80), .O(gate208inter1));
  and2  gate1109(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate1110(.a(s_80), .O(gate208inter3));
  inv1  gate1111(.a(s_81), .O(gate208inter4));
  nand2 gate1112(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate1113(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate1114(.a(G627), .O(gate208inter7));
  inv1  gate1115(.a(G637), .O(gate208inter8));
  nand2 gate1116(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate1117(.a(s_81), .b(gate208inter3), .O(gate208inter10));
  nor2  gate1118(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate1119(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate1120(.a(gate208inter12), .b(gate208inter1), .O(G687));
nand2 gate209( .a(G602), .b(G666), .O(G690) );

  xor2  gate2003(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate2004(.a(gate210inter0), .b(s_208), .O(gate210inter1));
  and2  gate2005(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate2006(.a(s_208), .O(gate210inter3));
  inv1  gate2007(.a(s_209), .O(gate210inter4));
  nand2 gate2008(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate2009(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate2010(.a(G607), .O(gate210inter7));
  inv1  gate2011(.a(G666), .O(gate210inter8));
  nand2 gate2012(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate2013(.a(s_209), .b(gate210inter3), .O(gate210inter10));
  nor2  gate2014(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate2015(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate2016(.a(gate210inter12), .b(gate210inter1), .O(G691));
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate1933(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate1934(.a(gate214inter0), .b(s_198), .O(gate214inter1));
  and2  gate1935(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate1936(.a(s_198), .O(gate214inter3));
  inv1  gate1937(.a(s_199), .O(gate214inter4));
  nand2 gate1938(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate1939(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate1940(.a(G612), .O(gate214inter7));
  inv1  gate1941(.a(G672), .O(gate214inter8));
  nand2 gate1942(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate1943(.a(s_199), .b(gate214inter3), .O(gate214inter10));
  nor2  gate1944(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate1945(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate1946(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate2031(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate2032(.a(gate216inter0), .b(s_212), .O(gate216inter1));
  and2  gate2033(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate2034(.a(s_212), .O(gate216inter3));
  inv1  gate2035(.a(s_213), .O(gate216inter4));
  nand2 gate2036(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate2037(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate2038(.a(G617), .O(gate216inter7));
  inv1  gate2039(.a(G675), .O(gate216inter8));
  nand2 gate2040(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate2041(.a(s_213), .b(gate216inter3), .O(gate216inter10));
  nor2  gate2042(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate2043(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate2044(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate2157(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate2158(.a(gate218inter0), .b(s_230), .O(gate218inter1));
  and2  gate2159(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate2160(.a(s_230), .O(gate218inter3));
  inv1  gate2161(.a(s_231), .O(gate218inter4));
  nand2 gate2162(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate2163(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate2164(.a(G627), .O(gate218inter7));
  inv1  gate2165(.a(G678), .O(gate218inter8));
  nand2 gate2166(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate2167(.a(s_231), .b(gate218inter3), .O(gate218inter10));
  nor2  gate2168(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate2169(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate2170(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate2437(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate2438(.a(gate228inter0), .b(s_270), .O(gate228inter1));
  and2  gate2439(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate2440(.a(s_270), .O(gate228inter3));
  inv1  gate2441(.a(s_271), .O(gate228inter4));
  nand2 gate2442(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate2443(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate2444(.a(G696), .O(gate228inter7));
  inv1  gate2445(.a(G697), .O(gate228inter8));
  nand2 gate2446(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate2447(.a(s_271), .b(gate228inter3), .O(gate228inter10));
  nor2  gate2448(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate2449(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate2450(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate1849(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate1850(.a(gate234inter0), .b(s_186), .O(gate234inter1));
  and2  gate1851(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate1852(.a(s_186), .O(gate234inter3));
  inv1  gate1853(.a(s_187), .O(gate234inter4));
  nand2 gate1854(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1855(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1856(.a(G245), .O(gate234inter7));
  inv1  gate1857(.a(G721), .O(gate234inter8));
  nand2 gate1858(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1859(.a(s_187), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1860(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1861(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1862(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate1905(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate1906(.a(gate240inter0), .b(s_194), .O(gate240inter1));
  and2  gate1907(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate1908(.a(s_194), .O(gate240inter3));
  inv1  gate1909(.a(s_195), .O(gate240inter4));
  nand2 gate1910(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate1911(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate1912(.a(G263), .O(gate240inter7));
  inv1  gate1913(.a(G715), .O(gate240inter8));
  nand2 gate1914(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate1915(.a(s_195), .b(gate240inter3), .O(gate240inter10));
  nor2  gate1916(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate1917(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate1918(.a(gate240inter12), .b(gate240inter1), .O(G751));

  xor2  gate1415(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate1416(.a(gate241inter0), .b(s_124), .O(gate241inter1));
  and2  gate1417(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate1418(.a(s_124), .O(gate241inter3));
  inv1  gate1419(.a(s_125), .O(gate241inter4));
  nand2 gate1420(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate1421(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate1422(.a(G242), .O(gate241inter7));
  inv1  gate1423(.a(G730), .O(gate241inter8));
  nand2 gate1424(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate1425(.a(s_125), .b(gate241inter3), .O(gate241inter10));
  nor2  gate1426(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate1427(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate1428(.a(gate241inter12), .b(gate241inter1), .O(G754));

  xor2  gate1499(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate1500(.a(gate242inter0), .b(s_136), .O(gate242inter1));
  and2  gate1501(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate1502(.a(s_136), .O(gate242inter3));
  inv1  gate1503(.a(s_137), .O(gate242inter4));
  nand2 gate1504(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate1505(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate1506(.a(G718), .O(gate242inter7));
  inv1  gate1507(.a(G730), .O(gate242inter8));
  nand2 gate1508(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate1509(.a(s_137), .b(gate242inter3), .O(gate242inter10));
  nor2  gate1510(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate1511(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate1512(.a(gate242inter12), .b(gate242inter1), .O(G755));

  xor2  gate925(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate926(.a(gate243inter0), .b(s_54), .O(gate243inter1));
  and2  gate927(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate928(.a(s_54), .O(gate243inter3));
  inv1  gate929(.a(s_55), .O(gate243inter4));
  nand2 gate930(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate931(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate932(.a(G245), .O(gate243inter7));
  inv1  gate933(.a(G733), .O(gate243inter8));
  nand2 gate934(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate935(.a(s_55), .b(gate243inter3), .O(gate243inter10));
  nor2  gate936(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate937(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate938(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate2213(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate2214(.a(gate245inter0), .b(s_238), .O(gate245inter1));
  and2  gate2215(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate2216(.a(s_238), .O(gate245inter3));
  inv1  gate2217(.a(s_239), .O(gate245inter4));
  nand2 gate2218(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate2219(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate2220(.a(G248), .O(gate245inter7));
  inv1  gate2221(.a(G736), .O(gate245inter8));
  nand2 gate2222(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate2223(.a(s_239), .b(gate245inter3), .O(gate245inter10));
  nor2  gate2224(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate2225(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate2226(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate1359(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate1360(.a(gate253inter0), .b(s_116), .O(gate253inter1));
  and2  gate1361(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate1362(.a(s_116), .O(gate253inter3));
  inv1  gate1363(.a(s_117), .O(gate253inter4));
  nand2 gate1364(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate1365(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate1366(.a(G260), .O(gate253inter7));
  inv1  gate1367(.a(G748), .O(gate253inter8));
  nand2 gate1368(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate1369(.a(s_117), .b(gate253inter3), .O(gate253inter10));
  nor2  gate1370(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate1371(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate1372(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );

  xor2  gate2339(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate2340(.a(gate256inter0), .b(s_256), .O(gate256inter1));
  and2  gate2341(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate2342(.a(s_256), .O(gate256inter3));
  inv1  gate2343(.a(s_257), .O(gate256inter4));
  nand2 gate2344(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate2345(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate2346(.a(G715), .O(gate256inter7));
  inv1  gate2347(.a(G751), .O(gate256inter8));
  nand2 gate2348(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate2349(.a(s_257), .b(gate256inter3), .O(gate256inter10));
  nor2  gate2350(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate2351(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate2352(.a(gate256inter12), .b(gate256inter1), .O(G769));

  xor2  gate1471(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate1472(.a(gate257inter0), .b(s_132), .O(gate257inter1));
  and2  gate1473(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate1474(.a(s_132), .O(gate257inter3));
  inv1  gate1475(.a(s_133), .O(gate257inter4));
  nand2 gate1476(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate1477(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate1478(.a(G754), .O(gate257inter7));
  inv1  gate1479(.a(G755), .O(gate257inter8));
  nand2 gate1480(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate1481(.a(s_133), .b(gate257inter3), .O(gate257inter10));
  nor2  gate1482(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate1483(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate1484(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );

  xor2  gate1079(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate1080(.a(gate260inter0), .b(s_76), .O(gate260inter1));
  and2  gate1081(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate1082(.a(s_76), .O(gate260inter3));
  inv1  gate1083(.a(s_77), .O(gate260inter4));
  nand2 gate1084(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate1085(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate1086(.a(G760), .O(gate260inter7));
  inv1  gate1087(.a(G761), .O(gate260inter8));
  nand2 gate1088(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate1089(.a(s_77), .b(gate260inter3), .O(gate260inter10));
  nor2  gate1090(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate1091(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate1092(.a(gate260inter12), .b(gate260inter1), .O(G779));

  xor2  gate1737(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate1738(.a(gate261inter0), .b(s_170), .O(gate261inter1));
  and2  gate1739(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate1740(.a(s_170), .O(gate261inter3));
  inv1  gate1741(.a(s_171), .O(gate261inter4));
  nand2 gate1742(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate1743(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate1744(.a(G762), .O(gate261inter7));
  inv1  gate1745(.a(G763), .O(gate261inter8));
  nand2 gate1746(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate1747(.a(s_171), .b(gate261inter3), .O(gate261inter10));
  nor2  gate1748(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate1749(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate1750(.a(gate261inter12), .b(gate261inter1), .O(G782));
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate589(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate590(.a(gate263inter0), .b(s_6), .O(gate263inter1));
  and2  gate591(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate592(.a(s_6), .O(gate263inter3));
  inv1  gate593(.a(s_7), .O(gate263inter4));
  nand2 gate594(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate595(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate596(.a(G766), .O(gate263inter7));
  inv1  gate597(.a(G767), .O(gate263inter8));
  nand2 gate598(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate599(.a(s_7), .b(gate263inter3), .O(gate263inter10));
  nor2  gate600(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate601(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate602(.a(gate263inter12), .b(gate263inter1), .O(G788));

  xor2  gate771(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate772(.a(gate264inter0), .b(s_32), .O(gate264inter1));
  and2  gate773(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate774(.a(s_32), .O(gate264inter3));
  inv1  gate775(.a(s_33), .O(gate264inter4));
  nand2 gate776(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate777(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate778(.a(G768), .O(gate264inter7));
  inv1  gate779(.a(G769), .O(gate264inter8));
  nand2 gate780(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate781(.a(s_33), .b(gate264inter3), .O(gate264inter10));
  nor2  gate782(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate783(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate784(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate2381(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate2382(.a(gate269inter0), .b(s_262), .O(gate269inter1));
  and2  gate2383(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate2384(.a(s_262), .O(gate269inter3));
  inv1  gate2385(.a(s_263), .O(gate269inter4));
  nand2 gate2386(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate2387(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate2388(.a(G654), .O(gate269inter7));
  inv1  gate2389(.a(G782), .O(gate269inter8));
  nand2 gate2390(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate2391(.a(s_263), .b(gate269inter3), .O(gate269inter10));
  nor2  gate2392(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate2393(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate2394(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate2129(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate2130(.a(gate271inter0), .b(s_226), .O(gate271inter1));
  and2  gate2131(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate2132(.a(s_226), .O(gate271inter3));
  inv1  gate2133(.a(s_227), .O(gate271inter4));
  nand2 gate2134(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate2135(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate2136(.a(G660), .O(gate271inter7));
  inv1  gate2137(.a(G788), .O(gate271inter8));
  nand2 gate2138(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate2139(.a(s_227), .b(gate271inter3), .O(gate271inter10));
  nor2  gate2140(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate2141(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate2142(.a(gate271inter12), .b(gate271inter1), .O(G812));

  xor2  gate2059(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate2060(.a(gate272inter0), .b(s_216), .O(gate272inter1));
  and2  gate2061(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate2062(.a(s_216), .O(gate272inter3));
  inv1  gate2063(.a(s_217), .O(gate272inter4));
  nand2 gate2064(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate2065(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate2066(.a(G663), .O(gate272inter7));
  inv1  gate2067(.a(G791), .O(gate272inter8));
  nand2 gate2068(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate2069(.a(s_217), .b(gate272inter3), .O(gate272inter10));
  nor2  gate2070(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate2071(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate2072(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );

  xor2  gate2395(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate2396(.a(gate277inter0), .b(s_264), .O(gate277inter1));
  and2  gate2397(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate2398(.a(s_264), .O(gate277inter3));
  inv1  gate2399(.a(s_265), .O(gate277inter4));
  nand2 gate2400(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate2401(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate2402(.a(G648), .O(gate277inter7));
  inv1  gate2403(.a(G800), .O(gate277inter8));
  nand2 gate2404(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate2405(.a(s_265), .b(gate277inter3), .O(gate277inter10));
  nor2  gate2406(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate2407(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate2408(.a(gate277inter12), .b(gate277inter1), .O(G822));

  xor2  gate1667(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate1668(.a(gate278inter0), .b(s_160), .O(gate278inter1));
  and2  gate1669(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate1670(.a(s_160), .O(gate278inter3));
  inv1  gate1671(.a(s_161), .O(gate278inter4));
  nand2 gate1672(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate1673(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate1674(.a(G776), .O(gate278inter7));
  inv1  gate1675(.a(G800), .O(gate278inter8));
  nand2 gate1676(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate1677(.a(s_161), .b(gate278inter3), .O(gate278inter10));
  nor2  gate1678(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate1679(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate1680(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );

  xor2  gate1611(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate1612(.a(gate281inter0), .b(s_152), .O(gate281inter1));
  and2  gate1613(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate1614(.a(s_152), .O(gate281inter3));
  inv1  gate1615(.a(s_153), .O(gate281inter4));
  nand2 gate1616(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate1617(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate1618(.a(G654), .O(gate281inter7));
  inv1  gate1619(.a(G806), .O(gate281inter8));
  nand2 gate1620(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate1621(.a(s_153), .b(gate281inter3), .O(gate281inter10));
  nor2  gate1622(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate1623(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate1624(.a(gate281inter12), .b(gate281inter1), .O(G826));

  xor2  gate1919(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate1920(.a(gate282inter0), .b(s_196), .O(gate282inter1));
  and2  gate1921(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate1922(.a(s_196), .O(gate282inter3));
  inv1  gate1923(.a(s_197), .O(gate282inter4));
  nand2 gate1924(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate1925(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate1926(.a(G782), .O(gate282inter7));
  inv1  gate1927(.a(G806), .O(gate282inter8));
  nand2 gate1928(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate1929(.a(s_197), .b(gate282inter3), .O(gate282inter10));
  nor2  gate1930(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate1931(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate1932(.a(gate282inter12), .b(gate282inter1), .O(G827));

  xor2  gate2227(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate2228(.a(gate283inter0), .b(s_240), .O(gate283inter1));
  and2  gate2229(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate2230(.a(s_240), .O(gate283inter3));
  inv1  gate2231(.a(s_241), .O(gate283inter4));
  nand2 gate2232(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate2233(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate2234(.a(G657), .O(gate283inter7));
  inv1  gate2235(.a(G809), .O(gate283inter8));
  nand2 gate2236(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate2237(.a(s_241), .b(gate283inter3), .O(gate283inter10));
  nor2  gate2238(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate2239(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate2240(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate2101(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate2102(.a(gate285inter0), .b(s_222), .O(gate285inter1));
  and2  gate2103(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate2104(.a(s_222), .O(gate285inter3));
  inv1  gate2105(.a(s_223), .O(gate285inter4));
  nand2 gate2106(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate2107(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate2108(.a(G660), .O(gate285inter7));
  inv1  gate2109(.a(G812), .O(gate285inter8));
  nand2 gate2110(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate2111(.a(s_223), .b(gate285inter3), .O(gate285inter10));
  nor2  gate2112(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate2113(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate2114(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate1597(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate1598(.a(gate287inter0), .b(s_150), .O(gate287inter1));
  and2  gate1599(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate1600(.a(s_150), .O(gate287inter3));
  inv1  gate1601(.a(s_151), .O(gate287inter4));
  nand2 gate1602(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate1603(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate1604(.a(G663), .O(gate287inter7));
  inv1  gate1605(.a(G815), .O(gate287inter8));
  nand2 gate1606(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate1607(.a(s_151), .b(gate287inter3), .O(gate287inter10));
  nor2  gate1608(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate1609(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate1610(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate1541(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate1542(.a(gate294inter0), .b(s_142), .O(gate294inter1));
  and2  gate1543(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate1544(.a(s_142), .O(gate294inter3));
  inv1  gate1545(.a(s_143), .O(gate294inter4));
  nand2 gate1546(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate1547(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate1548(.a(G832), .O(gate294inter7));
  inv1  gate1549(.a(G833), .O(gate294inter8));
  nand2 gate1550(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate1551(.a(s_143), .b(gate294inter3), .O(gate294inter10));
  nor2  gate1552(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate1553(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate1554(.a(gate294inter12), .b(gate294inter1), .O(G899));

  xor2  gate799(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate800(.a(gate295inter0), .b(s_36), .O(gate295inter1));
  and2  gate801(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate802(.a(s_36), .O(gate295inter3));
  inv1  gate803(.a(s_37), .O(gate295inter4));
  nand2 gate804(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate805(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate806(.a(G830), .O(gate295inter7));
  inv1  gate807(.a(G831), .O(gate295inter8));
  nand2 gate808(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate809(.a(s_37), .b(gate295inter3), .O(gate295inter10));
  nor2  gate810(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate811(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate812(.a(gate295inter12), .b(gate295inter1), .O(G912));
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate1765(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate1766(.a(gate390inter0), .b(s_174), .O(gate390inter1));
  and2  gate1767(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate1768(.a(s_174), .O(gate390inter3));
  inv1  gate1769(.a(s_175), .O(gate390inter4));
  nand2 gate1770(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate1771(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate1772(.a(G4), .O(gate390inter7));
  inv1  gate1773(.a(G1045), .O(gate390inter8));
  nand2 gate1774(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate1775(.a(s_175), .b(gate390inter3), .O(gate390inter10));
  nor2  gate1776(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate1777(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate1778(.a(gate390inter12), .b(gate390inter1), .O(G1141));

  xor2  gate1807(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate1808(.a(gate391inter0), .b(s_180), .O(gate391inter1));
  and2  gate1809(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate1810(.a(s_180), .O(gate391inter3));
  inv1  gate1811(.a(s_181), .O(gate391inter4));
  nand2 gate1812(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate1813(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate1814(.a(G5), .O(gate391inter7));
  inv1  gate1815(.a(G1048), .O(gate391inter8));
  nand2 gate1816(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate1817(.a(s_181), .b(gate391inter3), .O(gate391inter10));
  nor2  gate1818(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate1819(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate1820(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate1513(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate1514(.a(gate394inter0), .b(s_138), .O(gate394inter1));
  and2  gate1515(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate1516(.a(s_138), .O(gate394inter3));
  inv1  gate1517(.a(s_139), .O(gate394inter4));
  nand2 gate1518(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate1519(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate1520(.a(G8), .O(gate394inter7));
  inv1  gate1521(.a(G1057), .O(gate394inter8));
  nand2 gate1522(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate1523(.a(s_139), .b(gate394inter3), .O(gate394inter10));
  nor2  gate1524(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate1525(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate1526(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate1891(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate1892(.a(gate398inter0), .b(s_192), .O(gate398inter1));
  and2  gate1893(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate1894(.a(s_192), .O(gate398inter3));
  inv1  gate1895(.a(s_193), .O(gate398inter4));
  nand2 gate1896(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate1897(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate1898(.a(G12), .O(gate398inter7));
  inv1  gate1899(.a(G1069), .O(gate398inter8));
  nand2 gate1900(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate1901(.a(s_193), .b(gate398inter3), .O(gate398inter10));
  nor2  gate1902(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate1903(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate1904(.a(gate398inter12), .b(gate398inter1), .O(G1165));

  xor2  gate967(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate968(.a(gate399inter0), .b(s_60), .O(gate399inter1));
  and2  gate969(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate970(.a(s_60), .O(gate399inter3));
  inv1  gate971(.a(s_61), .O(gate399inter4));
  nand2 gate972(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate973(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate974(.a(G13), .O(gate399inter7));
  inv1  gate975(.a(G1072), .O(gate399inter8));
  nand2 gate976(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate977(.a(s_61), .b(gate399inter3), .O(gate399inter10));
  nor2  gate978(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate979(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate980(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate1989(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate1990(.a(gate406inter0), .b(s_206), .O(gate406inter1));
  and2  gate1991(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate1992(.a(s_206), .O(gate406inter3));
  inv1  gate1993(.a(s_207), .O(gate406inter4));
  nand2 gate1994(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate1995(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate1996(.a(G20), .O(gate406inter7));
  inv1  gate1997(.a(G1093), .O(gate406inter8));
  nand2 gate1998(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate1999(.a(s_207), .b(gate406inter3), .O(gate406inter10));
  nor2  gate2000(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate2001(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate2002(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );

  xor2  gate1975(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate1976(.a(gate412inter0), .b(s_204), .O(gate412inter1));
  and2  gate1977(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate1978(.a(s_204), .O(gate412inter3));
  inv1  gate1979(.a(s_205), .O(gate412inter4));
  nand2 gate1980(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate1981(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate1982(.a(G26), .O(gate412inter7));
  inv1  gate1983(.a(G1111), .O(gate412inter8));
  nand2 gate1984(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate1985(.a(s_205), .b(gate412inter3), .O(gate412inter10));
  nor2  gate1986(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate1987(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate1988(.a(gate412inter12), .b(gate412inter1), .O(G1207));

  xor2  gate1373(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate1374(.a(gate413inter0), .b(s_118), .O(gate413inter1));
  and2  gate1375(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate1376(.a(s_118), .O(gate413inter3));
  inv1  gate1377(.a(s_119), .O(gate413inter4));
  nand2 gate1378(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1379(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1380(.a(G27), .O(gate413inter7));
  inv1  gate1381(.a(G1114), .O(gate413inter8));
  nand2 gate1382(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1383(.a(s_119), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1384(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1385(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1386(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate2269(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate2270(.a(gate415inter0), .b(s_246), .O(gate415inter1));
  and2  gate2271(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate2272(.a(s_246), .O(gate415inter3));
  inv1  gate2273(.a(s_247), .O(gate415inter4));
  nand2 gate2274(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate2275(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate2276(.a(G29), .O(gate415inter7));
  inv1  gate2277(.a(G1120), .O(gate415inter8));
  nand2 gate2278(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate2279(.a(s_247), .b(gate415inter3), .O(gate415inter10));
  nor2  gate2280(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate2281(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate2282(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate1037(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1038(.a(gate420inter0), .b(s_70), .O(gate420inter1));
  and2  gate1039(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1040(.a(s_70), .O(gate420inter3));
  inv1  gate1041(.a(s_71), .O(gate420inter4));
  nand2 gate1042(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1043(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1044(.a(G1036), .O(gate420inter7));
  inv1  gate1045(.a(G1132), .O(gate420inter8));
  nand2 gate1046(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1047(.a(s_71), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1048(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1049(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1050(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate1275(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate1276(.a(gate431inter0), .b(s_104), .O(gate431inter1));
  and2  gate1277(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate1278(.a(s_104), .O(gate431inter3));
  inv1  gate1279(.a(s_105), .O(gate431inter4));
  nand2 gate1280(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate1281(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate1282(.a(G7), .O(gate431inter7));
  inv1  gate1283(.a(G1150), .O(gate431inter8));
  nand2 gate1284(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate1285(.a(s_105), .b(gate431inter3), .O(gate431inter10));
  nor2  gate1286(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate1287(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate1288(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate1093(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate1094(.a(gate433inter0), .b(s_78), .O(gate433inter1));
  and2  gate1095(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate1096(.a(s_78), .O(gate433inter3));
  inv1  gate1097(.a(s_79), .O(gate433inter4));
  nand2 gate1098(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate1099(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate1100(.a(G8), .O(gate433inter7));
  inv1  gate1101(.a(G1153), .O(gate433inter8));
  nand2 gate1102(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate1103(.a(s_79), .b(gate433inter3), .O(gate433inter10));
  nor2  gate1104(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate1105(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate1106(.a(gate433inter12), .b(gate433inter1), .O(G1242));

  xor2  gate855(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate856(.a(gate434inter0), .b(s_44), .O(gate434inter1));
  and2  gate857(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate858(.a(s_44), .O(gate434inter3));
  inv1  gate859(.a(s_45), .O(gate434inter4));
  nand2 gate860(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate861(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate862(.a(G1057), .O(gate434inter7));
  inv1  gate863(.a(G1153), .O(gate434inter8));
  nand2 gate864(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate865(.a(s_45), .b(gate434inter3), .O(gate434inter10));
  nor2  gate866(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate867(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate868(.a(gate434inter12), .b(gate434inter1), .O(G1243));

  xor2  gate701(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate702(.a(gate435inter0), .b(s_22), .O(gate435inter1));
  and2  gate703(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate704(.a(s_22), .O(gate435inter3));
  inv1  gate705(.a(s_23), .O(gate435inter4));
  nand2 gate706(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate707(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate708(.a(G9), .O(gate435inter7));
  inv1  gate709(.a(G1156), .O(gate435inter8));
  nand2 gate710(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate711(.a(s_23), .b(gate435inter3), .O(gate435inter10));
  nor2  gate712(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate713(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate714(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate617(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate618(.a(gate438inter0), .b(s_10), .O(gate438inter1));
  and2  gate619(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate620(.a(s_10), .O(gate438inter3));
  inv1  gate621(.a(s_11), .O(gate438inter4));
  nand2 gate622(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate623(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate624(.a(G1063), .O(gate438inter7));
  inv1  gate625(.a(G1159), .O(gate438inter8));
  nand2 gate626(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate627(.a(s_11), .b(gate438inter3), .O(gate438inter10));
  nor2  gate628(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate629(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate630(.a(gate438inter12), .b(gate438inter1), .O(G1247));

  xor2  gate1261(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate1262(.a(gate439inter0), .b(s_102), .O(gate439inter1));
  and2  gate1263(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate1264(.a(s_102), .O(gate439inter3));
  inv1  gate1265(.a(s_103), .O(gate439inter4));
  nand2 gate1266(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate1267(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate1268(.a(G11), .O(gate439inter7));
  inv1  gate1269(.a(G1162), .O(gate439inter8));
  nand2 gate1270(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate1271(.a(s_103), .b(gate439inter3), .O(gate439inter10));
  nor2  gate1272(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate1273(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate1274(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate1233(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate1234(.a(gate442inter0), .b(s_98), .O(gate442inter1));
  and2  gate1235(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate1236(.a(s_98), .O(gate442inter3));
  inv1  gate1237(.a(s_99), .O(gate442inter4));
  nand2 gate1238(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate1239(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate1240(.a(G1069), .O(gate442inter7));
  inv1  gate1241(.a(G1165), .O(gate442inter8));
  nand2 gate1242(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate1243(.a(s_99), .b(gate442inter3), .O(gate442inter10));
  nor2  gate1244(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate1245(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate1246(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate2045(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate2046(.a(gate444inter0), .b(s_214), .O(gate444inter1));
  and2  gate2047(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate2048(.a(s_214), .O(gate444inter3));
  inv1  gate2049(.a(s_215), .O(gate444inter4));
  nand2 gate2050(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate2051(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate2052(.a(G1072), .O(gate444inter7));
  inv1  gate2053(.a(G1168), .O(gate444inter8));
  nand2 gate2054(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate2055(.a(s_215), .b(gate444inter3), .O(gate444inter10));
  nor2  gate2056(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate2057(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate2058(.a(gate444inter12), .b(gate444inter1), .O(G1253));

  xor2  gate1961(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate1962(.a(gate445inter0), .b(s_202), .O(gate445inter1));
  and2  gate1963(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate1964(.a(s_202), .O(gate445inter3));
  inv1  gate1965(.a(s_203), .O(gate445inter4));
  nand2 gate1966(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate1967(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate1968(.a(G14), .O(gate445inter7));
  inv1  gate1969(.a(G1171), .O(gate445inter8));
  nand2 gate1970(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate1971(.a(s_203), .b(gate445inter3), .O(gate445inter10));
  nor2  gate1972(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate1973(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate1974(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );

  xor2  gate1947(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate1948(.a(gate447inter0), .b(s_200), .O(gate447inter1));
  and2  gate1949(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate1950(.a(s_200), .O(gate447inter3));
  inv1  gate1951(.a(s_201), .O(gate447inter4));
  nand2 gate1952(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate1953(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate1954(.a(G15), .O(gate447inter7));
  inv1  gate1955(.a(G1174), .O(gate447inter8));
  nand2 gate1956(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate1957(.a(s_201), .b(gate447inter3), .O(gate447inter10));
  nor2  gate1958(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate1959(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate1960(.a(gate447inter12), .b(gate447inter1), .O(G1256));

  xor2  gate2087(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate2088(.a(gate448inter0), .b(s_220), .O(gate448inter1));
  and2  gate2089(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate2090(.a(s_220), .O(gate448inter3));
  inv1  gate2091(.a(s_221), .O(gate448inter4));
  nand2 gate2092(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate2093(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate2094(.a(G1078), .O(gate448inter7));
  inv1  gate2095(.a(G1174), .O(gate448inter8));
  nand2 gate2096(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate2097(.a(s_221), .b(gate448inter3), .O(gate448inter10));
  nor2  gate2098(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate2099(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate2100(.a(gate448inter12), .b(gate448inter1), .O(G1257));

  xor2  gate911(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate912(.a(gate449inter0), .b(s_52), .O(gate449inter1));
  and2  gate913(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate914(.a(s_52), .O(gate449inter3));
  inv1  gate915(.a(s_53), .O(gate449inter4));
  nand2 gate916(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate917(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate918(.a(G16), .O(gate449inter7));
  inv1  gate919(.a(G1177), .O(gate449inter8));
  nand2 gate920(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate921(.a(s_53), .b(gate449inter3), .O(gate449inter10));
  nor2  gate922(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate923(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate924(.a(gate449inter12), .b(gate449inter1), .O(G1258));

  xor2  gate1555(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate1556(.a(gate450inter0), .b(s_144), .O(gate450inter1));
  and2  gate1557(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate1558(.a(s_144), .O(gate450inter3));
  inv1  gate1559(.a(s_145), .O(gate450inter4));
  nand2 gate1560(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate1561(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate1562(.a(G1081), .O(gate450inter7));
  inv1  gate1563(.a(G1177), .O(gate450inter8));
  nand2 gate1564(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate1565(.a(s_145), .b(gate450inter3), .O(gate450inter10));
  nor2  gate1566(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate1567(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate1568(.a(gate450inter12), .b(gate450inter1), .O(G1259));
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate1331(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate1332(.a(gate459inter0), .b(s_112), .O(gate459inter1));
  and2  gate1333(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate1334(.a(s_112), .O(gate459inter3));
  inv1  gate1335(.a(s_113), .O(gate459inter4));
  nand2 gate1336(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate1337(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate1338(.a(G21), .O(gate459inter7));
  inv1  gate1339(.a(G1192), .O(gate459inter8));
  nand2 gate1340(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate1341(.a(s_113), .b(gate459inter3), .O(gate459inter10));
  nor2  gate1342(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate1343(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate1344(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate2325(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate2326(.a(gate461inter0), .b(s_254), .O(gate461inter1));
  and2  gate2327(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate2328(.a(s_254), .O(gate461inter3));
  inv1  gate2329(.a(s_255), .O(gate461inter4));
  nand2 gate2330(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate2331(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate2332(.a(G22), .O(gate461inter7));
  inv1  gate2333(.a(G1195), .O(gate461inter8));
  nand2 gate2334(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate2335(.a(s_255), .b(gate461inter3), .O(gate461inter10));
  nor2  gate2336(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate2337(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate2338(.a(gate461inter12), .b(gate461inter1), .O(G1270));
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate1429(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate1430(.a(gate464inter0), .b(s_126), .O(gate464inter1));
  and2  gate1431(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate1432(.a(s_126), .O(gate464inter3));
  inv1  gate1433(.a(s_127), .O(gate464inter4));
  nand2 gate1434(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate1435(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate1436(.a(G1102), .O(gate464inter7));
  inv1  gate1437(.a(G1198), .O(gate464inter8));
  nand2 gate1438(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate1439(.a(s_127), .b(gate464inter3), .O(gate464inter10));
  nor2  gate1440(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate1441(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate1442(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate1793(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate1794(.a(gate467inter0), .b(s_178), .O(gate467inter1));
  and2  gate1795(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate1796(.a(s_178), .O(gate467inter3));
  inv1  gate1797(.a(s_179), .O(gate467inter4));
  nand2 gate1798(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate1799(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate1800(.a(G25), .O(gate467inter7));
  inv1  gate1801(.a(G1204), .O(gate467inter8));
  nand2 gate1802(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate1803(.a(s_179), .b(gate467inter3), .O(gate467inter10));
  nor2  gate1804(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate1805(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate1806(.a(gate467inter12), .b(gate467inter1), .O(G1276));

  xor2  gate645(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate646(.a(gate468inter0), .b(s_14), .O(gate468inter1));
  and2  gate647(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate648(.a(s_14), .O(gate468inter3));
  inv1  gate649(.a(s_15), .O(gate468inter4));
  nand2 gate650(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate651(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate652(.a(G1108), .O(gate468inter7));
  inv1  gate653(.a(G1204), .O(gate468inter8));
  nand2 gate654(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate655(.a(s_15), .b(gate468inter3), .O(gate468inter10));
  nor2  gate656(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate657(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate658(.a(gate468inter12), .b(gate468inter1), .O(G1277));

  xor2  gate995(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate996(.a(gate469inter0), .b(s_64), .O(gate469inter1));
  and2  gate997(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate998(.a(s_64), .O(gate469inter3));
  inv1  gate999(.a(s_65), .O(gate469inter4));
  nand2 gate1000(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate1001(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate1002(.a(G26), .O(gate469inter7));
  inv1  gate1003(.a(G1207), .O(gate469inter8));
  nand2 gate1004(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate1005(.a(s_65), .b(gate469inter3), .O(gate469inter10));
  nor2  gate1006(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate1007(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate1008(.a(gate469inter12), .b(gate469inter1), .O(G1278));
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate1709(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate1710(.a(gate477inter0), .b(s_166), .O(gate477inter1));
  and2  gate1711(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate1712(.a(s_166), .O(gate477inter3));
  inv1  gate1713(.a(s_167), .O(gate477inter4));
  nand2 gate1714(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate1715(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate1716(.a(G30), .O(gate477inter7));
  inv1  gate1717(.a(G1219), .O(gate477inter8));
  nand2 gate1718(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate1719(.a(s_167), .b(gate477inter3), .O(gate477inter10));
  nor2  gate1720(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate1721(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate1722(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate757(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate758(.a(gate482inter0), .b(s_30), .O(gate482inter1));
  and2  gate759(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate760(.a(s_30), .O(gate482inter3));
  inv1  gate761(.a(s_31), .O(gate482inter4));
  nand2 gate762(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate763(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate764(.a(G1129), .O(gate482inter7));
  inv1  gate765(.a(G1225), .O(gate482inter8));
  nand2 gate766(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate767(.a(s_31), .b(gate482inter3), .O(gate482inter10));
  nor2  gate768(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate769(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate770(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );

  xor2  gate1065(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate1066(.a(gate484inter0), .b(s_74), .O(gate484inter1));
  and2  gate1067(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate1068(.a(s_74), .O(gate484inter3));
  inv1  gate1069(.a(s_75), .O(gate484inter4));
  nand2 gate1070(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate1071(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate1072(.a(G1230), .O(gate484inter7));
  inv1  gate1073(.a(G1231), .O(gate484inter8));
  nand2 gate1074(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate1075(.a(s_75), .b(gate484inter3), .O(gate484inter10));
  nor2  gate1076(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate1077(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate1078(.a(gate484inter12), .b(gate484inter1), .O(G1293));

  xor2  gate1009(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate1010(.a(gate485inter0), .b(s_66), .O(gate485inter1));
  and2  gate1011(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate1012(.a(s_66), .O(gate485inter3));
  inv1  gate1013(.a(s_67), .O(gate485inter4));
  nand2 gate1014(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate1015(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate1016(.a(G1232), .O(gate485inter7));
  inv1  gate1017(.a(G1233), .O(gate485inter8));
  nand2 gate1018(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate1019(.a(s_67), .b(gate485inter3), .O(gate485inter10));
  nor2  gate1020(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate1021(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate1022(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate659(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate660(.a(gate488inter0), .b(s_16), .O(gate488inter1));
  and2  gate661(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate662(.a(s_16), .O(gate488inter3));
  inv1  gate663(.a(s_17), .O(gate488inter4));
  nand2 gate664(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate665(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate666(.a(G1238), .O(gate488inter7));
  inv1  gate667(.a(G1239), .O(gate488inter8));
  nand2 gate668(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate669(.a(s_17), .b(gate488inter3), .O(gate488inter10));
  nor2  gate670(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate671(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate672(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate2185(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate2186(.a(gate491inter0), .b(s_234), .O(gate491inter1));
  and2  gate2187(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate2188(.a(s_234), .O(gate491inter3));
  inv1  gate2189(.a(s_235), .O(gate491inter4));
  nand2 gate2190(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate2191(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate2192(.a(G1244), .O(gate491inter7));
  inv1  gate2193(.a(G1245), .O(gate491inter8));
  nand2 gate2194(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate2195(.a(s_235), .b(gate491inter3), .O(gate491inter10));
  nor2  gate2196(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate2197(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate2198(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate1247(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1248(.a(gate494inter0), .b(s_100), .O(gate494inter1));
  and2  gate1249(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1250(.a(s_100), .O(gate494inter3));
  inv1  gate1251(.a(s_101), .O(gate494inter4));
  nand2 gate1252(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1253(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1254(.a(G1250), .O(gate494inter7));
  inv1  gate1255(.a(G1251), .O(gate494inter8));
  nand2 gate1256(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1257(.a(s_101), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1258(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1259(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1260(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate1051(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate1052(.a(gate496inter0), .b(s_72), .O(gate496inter1));
  and2  gate1053(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate1054(.a(s_72), .O(gate496inter3));
  inv1  gate1055(.a(s_73), .O(gate496inter4));
  nand2 gate1056(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate1057(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate1058(.a(G1254), .O(gate496inter7));
  inv1  gate1059(.a(G1255), .O(gate496inter8));
  nand2 gate1060(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate1061(.a(s_73), .b(gate496inter3), .O(gate496inter10));
  nor2  gate1062(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate1063(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate1064(.a(gate496inter12), .b(gate496inter1), .O(G1305));

  xor2  gate1653(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate1654(.a(gate497inter0), .b(s_158), .O(gate497inter1));
  and2  gate1655(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate1656(.a(s_158), .O(gate497inter3));
  inv1  gate1657(.a(s_159), .O(gate497inter4));
  nand2 gate1658(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate1659(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate1660(.a(G1256), .O(gate497inter7));
  inv1  gate1661(.a(G1257), .O(gate497inter8));
  nand2 gate1662(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate1663(.a(s_159), .b(gate497inter3), .O(gate497inter10));
  nor2  gate1664(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate1665(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate1666(.a(gate497inter12), .b(gate497inter1), .O(G1306));

  xor2  gate1303(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate1304(.a(gate498inter0), .b(s_108), .O(gate498inter1));
  and2  gate1305(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate1306(.a(s_108), .O(gate498inter3));
  inv1  gate1307(.a(s_109), .O(gate498inter4));
  nand2 gate1308(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate1309(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate1310(.a(G1258), .O(gate498inter7));
  inv1  gate1311(.a(G1259), .O(gate498inter8));
  nand2 gate1312(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate1313(.a(s_109), .b(gate498inter3), .O(gate498inter10));
  nor2  gate1314(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate1315(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate1316(.a(gate498inter12), .b(gate498inter1), .O(G1307));

  xor2  gate1457(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate1458(.a(gate499inter0), .b(s_130), .O(gate499inter1));
  and2  gate1459(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate1460(.a(s_130), .O(gate499inter3));
  inv1  gate1461(.a(s_131), .O(gate499inter4));
  nand2 gate1462(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate1463(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate1464(.a(G1260), .O(gate499inter7));
  inv1  gate1465(.a(G1261), .O(gate499inter8));
  nand2 gate1466(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate1467(.a(s_131), .b(gate499inter3), .O(gate499inter10));
  nor2  gate1468(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate1469(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate1470(.a(gate499inter12), .b(gate499inter1), .O(G1308));

  xor2  gate575(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate576(.a(gate500inter0), .b(s_4), .O(gate500inter1));
  and2  gate577(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate578(.a(s_4), .O(gate500inter3));
  inv1  gate579(.a(s_5), .O(gate500inter4));
  nand2 gate580(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate581(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate582(.a(G1262), .O(gate500inter7));
  inv1  gate583(.a(G1263), .O(gate500inter8));
  nand2 gate584(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate585(.a(s_5), .b(gate500inter3), .O(gate500inter10));
  nor2  gate586(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate587(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate588(.a(gate500inter12), .b(gate500inter1), .O(G1309));
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );

  xor2  gate715(.a(G1267), .b(G1266), .O(gate502inter0));
  nand2 gate716(.a(gate502inter0), .b(s_24), .O(gate502inter1));
  and2  gate717(.a(G1267), .b(G1266), .O(gate502inter2));
  inv1  gate718(.a(s_24), .O(gate502inter3));
  inv1  gate719(.a(s_25), .O(gate502inter4));
  nand2 gate720(.a(gate502inter4), .b(gate502inter3), .O(gate502inter5));
  nor2  gate721(.a(gate502inter5), .b(gate502inter2), .O(gate502inter6));
  inv1  gate722(.a(G1266), .O(gate502inter7));
  inv1  gate723(.a(G1267), .O(gate502inter8));
  nand2 gate724(.a(gate502inter8), .b(gate502inter7), .O(gate502inter9));
  nand2 gate725(.a(s_25), .b(gate502inter3), .O(gate502inter10));
  nor2  gate726(.a(gate502inter10), .b(gate502inter9), .O(gate502inter11));
  nor2  gate727(.a(gate502inter11), .b(gate502inter6), .O(gate502inter12));
  nand2 gate728(.a(gate502inter12), .b(gate502inter1), .O(G1311));
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate2311(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate2312(.a(gate510inter0), .b(s_252), .O(gate510inter1));
  and2  gate2313(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate2314(.a(s_252), .O(gate510inter3));
  inv1  gate2315(.a(s_253), .O(gate510inter4));
  nand2 gate2316(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate2317(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate2318(.a(G1282), .O(gate510inter7));
  inv1  gate2319(.a(G1283), .O(gate510inter8));
  nand2 gate2320(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate2321(.a(s_253), .b(gate510inter3), .O(gate510inter10));
  nor2  gate2322(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate2323(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate2324(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate1401(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate1402(.a(gate514inter0), .b(s_122), .O(gate514inter1));
  and2  gate1403(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate1404(.a(s_122), .O(gate514inter3));
  inv1  gate1405(.a(s_123), .O(gate514inter4));
  nand2 gate1406(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate1407(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate1408(.a(G1290), .O(gate514inter7));
  inv1  gate1409(.a(G1291), .O(gate514inter8));
  nand2 gate1410(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate1411(.a(s_123), .b(gate514inter3), .O(gate514inter10));
  nor2  gate1412(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate1413(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate1414(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule