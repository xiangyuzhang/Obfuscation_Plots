module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate911(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate912(.a(gate12inter0), .b(s_52), .O(gate12inter1));
  and2  gate913(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate914(.a(s_52), .O(gate12inter3));
  inv1  gate915(.a(s_53), .O(gate12inter4));
  nand2 gate916(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate917(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate918(.a(G7), .O(gate12inter7));
  inv1  gate919(.a(G8), .O(gate12inter8));
  nand2 gate920(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate921(.a(s_53), .b(gate12inter3), .O(gate12inter10));
  nor2  gate922(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate923(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate924(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate1247(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate1248(.a(gate26inter0), .b(s_100), .O(gate26inter1));
  and2  gate1249(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate1250(.a(s_100), .O(gate26inter3));
  inv1  gate1251(.a(s_101), .O(gate26inter4));
  nand2 gate1252(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate1253(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate1254(.a(G9), .O(gate26inter7));
  inv1  gate1255(.a(G13), .O(gate26inter8));
  nand2 gate1256(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate1257(.a(s_101), .b(gate26inter3), .O(gate26inter10));
  nor2  gate1258(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate1259(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate1260(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate1373(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate1374(.a(gate34inter0), .b(s_118), .O(gate34inter1));
  and2  gate1375(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate1376(.a(s_118), .O(gate34inter3));
  inv1  gate1377(.a(s_119), .O(gate34inter4));
  nand2 gate1378(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate1379(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate1380(.a(G25), .O(gate34inter7));
  inv1  gate1381(.a(G29), .O(gate34inter8));
  nand2 gate1382(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate1383(.a(s_119), .b(gate34inter3), .O(gate34inter10));
  nor2  gate1384(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate1385(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate1386(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate967(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate968(.a(gate43inter0), .b(s_60), .O(gate43inter1));
  and2  gate969(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate970(.a(s_60), .O(gate43inter3));
  inv1  gate971(.a(s_61), .O(gate43inter4));
  nand2 gate972(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate973(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate974(.a(G3), .O(gate43inter7));
  inv1  gate975(.a(G269), .O(gate43inter8));
  nand2 gate976(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate977(.a(s_61), .b(gate43inter3), .O(gate43inter10));
  nor2  gate978(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate979(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate980(.a(gate43inter12), .b(gate43inter1), .O(G364));

  xor2  gate1289(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate1290(.a(gate44inter0), .b(s_106), .O(gate44inter1));
  and2  gate1291(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate1292(.a(s_106), .O(gate44inter3));
  inv1  gate1293(.a(s_107), .O(gate44inter4));
  nand2 gate1294(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate1295(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate1296(.a(G4), .O(gate44inter7));
  inv1  gate1297(.a(G269), .O(gate44inter8));
  nand2 gate1298(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate1299(.a(s_107), .b(gate44inter3), .O(gate44inter10));
  nor2  gate1300(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate1301(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate1302(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate1163(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate1164(.a(gate54inter0), .b(s_88), .O(gate54inter1));
  and2  gate1165(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate1166(.a(s_88), .O(gate54inter3));
  inv1  gate1167(.a(s_89), .O(gate54inter4));
  nand2 gate1168(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate1169(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate1170(.a(G14), .O(gate54inter7));
  inv1  gate1171(.a(G284), .O(gate54inter8));
  nand2 gate1172(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate1173(.a(s_89), .b(gate54inter3), .O(gate54inter10));
  nor2  gate1174(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate1175(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate1176(.a(gate54inter12), .b(gate54inter1), .O(G375));

  xor2  gate1065(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate1066(.a(gate55inter0), .b(s_74), .O(gate55inter1));
  and2  gate1067(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate1068(.a(s_74), .O(gate55inter3));
  inv1  gate1069(.a(s_75), .O(gate55inter4));
  nand2 gate1070(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate1071(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate1072(.a(G15), .O(gate55inter7));
  inv1  gate1073(.a(G287), .O(gate55inter8));
  nand2 gate1074(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate1075(.a(s_75), .b(gate55inter3), .O(gate55inter10));
  nor2  gate1076(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate1077(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate1078(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate1261(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate1262(.a(gate66inter0), .b(s_102), .O(gate66inter1));
  and2  gate1263(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate1264(.a(s_102), .O(gate66inter3));
  inv1  gate1265(.a(s_103), .O(gate66inter4));
  nand2 gate1266(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate1267(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate1268(.a(G26), .O(gate66inter7));
  inv1  gate1269(.a(G302), .O(gate66inter8));
  nand2 gate1270(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate1271(.a(s_103), .b(gate66inter3), .O(gate66inter10));
  nor2  gate1272(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate1273(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate1274(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate855(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate856(.a(gate74inter0), .b(s_44), .O(gate74inter1));
  and2  gate857(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate858(.a(s_44), .O(gate74inter3));
  inv1  gate859(.a(s_45), .O(gate74inter4));
  nand2 gate860(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate861(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate862(.a(G5), .O(gate74inter7));
  inv1  gate863(.a(G314), .O(gate74inter8));
  nand2 gate864(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate865(.a(s_45), .b(gate74inter3), .O(gate74inter10));
  nor2  gate866(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate867(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate868(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate1135(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate1136(.a(gate77inter0), .b(s_84), .O(gate77inter1));
  and2  gate1137(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate1138(.a(s_84), .O(gate77inter3));
  inv1  gate1139(.a(s_85), .O(gate77inter4));
  nand2 gate1140(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate1141(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate1142(.a(G2), .O(gate77inter7));
  inv1  gate1143(.a(G320), .O(gate77inter8));
  nand2 gate1144(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate1145(.a(s_85), .b(gate77inter3), .O(gate77inter10));
  nor2  gate1146(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate1147(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate1148(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );

  xor2  gate561(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate562(.a(gate84inter0), .b(s_2), .O(gate84inter1));
  and2  gate563(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate564(.a(s_2), .O(gate84inter3));
  inv1  gate565(.a(s_3), .O(gate84inter4));
  nand2 gate566(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate567(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate568(.a(G15), .O(gate84inter7));
  inv1  gate569(.a(G329), .O(gate84inter8));
  nand2 gate570(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate571(.a(s_3), .b(gate84inter3), .O(gate84inter10));
  nor2  gate572(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate573(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate574(.a(gate84inter12), .b(gate84inter1), .O(G405));
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate1149(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate1150(.a(gate90inter0), .b(s_86), .O(gate90inter1));
  and2  gate1151(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate1152(.a(s_86), .O(gate90inter3));
  inv1  gate1153(.a(s_87), .O(gate90inter4));
  nand2 gate1154(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate1155(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate1156(.a(G21), .O(gate90inter7));
  inv1  gate1157(.a(G338), .O(gate90inter8));
  nand2 gate1158(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate1159(.a(s_87), .b(gate90inter3), .O(gate90inter10));
  nor2  gate1160(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate1161(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate1162(.a(gate90inter12), .b(gate90inter1), .O(G411));
nand2 gate91( .a(G25), .b(G341), .O(G412) );

  xor2  gate1317(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate1318(.a(gate92inter0), .b(s_110), .O(gate92inter1));
  and2  gate1319(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate1320(.a(s_110), .O(gate92inter3));
  inv1  gate1321(.a(s_111), .O(gate92inter4));
  nand2 gate1322(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate1323(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate1324(.a(G29), .O(gate92inter7));
  inv1  gate1325(.a(G341), .O(gate92inter8));
  nand2 gate1326(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate1327(.a(s_111), .b(gate92inter3), .O(gate92inter10));
  nor2  gate1328(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate1329(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate1330(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );

  xor2  gate1345(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate1346(.a(gate101inter0), .b(s_114), .O(gate101inter1));
  and2  gate1347(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate1348(.a(s_114), .O(gate101inter3));
  inv1  gate1349(.a(s_115), .O(gate101inter4));
  nand2 gate1350(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate1351(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate1352(.a(G20), .O(gate101inter7));
  inv1  gate1353(.a(G356), .O(gate101inter8));
  nand2 gate1354(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate1355(.a(s_115), .b(gate101inter3), .O(gate101inter10));
  nor2  gate1356(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate1357(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate1358(.a(gate101inter12), .b(gate101inter1), .O(G422));
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate687(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate688(.a(gate106inter0), .b(s_20), .O(gate106inter1));
  and2  gate689(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate690(.a(s_20), .O(gate106inter3));
  inv1  gate691(.a(s_21), .O(gate106inter4));
  nand2 gate692(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate693(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate694(.a(G364), .O(gate106inter7));
  inv1  gate695(.a(G365), .O(gate106inter8));
  nand2 gate696(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate697(.a(s_21), .b(gate106inter3), .O(gate106inter10));
  nor2  gate698(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate699(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate700(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );

  xor2  gate1219(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate1220(.a(gate111inter0), .b(s_96), .O(gate111inter1));
  and2  gate1221(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate1222(.a(s_96), .O(gate111inter3));
  inv1  gate1223(.a(s_97), .O(gate111inter4));
  nand2 gate1224(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate1225(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate1226(.a(G374), .O(gate111inter7));
  inv1  gate1227(.a(G375), .O(gate111inter8));
  nand2 gate1228(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate1229(.a(s_97), .b(gate111inter3), .O(gate111inter10));
  nor2  gate1230(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate1231(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate1232(.a(gate111inter12), .b(gate111inter1), .O(G444));
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );

  xor2  gate1401(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate1402(.a(gate114inter0), .b(s_122), .O(gate114inter1));
  and2  gate1403(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate1404(.a(s_122), .O(gate114inter3));
  inv1  gate1405(.a(s_123), .O(gate114inter4));
  nand2 gate1406(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate1407(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate1408(.a(G380), .O(gate114inter7));
  inv1  gate1409(.a(G381), .O(gate114inter8));
  nand2 gate1410(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate1411(.a(s_123), .b(gate114inter3), .O(gate114inter10));
  nor2  gate1412(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate1413(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate1414(.a(gate114inter12), .b(gate114inter1), .O(G453));
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate827(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate828(.a(gate118inter0), .b(s_40), .O(gate118inter1));
  and2  gate829(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate830(.a(s_40), .O(gate118inter3));
  inv1  gate831(.a(s_41), .O(gate118inter4));
  nand2 gate832(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate833(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate834(.a(G388), .O(gate118inter7));
  inv1  gate835(.a(G389), .O(gate118inter8));
  nand2 gate836(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate837(.a(s_41), .b(gate118inter3), .O(gate118inter10));
  nor2  gate838(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate839(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate840(.a(gate118inter12), .b(gate118inter1), .O(G465));
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );

  xor2  gate1009(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate1010(.a(gate122inter0), .b(s_66), .O(gate122inter1));
  and2  gate1011(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate1012(.a(s_66), .O(gate122inter3));
  inv1  gate1013(.a(s_67), .O(gate122inter4));
  nand2 gate1014(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate1015(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate1016(.a(G396), .O(gate122inter7));
  inv1  gate1017(.a(G397), .O(gate122inter8));
  nand2 gate1018(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate1019(.a(s_67), .b(gate122inter3), .O(gate122inter10));
  nor2  gate1020(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate1021(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate1022(.a(gate122inter12), .b(gate122inter1), .O(G477));
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate813(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate814(.a(gate136inter0), .b(s_38), .O(gate136inter1));
  and2  gate815(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate816(.a(s_38), .O(gate136inter3));
  inv1  gate817(.a(s_39), .O(gate136inter4));
  nand2 gate818(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate819(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate820(.a(G424), .O(gate136inter7));
  inv1  gate821(.a(G425), .O(gate136inter8));
  nand2 gate822(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate823(.a(s_39), .b(gate136inter3), .O(gate136inter10));
  nor2  gate824(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate825(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate826(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );

  xor2  gate1303(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate1304(.a(gate139inter0), .b(s_108), .O(gate139inter1));
  and2  gate1305(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate1306(.a(s_108), .O(gate139inter3));
  inv1  gate1307(.a(s_109), .O(gate139inter4));
  nand2 gate1308(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate1309(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate1310(.a(G438), .O(gate139inter7));
  inv1  gate1311(.a(G441), .O(gate139inter8));
  nand2 gate1312(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate1313(.a(s_109), .b(gate139inter3), .O(gate139inter10));
  nor2  gate1314(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate1315(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate1316(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate1331(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1332(.a(gate148inter0), .b(s_112), .O(gate148inter1));
  and2  gate1333(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1334(.a(s_112), .O(gate148inter3));
  inv1  gate1335(.a(s_113), .O(gate148inter4));
  nand2 gate1336(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1337(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1338(.a(G492), .O(gate148inter7));
  inv1  gate1339(.a(G495), .O(gate148inter8));
  nand2 gate1340(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1341(.a(s_113), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1342(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1343(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1344(.a(gate148inter12), .b(gate148inter1), .O(G555));

  xor2  gate799(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate800(.a(gate149inter0), .b(s_36), .O(gate149inter1));
  and2  gate801(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate802(.a(s_36), .O(gate149inter3));
  inv1  gate803(.a(s_37), .O(gate149inter4));
  nand2 gate804(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate805(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate806(.a(G498), .O(gate149inter7));
  inv1  gate807(.a(G501), .O(gate149inter8));
  nand2 gate808(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate809(.a(s_37), .b(gate149inter3), .O(gate149inter10));
  nor2  gate810(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate811(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate812(.a(gate149inter12), .b(gate149inter1), .O(G558));

  xor2  gate995(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate996(.a(gate150inter0), .b(s_64), .O(gate150inter1));
  and2  gate997(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate998(.a(s_64), .O(gate150inter3));
  inv1  gate999(.a(s_65), .O(gate150inter4));
  nand2 gate1000(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate1001(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate1002(.a(G504), .O(gate150inter7));
  inv1  gate1003(.a(G507), .O(gate150inter8));
  nand2 gate1004(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate1005(.a(s_65), .b(gate150inter3), .O(gate150inter10));
  nor2  gate1006(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate1007(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate1008(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );

  xor2  gate785(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate786(.a(gate158inter0), .b(s_34), .O(gate158inter1));
  and2  gate787(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate788(.a(s_34), .O(gate158inter3));
  inv1  gate789(.a(s_35), .O(gate158inter4));
  nand2 gate790(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate791(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate792(.a(G441), .O(gate158inter7));
  inv1  gate793(.a(G528), .O(gate158inter8));
  nand2 gate794(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate795(.a(s_35), .b(gate158inter3), .O(gate158inter10));
  nor2  gate796(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate797(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate798(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate869(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate870(.a(gate162inter0), .b(s_46), .O(gate162inter1));
  and2  gate871(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate872(.a(s_46), .O(gate162inter3));
  inv1  gate873(.a(s_47), .O(gate162inter4));
  nand2 gate874(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate875(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate876(.a(G453), .O(gate162inter7));
  inv1  gate877(.a(G534), .O(gate162inter8));
  nand2 gate878(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate879(.a(s_47), .b(gate162inter3), .O(gate162inter10));
  nor2  gate880(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate881(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate882(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );

  xor2  gate645(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate646(.a(gate166inter0), .b(s_14), .O(gate166inter1));
  and2  gate647(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate648(.a(s_14), .O(gate166inter3));
  inv1  gate649(.a(s_15), .O(gate166inter4));
  nand2 gate650(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate651(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate652(.a(G465), .O(gate166inter7));
  inv1  gate653(.a(G540), .O(gate166inter8));
  nand2 gate654(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate655(.a(s_15), .b(gate166inter3), .O(gate166inter10));
  nor2  gate656(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate657(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate658(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );

  xor2  gate883(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate884(.a(gate169inter0), .b(s_48), .O(gate169inter1));
  and2  gate885(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate886(.a(s_48), .O(gate169inter3));
  inv1  gate887(.a(s_49), .O(gate169inter4));
  nand2 gate888(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate889(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate890(.a(G474), .O(gate169inter7));
  inv1  gate891(.a(G546), .O(gate169inter8));
  nand2 gate892(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate893(.a(s_49), .b(gate169inter3), .O(gate169inter10));
  nor2  gate894(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate895(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate896(.a(gate169inter12), .b(gate169inter1), .O(G586));
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate1429(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate1430(.a(gate174inter0), .b(s_126), .O(gate174inter1));
  and2  gate1431(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate1432(.a(s_126), .O(gate174inter3));
  inv1  gate1433(.a(s_127), .O(gate174inter4));
  nand2 gate1434(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate1435(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate1436(.a(G489), .O(gate174inter7));
  inv1  gate1437(.a(G552), .O(gate174inter8));
  nand2 gate1438(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate1439(.a(s_127), .b(gate174inter3), .O(gate174inter10));
  nor2  gate1440(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate1441(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate1442(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );

  xor2  gate1093(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate1094(.a(gate189inter0), .b(s_78), .O(gate189inter1));
  and2  gate1095(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate1096(.a(s_78), .O(gate189inter3));
  inv1  gate1097(.a(s_79), .O(gate189inter4));
  nand2 gate1098(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate1099(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate1100(.a(G578), .O(gate189inter7));
  inv1  gate1101(.a(G579), .O(gate189inter8));
  nand2 gate1102(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate1103(.a(s_79), .b(gate189inter3), .O(gate189inter10));
  nor2  gate1104(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate1105(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate1106(.a(gate189inter12), .b(gate189inter1), .O(G622));
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate841(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate842(.a(gate193inter0), .b(s_42), .O(gate193inter1));
  and2  gate843(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate844(.a(s_42), .O(gate193inter3));
  inv1  gate845(.a(s_43), .O(gate193inter4));
  nand2 gate846(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate847(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate848(.a(G586), .O(gate193inter7));
  inv1  gate849(.a(G587), .O(gate193inter8));
  nand2 gate850(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate851(.a(s_43), .b(gate193inter3), .O(gate193inter10));
  nor2  gate852(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate853(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate854(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate729(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate730(.a(gate195inter0), .b(s_26), .O(gate195inter1));
  and2  gate731(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate732(.a(s_26), .O(gate195inter3));
  inv1  gate733(.a(s_27), .O(gate195inter4));
  nand2 gate734(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate735(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate736(.a(G590), .O(gate195inter7));
  inv1  gate737(.a(G591), .O(gate195inter8));
  nand2 gate738(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate739(.a(s_27), .b(gate195inter3), .O(gate195inter10));
  nor2  gate740(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate741(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate742(.a(gate195inter12), .b(gate195inter1), .O(G648));

  xor2  gate589(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate590(.a(gate196inter0), .b(s_6), .O(gate196inter1));
  and2  gate591(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate592(.a(s_6), .O(gate196inter3));
  inv1  gate593(.a(s_7), .O(gate196inter4));
  nand2 gate594(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate595(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate596(.a(G592), .O(gate196inter7));
  inv1  gate597(.a(G593), .O(gate196inter8));
  nand2 gate598(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate599(.a(s_7), .b(gate196inter3), .O(gate196inter10));
  nor2  gate600(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate601(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate602(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate547(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate548(.a(gate203inter0), .b(s_0), .O(gate203inter1));
  and2  gate549(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate550(.a(s_0), .O(gate203inter3));
  inv1  gate551(.a(s_1), .O(gate203inter4));
  nand2 gate552(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate553(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate554(.a(G602), .O(gate203inter7));
  inv1  gate555(.a(G612), .O(gate203inter8));
  nand2 gate556(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate557(.a(s_1), .b(gate203inter3), .O(gate203inter10));
  nor2  gate558(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate559(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate560(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate659(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate660(.a(gate206inter0), .b(s_16), .O(gate206inter1));
  and2  gate661(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate662(.a(s_16), .O(gate206inter3));
  inv1  gate663(.a(s_17), .O(gate206inter4));
  nand2 gate664(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate665(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate666(.a(G632), .O(gate206inter7));
  inv1  gate667(.a(G637), .O(gate206inter8));
  nand2 gate668(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate669(.a(s_17), .b(gate206inter3), .O(gate206inter10));
  nor2  gate670(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate671(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate672(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );

  xor2  gate603(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate604(.a(gate210inter0), .b(s_8), .O(gate210inter1));
  and2  gate605(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate606(.a(s_8), .O(gate210inter3));
  inv1  gate607(.a(s_9), .O(gate210inter4));
  nand2 gate608(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate609(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate610(.a(G607), .O(gate210inter7));
  inv1  gate611(.a(G666), .O(gate210inter8));
  nand2 gate612(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate613(.a(s_9), .b(gate210inter3), .O(gate210inter10));
  nor2  gate614(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate615(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate616(.a(gate210inter12), .b(gate210inter1), .O(G691));
nand2 gate211( .a(G612), .b(G669), .O(G692) );

  xor2  gate575(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate576(.a(gate212inter0), .b(s_4), .O(gate212inter1));
  and2  gate577(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate578(.a(s_4), .O(gate212inter3));
  inv1  gate579(.a(s_5), .O(gate212inter4));
  nand2 gate580(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate581(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate582(.a(G617), .O(gate212inter7));
  inv1  gate583(.a(G669), .O(gate212inter8));
  nand2 gate584(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate585(.a(s_5), .b(gate212inter3), .O(gate212inter10));
  nor2  gate586(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate587(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate588(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate743(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate744(.a(gate216inter0), .b(s_28), .O(gate216inter1));
  and2  gate745(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate746(.a(s_28), .O(gate216inter3));
  inv1  gate747(.a(s_29), .O(gate216inter4));
  nand2 gate748(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate749(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate750(.a(G617), .O(gate216inter7));
  inv1  gate751(.a(G675), .O(gate216inter8));
  nand2 gate752(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate753(.a(s_29), .b(gate216inter3), .O(gate216inter10));
  nor2  gate754(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate755(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate756(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate1023(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate1024(.a(gate223inter0), .b(s_68), .O(gate223inter1));
  and2  gate1025(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate1026(.a(s_68), .O(gate223inter3));
  inv1  gate1027(.a(s_69), .O(gate223inter4));
  nand2 gate1028(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate1029(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate1030(.a(G627), .O(gate223inter7));
  inv1  gate1031(.a(G687), .O(gate223inter8));
  nand2 gate1032(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate1033(.a(s_69), .b(gate223inter3), .O(gate223inter10));
  nor2  gate1034(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate1035(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate1036(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );

  xor2  gate1121(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate1122(.a(gate238inter0), .b(s_82), .O(gate238inter1));
  and2  gate1123(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate1124(.a(s_82), .O(gate238inter3));
  inv1  gate1125(.a(s_83), .O(gate238inter4));
  nand2 gate1126(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate1127(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate1128(.a(G257), .O(gate238inter7));
  inv1  gate1129(.a(G709), .O(gate238inter8));
  nand2 gate1130(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate1131(.a(s_83), .b(gate238inter3), .O(gate238inter10));
  nor2  gate1132(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate1133(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate1134(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate1415(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate1416(.a(gate240inter0), .b(s_124), .O(gate240inter1));
  and2  gate1417(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate1418(.a(s_124), .O(gate240inter3));
  inv1  gate1419(.a(s_125), .O(gate240inter4));
  nand2 gate1420(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate1421(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate1422(.a(G263), .O(gate240inter7));
  inv1  gate1423(.a(G715), .O(gate240inter8));
  nand2 gate1424(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate1425(.a(s_125), .b(gate240inter3), .O(gate240inter10));
  nor2  gate1426(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate1427(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate1428(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );

  xor2  gate1443(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate1444(.a(gate246inter0), .b(s_128), .O(gate246inter1));
  and2  gate1445(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate1446(.a(s_128), .O(gate246inter3));
  inv1  gate1447(.a(s_129), .O(gate246inter4));
  nand2 gate1448(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate1449(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate1450(.a(G724), .O(gate246inter7));
  inv1  gate1451(.a(G736), .O(gate246inter8));
  nand2 gate1452(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate1453(.a(s_129), .b(gate246inter3), .O(gate246inter10));
  nor2  gate1454(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate1455(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate1456(.a(gate246inter12), .b(gate246inter1), .O(G759));
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate1275(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate1276(.a(gate250inter0), .b(s_104), .O(gate250inter1));
  and2  gate1277(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate1278(.a(s_104), .O(gate250inter3));
  inv1  gate1279(.a(s_105), .O(gate250inter4));
  nand2 gate1280(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate1281(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate1282(.a(G706), .O(gate250inter7));
  inv1  gate1283(.a(G742), .O(gate250inter8));
  nand2 gate1284(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate1285(.a(s_105), .b(gate250inter3), .O(gate250inter10));
  nor2  gate1286(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate1287(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate1288(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate1177(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate1178(.a(gate253inter0), .b(s_90), .O(gate253inter1));
  and2  gate1179(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate1180(.a(s_90), .O(gate253inter3));
  inv1  gate1181(.a(s_91), .O(gate253inter4));
  nand2 gate1182(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate1183(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate1184(.a(G260), .O(gate253inter7));
  inv1  gate1185(.a(G748), .O(gate253inter8));
  nand2 gate1186(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate1187(.a(s_91), .b(gate253inter3), .O(gate253inter10));
  nor2  gate1188(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate1189(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate1190(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate953(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate954(.a(gate263inter0), .b(s_58), .O(gate263inter1));
  and2  gate955(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate956(.a(s_58), .O(gate263inter3));
  inv1  gate957(.a(s_59), .O(gate263inter4));
  nand2 gate958(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate959(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate960(.a(G766), .O(gate263inter7));
  inv1  gate961(.a(G767), .O(gate263inter8));
  nand2 gate962(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate963(.a(s_59), .b(gate263inter3), .O(gate263inter10));
  nor2  gate964(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate965(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate966(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate897(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate898(.a(gate276inter0), .b(s_50), .O(gate276inter1));
  and2  gate899(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate900(.a(s_50), .O(gate276inter3));
  inv1  gate901(.a(s_51), .O(gate276inter4));
  nand2 gate902(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate903(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate904(.a(G773), .O(gate276inter7));
  inv1  gate905(.a(G797), .O(gate276inter8));
  nand2 gate906(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate907(.a(s_51), .b(gate276inter3), .O(gate276inter10));
  nor2  gate908(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate909(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate910(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );

  xor2  gate757(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate758(.a(gate281inter0), .b(s_30), .O(gate281inter1));
  and2  gate759(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate760(.a(s_30), .O(gate281inter3));
  inv1  gate761(.a(s_31), .O(gate281inter4));
  nand2 gate762(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate763(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate764(.a(G654), .O(gate281inter7));
  inv1  gate765(.a(G806), .O(gate281inter8));
  nand2 gate766(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate767(.a(s_31), .b(gate281inter3), .O(gate281inter10));
  nor2  gate768(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate769(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate770(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate1191(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate1192(.a(gate285inter0), .b(s_92), .O(gate285inter1));
  and2  gate1193(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate1194(.a(s_92), .O(gate285inter3));
  inv1  gate1195(.a(s_93), .O(gate285inter4));
  nand2 gate1196(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate1197(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate1198(.a(G660), .O(gate285inter7));
  inv1  gate1199(.a(G812), .O(gate285inter8));
  nand2 gate1200(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate1201(.a(s_93), .b(gate285inter3), .O(gate285inter10));
  nor2  gate1202(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate1203(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate1204(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate1457(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate1458(.a(gate287inter0), .b(s_130), .O(gate287inter1));
  and2  gate1459(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate1460(.a(s_130), .O(gate287inter3));
  inv1  gate1461(.a(s_131), .O(gate287inter4));
  nand2 gate1462(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate1463(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate1464(.a(G663), .O(gate287inter7));
  inv1  gate1465(.a(G815), .O(gate287inter8));
  nand2 gate1466(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate1467(.a(s_131), .b(gate287inter3), .O(gate287inter10));
  nor2  gate1468(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate1469(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate1470(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate715(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate716(.a(gate391inter0), .b(s_24), .O(gate391inter1));
  and2  gate717(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate718(.a(s_24), .O(gate391inter3));
  inv1  gate719(.a(s_25), .O(gate391inter4));
  nand2 gate720(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate721(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate722(.a(G5), .O(gate391inter7));
  inv1  gate723(.a(G1048), .O(gate391inter8));
  nand2 gate724(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate725(.a(s_25), .b(gate391inter3), .O(gate391inter10));
  nor2  gate726(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate727(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate728(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate1079(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1080(.a(gate395inter0), .b(s_76), .O(gate395inter1));
  and2  gate1081(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1082(.a(s_76), .O(gate395inter3));
  inv1  gate1083(.a(s_77), .O(gate395inter4));
  nand2 gate1084(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1085(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1086(.a(G9), .O(gate395inter7));
  inv1  gate1087(.a(G1060), .O(gate395inter8));
  nand2 gate1088(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1089(.a(s_77), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1090(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1091(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1092(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate925(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate926(.a(gate398inter0), .b(s_54), .O(gate398inter1));
  and2  gate927(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate928(.a(s_54), .O(gate398inter3));
  inv1  gate929(.a(s_55), .O(gate398inter4));
  nand2 gate930(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate931(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate932(.a(G12), .O(gate398inter7));
  inv1  gate933(.a(G1069), .O(gate398inter8));
  nand2 gate934(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate935(.a(s_55), .b(gate398inter3), .O(gate398inter10));
  nor2  gate936(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate937(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate938(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate1205(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate1206(.a(gate411inter0), .b(s_94), .O(gate411inter1));
  and2  gate1207(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate1208(.a(s_94), .O(gate411inter3));
  inv1  gate1209(.a(s_95), .O(gate411inter4));
  nand2 gate1210(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate1211(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate1212(.a(G25), .O(gate411inter7));
  inv1  gate1213(.a(G1108), .O(gate411inter8));
  nand2 gate1214(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate1215(.a(s_95), .b(gate411inter3), .O(gate411inter10));
  nor2  gate1216(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate1217(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate1218(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );

  xor2  gate1387(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate1388(.a(gate426inter0), .b(s_120), .O(gate426inter1));
  and2  gate1389(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate1390(.a(s_120), .O(gate426inter3));
  inv1  gate1391(.a(s_121), .O(gate426inter4));
  nand2 gate1392(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate1393(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate1394(.a(G1045), .O(gate426inter7));
  inv1  gate1395(.a(G1141), .O(gate426inter8));
  nand2 gate1396(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate1397(.a(s_121), .b(gate426inter3), .O(gate426inter10));
  nor2  gate1398(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate1399(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate1400(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate981(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate982(.a(gate433inter0), .b(s_62), .O(gate433inter1));
  and2  gate983(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate984(.a(s_62), .O(gate433inter3));
  inv1  gate985(.a(s_63), .O(gate433inter4));
  nand2 gate986(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate987(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate988(.a(G8), .O(gate433inter7));
  inv1  gate989(.a(G1153), .O(gate433inter8));
  nand2 gate990(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate991(.a(s_63), .b(gate433inter3), .O(gate433inter10));
  nor2  gate992(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate993(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate994(.a(gate433inter12), .b(gate433inter1), .O(G1242));

  xor2  gate771(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate772(.a(gate434inter0), .b(s_32), .O(gate434inter1));
  and2  gate773(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate774(.a(s_32), .O(gate434inter3));
  inv1  gate775(.a(s_33), .O(gate434inter4));
  nand2 gate776(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate777(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate778(.a(G1057), .O(gate434inter7));
  inv1  gate779(.a(G1153), .O(gate434inter8));
  nand2 gate780(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate781(.a(s_33), .b(gate434inter3), .O(gate434inter10));
  nor2  gate782(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate783(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate784(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate673(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate674(.a(gate445inter0), .b(s_18), .O(gate445inter1));
  and2  gate675(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate676(.a(s_18), .O(gate445inter3));
  inv1  gate677(.a(s_19), .O(gate445inter4));
  nand2 gate678(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate679(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate680(.a(G14), .O(gate445inter7));
  inv1  gate681(.a(G1171), .O(gate445inter8));
  nand2 gate682(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate683(.a(s_19), .b(gate445inter3), .O(gate445inter10));
  nor2  gate684(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate685(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate686(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate1051(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate1052(.a(gate457inter0), .b(s_72), .O(gate457inter1));
  and2  gate1053(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate1054(.a(s_72), .O(gate457inter3));
  inv1  gate1055(.a(s_73), .O(gate457inter4));
  nand2 gate1056(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate1057(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate1058(.a(G20), .O(gate457inter7));
  inv1  gate1059(.a(G1189), .O(gate457inter8));
  nand2 gate1060(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate1061(.a(s_73), .b(gate457inter3), .O(gate457inter10));
  nor2  gate1062(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate1063(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate1064(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate1233(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate1234(.a(gate472inter0), .b(s_98), .O(gate472inter1));
  and2  gate1235(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate1236(.a(s_98), .O(gate472inter3));
  inv1  gate1237(.a(s_99), .O(gate472inter4));
  nand2 gate1238(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate1239(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate1240(.a(G1114), .O(gate472inter7));
  inv1  gate1241(.a(G1210), .O(gate472inter8));
  nand2 gate1242(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate1243(.a(s_99), .b(gate472inter3), .O(gate472inter10));
  nor2  gate1244(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate1245(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate1246(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate1107(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate1108(.a(gate493inter0), .b(s_80), .O(gate493inter1));
  and2  gate1109(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate1110(.a(s_80), .O(gate493inter3));
  inv1  gate1111(.a(s_81), .O(gate493inter4));
  nand2 gate1112(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate1113(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate1114(.a(G1248), .O(gate493inter7));
  inv1  gate1115(.a(G1249), .O(gate493inter8));
  nand2 gate1116(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate1117(.a(s_81), .b(gate493inter3), .O(gate493inter10));
  nor2  gate1118(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate1119(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate1120(.a(gate493inter12), .b(gate493inter1), .O(G1302));
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate631(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate632(.a(gate501inter0), .b(s_12), .O(gate501inter1));
  and2  gate633(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate634(.a(s_12), .O(gate501inter3));
  inv1  gate635(.a(s_13), .O(gate501inter4));
  nand2 gate636(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate637(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate638(.a(G1264), .O(gate501inter7));
  inv1  gate639(.a(G1265), .O(gate501inter8));
  nand2 gate640(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate641(.a(s_13), .b(gate501inter3), .O(gate501inter10));
  nor2  gate642(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate643(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate644(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );

  xor2  gate617(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate618(.a(gate505inter0), .b(s_10), .O(gate505inter1));
  and2  gate619(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate620(.a(s_10), .O(gate505inter3));
  inv1  gate621(.a(s_11), .O(gate505inter4));
  nand2 gate622(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate623(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate624(.a(G1272), .O(gate505inter7));
  inv1  gate625(.a(G1273), .O(gate505inter8));
  nand2 gate626(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate627(.a(s_11), .b(gate505inter3), .O(gate505inter10));
  nor2  gate628(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate629(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate630(.a(gate505inter12), .b(gate505inter1), .O(G1314));
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate939(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate940(.a(gate508inter0), .b(s_56), .O(gate508inter1));
  and2  gate941(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate942(.a(s_56), .O(gate508inter3));
  inv1  gate943(.a(s_57), .O(gate508inter4));
  nand2 gate944(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate945(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate946(.a(G1278), .O(gate508inter7));
  inv1  gate947(.a(G1279), .O(gate508inter8));
  nand2 gate948(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate949(.a(s_57), .b(gate508inter3), .O(gate508inter10));
  nor2  gate950(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate951(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate952(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate1359(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate1360(.a(gate510inter0), .b(s_116), .O(gate510inter1));
  and2  gate1361(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate1362(.a(s_116), .O(gate510inter3));
  inv1  gate1363(.a(s_117), .O(gate510inter4));
  nand2 gate1364(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate1365(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate1366(.a(G1282), .O(gate510inter7));
  inv1  gate1367(.a(G1283), .O(gate510inter8));
  nand2 gate1368(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate1369(.a(s_117), .b(gate510inter3), .O(gate510inter10));
  nor2  gate1370(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate1371(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate1372(.a(gate510inter12), .b(gate510inter1), .O(G1319));

  xor2  gate1037(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate1038(.a(gate511inter0), .b(s_70), .O(gate511inter1));
  and2  gate1039(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate1040(.a(s_70), .O(gate511inter3));
  inv1  gate1041(.a(s_71), .O(gate511inter4));
  nand2 gate1042(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate1043(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate1044(.a(G1284), .O(gate511inter7));
  inv1  gate1045(.a(G1285), .O(gate511inter8));
  nand2 gate1046(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate1047(.a(s_71), .b(gate511inter3), .O(gate511inter10));
  nor2  gate1048(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate1049(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate1050(.a(gate511inter12), .b(gate511inter1), .O(G1320));

  xor2  gate701(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate702(.a(gate512inter0), .b(s_22), .O(gate512inter1));
  and2  gate703(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate704(.a(s_22), .O(gate512inter3));
  inv1  gate705(.a(s_23), .O(gate512inter4));
  nand2 gate706(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate707(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate708(.a(G1286), .O(gate512inter7));
  inv1  gate709(.a(G1287), .O(gate512inter8));
  nand2 gate710(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate711(.a(s_23), .b(gate512inter3), .O(gate512inter10));
  nor2  gate712(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate713(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate714(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule