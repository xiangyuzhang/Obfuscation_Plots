module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate715(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate716(.a(gate11inter0), .b(s_24), .O(gate11inter1));
  and2  gate717(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate718(.a(s_24), .O(gate11inter3));
  inv1  gate719(.a(s_25), .O(gate11inter4));
  nand2 gate720(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate721(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate722(.a(G5), .O(gate11inter7));
  inv1  gate723(.a(G6), .O(gate11inter8));
  nand2 gate724(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate725(.a(s_25), .b(gate11inter3), .O(gate11inter10));
  nor2  gate726(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate727(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate728(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );

  xor2  gate701(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate702(.a(gate30inter0), .b(s_22), .O(gate30inter1));
  and2  gate703(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate704(.a(s_22), .O(gate30inter3));
  inv1  gate705(.a(s_23), .O(gate30inter4));
  nand2 gate706(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate707(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate708(.a(G11), .O(gate30inter7));
  inv1  gate709(.a(G15), .O(gate30inter8));
  nand2 gate710(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate711(.a(s_23), .b(gate30inter3), .O(gate30inter10));
  nor2  gate712(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate713(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate714(.a(gate30inter12), .b(gate30inter1), .O(G329));
nand2 gate31( .a(G4), .b(G8), .O(G332) );

  xor2  gate771(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate772(.a(gate32inter0), .b(s_32), .O(gate32inter1));
  and2  gate773(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate774(.a(s_32), .O(gate32inter3));
  inv1  gate775(.a(s_33), .O(gate32inter4));
  nand2 gate776(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate777(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate778(.a(G12), .O(gate32inter7));
  inv1  gate779(.a(G16), .O(gate32inter8));
  nand2 gate780(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate781(.a(s_33), .b(gate32inter3), .O(gate32inter10));
  nor2  gate782(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate783(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate784(.a(gate32inter12), .b(gate32inter1), .O(G335));
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );

  xor2  gate645(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate646(.a(gate35inter0), .b(s_14), .O(gate35inter1));
  and2  gate647(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate648(.a(s_14), .O(gate35inter3));
  inv1  gate649(.a(s_15), .O(gate35inter4));
  nand2 gate650(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate651(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate652(.a(G18), .O(gate35inter7));
  inv1  gate653(.a(G22), .O(gate35inter8));
  nand2 gate654(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate655(.a(s_15), .b(gate35inter3), .O(gate35inter10));
  nor2  gate656(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate657(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate658(.a(gate35inter12), .b(gate35inter1), .O(G344));
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate883(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate884(.a(gate38inter0), .b(s_48), .O(gate38inter1));
  and2  gate885(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate886(.a(s_48), .O(gate38inter3));
  inv1  gate887(.a(s_49), .O(gate38inter4));
  nand2 gate888(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate889(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate890(.a(G27), .O(gate38inter7));
  inv1  gate891(.a(G31), .O(gate38inter8));
  nand2 gate892(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate893(.a(s_49), .b(gate38inter3), .O(gate38inter10));
  nor2  gate894(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate895(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate896(.a(gate38inter12), .b(gate38inter1), .O(G353));
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );

  xor2  gate1247(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate1248(.a(gate42inter0), .b(s_100), .O(gate42inter1));
  and2  gate1249(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate1250(.a(s_100), .O(gate42inter3));
  inv1  gate1251(.a(s_101), .O(gate42inter4));
  nand2 gate1252(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate1253(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate1254(.a(G2), .O(gate42inter7));
  inv1  gate1255(.a(G266), .O(gate42inter8));
  nand2 gate1256(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate1257(.a(s_101), .b(gate42inter3), .O(gate42inter10));
  nor2  gate1258(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate1259(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate1260(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );

  xor2  gate981(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate982(.a(gate44inter0), .b(s_62), .O(gate44inter1));
  and2  gate983(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate984(.a(s_62), .O(gate44inter3));
  inv1  gate985(.a(s_63), .O(gate44inter4));
  nand2 gate986(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate987(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate988(.a(G4), .O(gate44inter7));
  inv1  gate989(.a(G269), .O(gate44inter8));
  nand2 gate990(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate991(.a(s_63), .b(gate44inter3), .O(gate44inter10));
  nor2  gate992(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate993(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate994(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );

  xor2  gate1079(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate1080(.a(gate56inter0), .b(s_76), .O(gate56inter1));
  and2  gate1081(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate1082(.a(s_76), .O(gate56inter3));
  inv1  gate1083(.a(s_77), .O(gate56inter4));
  nand2 gate1084(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate1085(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate1086(.a(G16), .O(gate56inter7));
  inv1  gate1087(.a(G287), .O(gate56inter8));
  nand2 gate1088(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate1089(.a(s_77), .b(gate56inter3), .O(gate56inter10));
  nor2  gate1090(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate1091(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate1092(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate1093(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate1094(.a(gate63inter0), .b(s_78), .O(gate63inter1));
  and2  gate1095(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate1096(.a(s_78), .O(gate63inter3));
  inv1  gate1097(.a(s_79), .O(gate63inter4));
  nand2 gate1098(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate1099(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate1100(.a(G23), .O(gate63inter7));
  inv1  gate1101(.a(G299), .O(gate63inter8));
  nand2 gate1102(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate1103(.a(s_79), .b(gate63inter3), .O(gate63inter10));
  nor2  gate1104(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate1105(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate1106(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate841(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate842(.a(gate66inter0), .b(s_42), .O(gate66inter1));
  and2  gate843(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate844(.a(s_42), .O(gate66inter3));
  inv1  gate845(.a(s_43), .O(gate66inter4));
  nand2 gate846(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate847(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate848(.a(G26), .O(gate66inter7));
  inv1  gate849(.a(G302), .O(gate66inter8));
  nand2 gate850(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate851(.a(s_43), .b(gate66inter3), .O(gate66inter10));
  nor2  gate852(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate853(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate854(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate1177(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate1178(.a(gate77inter0), .b(s_90), .O(gate77inter1));
  and2  gate1179(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate1180(.a(s_90), .O(gate77inter3));
  inv1  gate1181(.a(s_91), .O(gate77inter4));
  nand2 gate1182(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate1183(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate1184(.a(G2), .O(gate77inter7));
  inv1  gate1185(.a(G320), .O(gate77inter8));
  nand2 gate1186(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate1187(.a(s_91), .b(gate77inter3), .O(gate77inter10));
  nor2  gate1188(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate1189(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate1190(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );

  xor2  gate687(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate688(.a(gate105inter0), .b(s_20), .O(gate105inter1));
  and2  gate689(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate690(.a(s_20), .O(gate105inter3));
  inv1  gate691(.a(s_21), .O(gate105inter4));
  nand2 gate692(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate693(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate694(.a(G362), .O(gate105inter7));
  inv1  gate695(.a(G363), .O(gate105inter8));
  nand2 gate696(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate697(.a(s_21), .b(gate105inter3), .O(gate105inter10));
  nor2  gate698(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate699(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate700(.a(gate105inter12), .b(gate105inter1), .O(G426));
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate897(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate898(.a(gate108inter0), .b(s_50), .O(gate108inter1));
  and2  gate899(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate900(.a(s_50), .O(gate108inter3));
  inv1  gate901(.a(s_51), .O(gate108inter4));
  nand2 gate902(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate903(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate904(.a(G368), .O(gate108inter7));
  inv1  gate905(.a(G369), .O(gate108inter8));
  nand2 gate906(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate907(.a(s_51), .b(gate108inter3), .O(gate108inter10));
  nor2  gate908(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate909(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate910(.a(gate108inter12), .b(gate108inter1), .O(G435));

  xor2  gate1107(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate1108(.a(gate109inter0), .b(s_80), .O(gate109inter1));
  and2  gate1109(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate1110(.a(s_80), .O(gate109inter3));
  inv1  gate1111(.a(s_81), .O(gate109inter4));
  nand2 gate1112(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate1113(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate1114(.a(G370), .O(gate109inter7));
  inv1  gate1115(.a(G371), .O(gate109inter8));
  nand2 gate1116(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate1117(.a(s_81), .b(gate109inter3), .O(gate109inter10));
  nor2  gate1118(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate1119(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate1120(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );

  xor2  gate785(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate786(.a(gate122inter0), .b(s_34), .O(gate122inter1));
  and2  gate787(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate788(.a(s_34), .O(gate122inter3));
  inv1  gate789(.a(s_35), .O(gate122inter4));
  nand2 gate790(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate791(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate792(.a(G396), .O(gate122inter7));
  inv1  gate793(.a(G397), .O(gate122inter8));
  nand2 gate794(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate795(.a(s_35), .b(gate122inter3), .O(gate122inter10));
  nor2  gate796(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate797(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate798(.a(gate122inter12), .b(gate122inter1), .O(G477));
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );

  xor2  gate1163(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate1164(.a(gate133inter0), .b(s_88), .O(gate133inter1));
  and2  gate1165(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate1166(.a(s_88), .O(gate133inter3));
  inv1  gate1167(.a(s_89), .O(gate133inter4));
  nand2 gate1168(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate1169(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate1170(.a(G418), .O(gate133inter7));
  inv1  gate1171(.a(G419), .O(gate133inter8));
  nand2 gate1172(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate1173(.a(s_89), .b(gate133inter3), .O(gate133inter10));
  nor2  gate1174(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate1175(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate1176(.a(gate133inter12), .b(gate133inter1), .O(G510));
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate659(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate660(.a(gate144inter0), .b(s_16), .O(gate144inter1));
  and2  gate661(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate662(.a(s_16), .O(gate144inter3));
  inv1  gate663(.a(s_17), .O(gate144inter4));
  nand2 gate664(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate665(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate666(.a(G468), .O(gate144inter7));
  inv1  gate667(.a(G471), .O(gate144inter8));
  nand2 gate668(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate669(.a(s_17), .b(gate144inter3), .O(gate144inter10));
  nor2  gate670(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate671(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate672(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate967(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate968(.a(gate150inter0), .b(s_60), .O(gate150inter1));
  and2  gate969(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate970(.a(s_60), .O(gate150inter3));
  inv1  gate971(.a(s_61), .O(gate150inter4));
  nand2 gate972(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate973(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate974(.a(G504), .O(gate150inter7));
  inv1  gate975(.a(G507), .O(gate150inter8));
  nand2 gate976(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate977(.a(s_61), .b(gate150inter3), .O(gate150inter10));
  nor2  gate978(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate979(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate980(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate589(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate590(.a(gate160inter0), .b(s_6), .O(gate160inter1));
  and2  gate591(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate592(.a(s_6), .O(gate160inter3));
  inv1  gate593(.a(s_7), .O(gate160inter4));
  nand2 gate594(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate595(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate596(.a(G447), .O(gate160inter7));
  inv1  gate597(.a(G531), .O(gate160inter8));
  nand2 gate598(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate599(.a(s_7), .b(gate160inter3), .O(gate160inter10));
  nor2  gate600(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate601(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate602(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );

  xor2  gate1205(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate1206(.a(gate171inter0), .b(s_94), .O(gate171inter1));
  and2  gate1207(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate1208(.a(s_94), .O(gate171inter3));
  inv1  gate1209(.a(s_95), .O(gate171inter4));
  nand2 gate1210(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate1211(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate1212(.a(G480), .O(gate171inter7));
  inv1  gate1213(.a(G549), .O(gate171inter8));
  nand2 gate1214(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate1215(.a(s_95), .b(gate171inter3), .O(gate171inter10));
  nor2  gate1216(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate1217(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate1218(.a(gate171inter12), .b(gate171inter1), .O(G588));
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );

  xor2  gate631(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate632(.a(gate179inter0), .b(s_12), .O(gate179inter1));
  and2  gate633(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate634(.a(s_12), .O(gate179inter3));
  inv1  gate635(.a(s_13), .O(gate179inter4));
  nand2 gate636(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate637(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate638(.a(G504), .O(gate179inter7));
  inv1  gate639(.a(G561), .O(gate179inter8));
  nand2 gate640(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate641(.a(s_13), .b(gate179inter3), .O(gate179inter10));
  nor2  gate642(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate643(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate644(.a(gate179inter12), .b(gate179inter1), .O(G596));
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate869(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate870(.a(gate197inter0), .b(s_46), .O(gate197inter1));
  and2  gate871(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate872(.a(s_46), .O(gate197inter3));
  inv1  gate873(.a(s_47), .O(gate197inter4));
  nand2 gate874(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate875(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate876(.a(G594), .O(gate197inter7));
  inv1  gate877(.a(G595), .O(gate197inter8));
  nand2 gate878(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate879(.a(s_47), .b(gate197inter3), .O(gate197inter10));
  nor2  gate880(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate881(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate882(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate757(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate758(.a(gate201inter0), .b(s_30), .O(gate201inter1));
  and2  gate759(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate760(.a(s_30), .O(gate201inter3));
  inv1  gate761(.a(s_31), .O(gate201inter4));
  nand2 gate762(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate763(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate764(.a(G602), .O(gate201inter7));
  inv1  gate765(.a(G607), .O(gate201inter8));
  nand2 gate766(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate767(.a(s_31), .b(gate201inter3), .O(gate201inter10));
  nor2  gate768(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate769(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate770(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate575(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate576(.a(gate205inter0), .b(s_4), .O(gate205inter1));
  and2  gate577(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate578(.a(s_4), .O(gate205inter3));
  inv1  gate579(.a(s_5), .O(gate205inter4));
  nand2 gate580(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate581(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate582(.a(G622), .O(gate205inter7));
  inv1  gate583(.a(G627), .O(gate205inter8));
  nand2 gate584(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate585(.a(s_5), .b(gate205inter3), .O(gate205inter10));
  nor2  gate586(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate587(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate588(.a(gate205inter12), .b(gate205inter1), .O(G678));

  xor2  gate1065(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate1066(.a(gate206inter0), .b(s_74), .O(gate206inter1));
  and2  gate1067(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate1068(.a(s_74), .O(gate206inter3));
  inv1  gate1069(.a(s_75), .O(gate206inter4));
  nand2 gate1070(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate1071(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate1072(.a(G632), .O(gate206inter7));
  inv1  gate1073(.a(G637), .O(gate206inter8));
  nand2 gate1074(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate1075(.a(s_75), .b(gate206inter3), .O(gate206inter10));
  nor2  gate1076(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate1077(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate1078(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate799(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate800(.a(gate216inter0), .b(s_36), .O(gate216inter1));
  and2  gate801(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate802(.a(s_36), .O(gate216inter3));
  inv1  gate803(.a(s_37), .O(gate216inter4));
  nand2 gate804(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate805(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate806(.a(G617), .O(gate216inter7));
  inv1  gate807(.a(G675), .O(gate216inter8));
  nand2 gate808(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate809(.a(s_37), .b(gate216inter3), .O(gate216inter10));
  nor2  gate810(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate811(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate812(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate911(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate912(.a(gate219inter0), .b(s_52), .O(gate219inter1));
  and2  gate913(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate914(.a(s_52), .O(gate219inter3));
  inv1  gate915(.a(s_53), .O(gate219inter4));
  nand2 gate916(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate917(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate918(.a(G632), .O(gate219inter7));
  inv1  gate919(.a(G681), .O(gate219inter8));
  nand2 gate920(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate921(.a(s_53), .b(gate219inter3), .O(gate219inter10));
  nor2  gate922(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate923(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate924(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate1219(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate1220(.a(gate226inter0), .b(s_96), .O(gate226inter1));
  and2  gate1221(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate1222(.a(s_96), .O(gate226inter3));
  inv1  gate1223(.a(s_97), .O(gate226inter4));
  nand2 gate1224(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate1225(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate1226(.a(G692), .O(gate226inter7));
  inv1  gate1227(.a(G693), .O(gate226inter8));
  nand2 gate1228(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate1229(.a(s_97), .b(gate226inter3), .O(gate226inter10));
  nor2  gate1230(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate1231(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate1232(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate827(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate828(.a(gate231inter0), .b(s_40), .O(gate231inter1));
  and2  gate829(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate830(.a(s_40), .O(gate231inter3));
  inv1  gate831(.a(s_41), .O(gate231inter4));
  nand2 gate832(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate833(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate834(.a(G702), .O(gate231inter7));
  inv1  gate835(.a(G703), .O(gate231inter8));
  nand2 gate836(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate837(.a(s_41), .b(gate231inter3), .O(gate231inter10));
  nor2  gate838(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate839(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate840(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );

  xor2  gate1051(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate1052(.a(gate234inter0), .b(s_72), .O(gate234inter1));
  and2  gate1053(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate1054(.a(s_72), .O(gate234inter3));
  inv1  gate1055(.a(s_73), .O(gate234inter4));
  nand2 gate1056(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1057(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1058(.a(G245), .O(gate234inter7));
  inv1  gate1059(.a(G721), .O(gate234inter8));
  nand2 gate1060(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1061(.a(s_73), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1062(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1063(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1064(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate953(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate954(.a(gate243inter0), .b(s_58), .O(gate243inter1));
  and2  gate955(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate956(.a(s_58), .O(gate243inter3));
  inv1  gate957(.a(s_59), .O(gate243inter4));
  nand2 gate958(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate959(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate960(.a(G245), .O(gate243inter7));
  inv1  gate961(.a(G733), .O(gate243inter8));
  nand2 gate962(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate963(.a(s_59), .b(gate243inter3), .O(gate243inter10));
  nor2  gate964(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate965(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate966(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate1191(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate1192(.a(gate249inter0), .b(s_92), .O(gate249inter1));
  and2  gate1193(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate1194(.a(s_92), .O(gate249inter3));
  inv1  gate1195(.a(s_93), .O(gate249inter4));
  nand2 gate1196(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate1197(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate1198(.a(G254), .O(gate249inter7));
  inv1  gate1199(.a(G742), .O(gate249inter8));
  nand2 gate1200(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate1201(.a(s_93), .b(gate249inter3), .O(gate249inter10));
  nor2  gate1202(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate1203(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate1204(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );

  xor2  gate729(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate730(.a(gate273inter0), .b(s_26), .O(gate273inter1));
  and2  gate731(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate732(.a(s_26), .O(gate273inter3));
  inv1  gate733(.a(s_27), .O(gate273inter4));
  nand2 gate734(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate735(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate736(.a(G642), .O(gate273inter7));
  inv1  gate737(.a(G794), .O(gate273inter8));
  nand2 gate738(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate739(.a(s_27), .b(gate273inter3), .O(gate273inter10));
  nor2  gate740(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate741(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate742(.a(gate273inter12), .b(gate273inter1), .O(G818));
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate855(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate856(.a(gate278inter0), .b(s_44), .O(gate278inter1));
  and2  gate857(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate858(.a(s_44), .O(gate278inter3));
  inv1  gate859(.a(s_45), .O(gate278inter4));
  nand2 gate860(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate861(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate862(.a(G776), .O(gate278inter7));
  inv1  gate863(.a(G800), .O(gate278inter8));
  nand2 gate864(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate865(.a(s_45), .b(gate278inter3), .O(gate278inter10));
  nor2  gate866(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate867(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate868(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate925(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate926(.a(gate287inter0), .b(s_54), .O(gate287inter1));
  and2  gate927(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate928(.a(s_54), .O(gate287inter3));
  inv1  gate929(.a(s_55), .O(gate287inter4));
  nand2 gate930(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate931(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate932(.a(G663), .O(gate287inter7));
  inv1  gate933(.a(G815), .O(gate287inter8));
  nand2 gate934(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate935(.a(s_55), .b(gate287inter3), .O(gate287inter10));
  nor2  gate936(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate937(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate938(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate1037(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate1038(.a(gate390inter0), .b(s_70), .O(gate390inter1));
  and2  gate1039(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate1040(.a(s_70), .O(gate390inter3));
  inv1  gate1041(.a(s_71), .O(gate390inter4));
  nand2 gate1042(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate1043(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate1044(.a(G4), .O(gate390inter7));
  inv1  gate1045(.a(G1045), .O(gate390inter8));
  nand2 gate1046(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate1047(.a(s_71), .b(gate390inter3), .O(gate390inter10));
  nor2  gate1048(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate1049(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate1050(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );

  xor2  gate547(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate548(.a(gate418inter0), .b(s_0), .O(gate418inter1));
  and2  gate549(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate550(.a(s_0), .O(gate418inter3));
  inv1  gate551(.a(s_1), .O(gate418inter4));
  nand2 gate552(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate553(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate554(.a(G32), .O(gate418inter7));
  inv1  gate555(.a(G1129), .O(gate418inter8));
  nand2 gate556(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate557(.a(s_1), .b(gate418inter3), .O(gate418inter10));
  nor2  gate558(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate559(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate560(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate813(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate814(.a(gate422inter0), .b(s_38), .O(gate422inter1));
  and2  gate815(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate816(.a(s_38), .O(gate422inter3));
  inv1  gate817(.a(s_39), .O(gate422inter4));
  nand2 gate818(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate819(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate820(.a(G1039), .O(gate422inter7));
  inv1  gate821(.a(G1135), .O(gate422inter8));
  nand2 gate822(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate823(.a(s_39), .b(gate422inter3), .O(gate422inter10));
  nor2  gate824(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate825(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate826(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate617(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate618(.a(gate425inter0), .b(s_10), .O(gate425inter1));
  and2  gate619(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate620(.a(s_10), .O(gate425inter3));
  inv1  gate621(.a(s_11), .O(gate425inter4));
  nand2 gate622(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate623(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate624(.a(G4), .O(gate425inter7));
  inv1  gate625(.a(G1141), .O(gate425inter8));
  nand2 gate626(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate627(.a(s_11), .b(gate425inter3), .O(gate425inter10));
  nor2  gate628(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate629(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate630(.a(gate425inter12), .b(gate425inter1), .O(G1234));

  xor2  gate1149(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate1150(.a(gate426inter0), .b(s_86), .O(gate426inter1));
  and2  gate1151(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate1152(.a(s_86), .O(gate426inter3));
  inv1  gate1153(.a(s_87), .O(gate426inter4));
  nand2 gate1154(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate1155(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate1156(.a(G1045), .O(gate426inter7));
  inv1  gate1157(.a(G1141), .O(gate426inter8));
  nand2 gate1158(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate1159(.a(s_87), .b(gate426inter3), .O(gate426inter10));
  nor2  gate1160(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate1161(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate1162(.a(gate426inter12), .b(gate426inter1), .O(G1235));

  xor2  gate1023(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate1024(.a(gate427inter0), .b(s_68), .O(gate427inter1));
  and2  gate1025(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate1026(.a(s_68), .O(gate427inter3));
  inv1  gate1027(.a(s_69), .O(gate427inter4));
  nand2 gate1028(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate1029(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate1030(.a(G5), .O(gate427inter7));
  inv1  gate1031(.a(G1144), .O(gate427inter8));
  nand2 gate1032(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate1033(.a(s_69), .b(gate427inter3), .O(gate427inter10));
  nor2  gate1034(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate1035(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate1036(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate1009(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate1010(.a(gate430inter0), .b(s_66), .O(gate430inter1));
  and2  gate1011(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate1012(.a(s_66), .O(gate430inter3));
  inv1  gate1013(.a(s_67), .O(gate430inter4));
  nand2 gate1014(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate1015(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate1016(.a(G1051), .O(gate430inter7));
  inv1  gate1017(.a(G1147), .O(gate430inter8));
  nand2 gate1018(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate1019(.a(s_67), .b(gate430inter3), .O(gate430inter10));
  nor2  gate1020(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate1021(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate1022(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );

  xor2  gate743(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate744(.a(gate449inter0), .b(s_28), .O(gate449inter1));
  and2  gate745(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate746(.a(s_28), .O(gate449inter3));
  inv1  gate747(.a(s_29), .O(gate449inter4));
  nand2 gate748(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate749(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate750(.a(G16), .O(gate449inter7));
  inv1  gate751(.a(G1177), .O(gate449inter8));
  nand2 gate752(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate753(.a(s_29), .b(gate449inter3), .O(gate449inter10));
  nor2  gate754(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate755(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate756(.a(gate449inter12), .b(gate449inter1), .O(G1258));

  xor2  gate995(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate996(.a(gate450inter0), .b(s_64), .O(gate450inter1));
  and2  gate997(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate998(.a(s_64), .O(gate450inter3));
  inv1  gate999(.a(s_65), .O(gate450inter4));
  nand2 gate1000(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate1001(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate1002(.a(G1081), .O(gate450inter7));
  inv1  gate1003(.a(G1177), .O(gate450inter8));
  nand2 gate1004(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate1005(.a(s_65), .b(gate450inter3), .O(gate450inter10));
  nor2  gate1006(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate1007(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate1008(.a(gate450inter12), .b(gate450inter1), .O(G1259));
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate1233(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate1234(.a(gate464inter0), .b(s_98), .O(gate464inter1));
  and2  gate1235(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate1236(.a(s_98), .O(gate464inter3));
  inv1  gate1237(.a(s_99), .O(gate464inter4));
  nand2 gate1238(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate1239(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate1240(.a(G1102), .O(gate464inter7));
  inv1  gate1241(.a(G1198), .O(gate464inter8));
  nand2 gate1242(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate1243(.a(s_99), .b(gate464inter3), .O(gate464inter10));
  nor2  gate1244(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate1245(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate1246(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );

  xor2  gate1135(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate1136(.a(gate479inter0), .b(s_84), .O(gate479inter1));
  and2  gate1137(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate1138(.a(s_84), .O(gate479inter3));
  inv1  gate1139(.a(s_85), .O(gate479inter4));
  nand2 gate1140(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate1141(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate1142(.a(G31), .O(gate479inter7));
  inv1  gate1143(.a(G1222), .O(gate479inter8));
  nand2 gate1144(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate1145(.a(s_85), .b(gate479inter3), .O(gate479inter10));
  nor2  gate1146(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate1147(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate1148(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate939(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate940(.a(gate481inter0), .b(s_56), .O(gate481inter1));
  and2  gate941(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate942(.a(s_56), .O(gate481inter3));
  inv1  gate943(.a(s_57), .O(gate481inter4));
  nand2 gate944(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate945(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate946(.a(G32), .O(gate481inter7));
  inv1  gate947(.a(G1225), .O(gate481inter8));
  nand2 gate948(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate949(.a(s_57), .b(gate481inter3), .O(gate481inter10));
  nor2  gate950(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate951(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate952(.a(gate481inter12), .b(gate481inter1), .O(G1290));

  xor2  gate603(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate604(.a(gate482inter0), .b(s_8), .O(gate482inter1));
  and2  gate605(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate606(.a(s_8), .O(gate482inter3));
  inv1  gate607(.a(s_9), .O(gate482inter4));
  nand2 gate608(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate609(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate610(.a(G1129), .O(gate482inter7));
  inv1  gate611(.a(G1225), .O(gate482inter8));
  nand2 gate612(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate613(.a(s_9), .b(gate482inter3), .O(gate482inter10));
  nor2  gate614(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate615(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate616(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate1121(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate1122(.a(gate487inter0), .b(s_82), .O(gate487inter1));
  and2  gate1123(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate1124(.a(s_82), .O(gate487inter3));
  inv1  gate1125(.a(s_83), .O(gate487inter4));
  nand2 gate1126(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate1127(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate1128(.a(G1236), .O(gate487inter7));
  inv1  gate1129(.a(G1237), .O(gate487inter8));
  nand2 gate1130(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate1131(.a(s_83), .b(gate487inter3), .O(gate487inter10));
  nor2  gate1132(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate1133(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate1134(.a(gate487inter12), .b(gate487inter1), .O(G1296));
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );

  xor2  gate673(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate674(.a(gate495inter0), .b(s_18), .O(gate495inter1));
  and2  gate675(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate676(.a(s_18), .O(gate495inter3));
  inv1  gate677(.a(s_19), .O(gate495inter4));
  nand2 gate678(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate679(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate680(.a(G1252), .O(gate495inter7));
  inv1  gate681(.a(G1253), .O(gate495inter8));
  nand2 gate682(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate683(.a(s_19), .b(gate495inter3), .O(gate495inter10));
  nor2  gate684(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate685(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate686(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate561(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate562(.a(gate508inter0), .b(s_2), .O(gate508inter1));
  and2  gate563(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate564(.a(s_2), .O(gate508inter3));
  inv1  gate565(.a(s_3), .O(gate508inter4));
  nand2 gate566(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate567(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate568(.a(G1278), .O(gate508inter7));
  inv1  gate569(.a(G1279), .O(gate508inter8));
  nand2 gate570(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate571(.a(s_3), .b(gate508inter3), .O(gate508inter10));
  nor2  gate572(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate573(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate574(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule