module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate1891(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate1892(.a(gate12inter0), .b(s_192), .O(gate12inter1));
  and2  gate1893(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate1894(.a(s_192), .O(gate12inter3));
  inv1  gate1895(.a(s_193), .O(gate12inter4));
  nand2 gate1896(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate1897(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate1898(.a(G7), .O(gate12inter7));
  inv1  gate1899(.a(G8), .O(gate12inter8));
  nand2 gate1900(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate1901(.a(s_193), .b(gate12inter3), .O(gate12inter10));
  nor2  gate1902(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate1903(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate1904(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );

  xor2  gate1401(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate1402(.a(gate14inter0), .b(s_122), .O(gate14inter1));
  and2  gate1403(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate1404(.a(s_122), .O(gate14inter3));
  inv1  gate1405(.a(s_123), .O(gate14inter4));
  nand2 gate1406(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate1407(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate1408(.a(G11), .O(gate14inter7));
  inv1  gate1409(.a(G12), .O(gate14inter8));
  nand2 gate1410(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate1411(.a(s_123), .b(gate14inter3), .O(gate14inter10));
  nor2  gate1412(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate1413(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate1414(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate701(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate702(.a(gate16inter0), .b(s_22), .O(gate16inter1));
  and2  gate703(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate704(.a(s_22), .O(gate16inter3));
  inv1  gate705(.a(s_23), .O(gate16inter4));
  nand2 gate706(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate707(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate708(.a(G15), .O(gate16inter7));
  inv1  gate709(.a(G16), .O(gate16inter8));
  nand2 gate710(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate711(.a(s_23), .b(gate16inter3), .O(gate16inter10));
  nor2  gate712(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate713(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate714(.a(gate16inter12), .b(gate16inter1), .O(G287));

  xor2  gate1835(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate1836(.a(gate17inter0), .b(s_184), .O(gate17inter1));
  and2  gate1837(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate1838(.a(s_184), .O(gate17inter3));
  inv1  gate1839(.a(s_185), .O(gate17inter4));
  nand2 gate1840(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate1841(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate1842(.a(G17), .O(gate17inter7));
  inv1  gate1843(.a(G18), .O(gate17inter8));
  nand2 gate1844(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate1845(.a(s_185), .b(gate17inter3), .O(gate17inter10));
  nor2  gate1846(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate1847(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate1848(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate1331(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate1332(.a(gate26inter0), .b(s_112), .O(gate26inter1));
  and2  gate1333(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate1334(.a(s_112), .O(gate26inter3));
  inv1  gate1335(.a(s_113), .O(gate26inter4));
  nand2 gate1336(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate1337(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate1338(.a(G9), .O(gate26inter7));
  inv1  gate1339(.a(G13), .O(gate26inter8));
  nand2 gate1340(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate1341(.a(s_113), .b(gate26inter3), .O(gate26inter10));
  nor2  gate1342(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate1343(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate1344(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate1989(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate1990(.a(gate28inter0), .b(s_206), .O(gate28inter1));
  and2  gate1991(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate1992(.a(s_206), .O(gate28inter3));
  inv1  gate1993(.a(s_207), .O(gate28inter4));
  nand2 gate1994(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate1995(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate1996(.a(G10), .O(gate28inter7));
  inv1  gate1997(.a(G14), .O(gate28inter8));
  nand2 gate1998(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate1999(.a(s_207), .b(gate28inter3), .O(gate28inter10));
  nor2  gate2000(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate2001(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate2002(.a(gate28inter12), .b(gate28inter1), .O(G323));
nand2 gate29( .a(G3), .b(G7), .O(G326) );

  xor2  gate1247(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate1248(.a(gate30inter0), .b(s_100), .O(gate30inter1));
  and2  gate1249(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate1250(.a(s_100), .O(gate30inter3));
  inv1  gate1251(.a(s_101), .O(gate30inter4));
  nand2 gate1252(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate1253(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate1254(.a(G11), .O(gate30inter7));
  inv1  gate1255(.a(G15), .O(gate30inter8));
  nand2 gate1256(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate1257(.a(s_101), .b(gate30inter3), .O(gate30inter10));
  nor2  gate1258(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate1259(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate1260(.a(gate30inter12), .b(gate30inter1), .O(G329));
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate1919(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate1920(.a(gate33inter0), .b(s_196), .O(gate33inter1));
  and2  gate1921(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate1922(.a(s_196), .O(gate33inter3));
  inv1  gate1923(.a(s_197), .O(gate33inter4));
  nand2 gate1924(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate1925(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate1926(.a(G17), .O(gate33inter7));
  inv1  gate1927(.a(G21), .O(gate33inter8));
  nand2 gate1928(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate1929(.a(s_197), .b(gate33inter3), .O(gate33inter10));
  nor2  gate1930(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate1931(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate1932(.a(gate33inter12), .b(gate33inter1), .O(G338));
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate1723(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate1724(.a(gate37inter0), .b(s_168), .O(gate37inter1));
  and2  gate1725(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate1726(.a(s_168), .O(gate37inter3));
  inv1  gate1727(.a(s_169), .O(gate37inter4));
  nand2 gate1728(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate1729(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate1730(.a(G19), .O(gate37inter7));
  inv1  gate1731(.a(G23), .O(gate37inter8));
  nand2 gate1732(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate1733(.a(s_169), .b(gate37inter3), .O(gate37inter10));
  nor2  gate1734(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate1735(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate1736(.a(gate37inter12), .b(gate37inter1), .O(G350));

  xor2  gate799(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate800(.a(gate38inter0), .b(s_36), .O(gate38inter1));
  and2  gate801(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate802(.a(s_36), .O(gate38inter3));
  inv1  gate803(.a(s_37), .O(gate38inter4));
  nand2 gate804(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate805(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate806(.a(G27), .O(gate38inter7));
  inv1  gate807(.a(G31), .O(gate38inter8));
  nand2 gate808(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate809(.a(s_37), .b(gate38inter3), .O(gate38inter10));
  nor2  gate810(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate811(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate812(.a(gate38inter12), .b(gate38inter1), .O(G353));
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate575(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate576(.a(gate51inter0), .b(s_4), .O(gate51inter1));
  and2  gate577(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate578(.a(s_4), .O(gate51inter3));
  inv1  gate579(.a(s_5), .O(gate51inter4));
  nand2 gate580(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate581(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate582(.a(G11), .O(gate51inter7));
  inv1  gate583(.a(G281), .O(gate51inter8));
  nand2 gate584(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate585(.a(s_5), .b(gate51inter3), .O(gate51inter10));
  nor2  gate586(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate587(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate588(.a(gate51inter12), .b(gate51inter1), .O(G372));
nand2 gate52( .a(G12), .b(G281), .O(G373) );

  xor2  gate911(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate912(.a(gate53inter0), .b(s_52), .O(gate53inter1));
  and2  gate913(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate914(.a(s_52), .O(gate53inter3));
  inv1  gate915(.a(s_53), .O(gate53inter4));
  nand2 gate916(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate917(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate918(.a(G13), .O(gate53inter7));
  inv1  gate919(.a(G284), .O(gate53inter8));
  nand2 gate920(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate921(.a(s_53), .b(gate53inter3), .O(gate53inter10));
  nor2  gate922(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate923(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate924(.a(gate53inter12), .b(gate53inter1), .O(G374));
nand2 gate54( .a(G14), .b(G284), .O(G375) );

  xor2  gate1009(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate1010(.a(gate55inter0), .b(s_66), .O(gate55inter1));
  and2  gate1011(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate1012(.a(s_66), .O(gate55inter3));
  inv1  gate1013(.a(s_67), .O(gate55inter4));
  nand2 gate1014(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate1015(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate1016(.a(G15), .O(gate55inter7));
  inv1  gate1017(.a(G287), .O(gate55inter8));
  nand2 gate1018(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate1019(.a(s_67), .b(gate55inter3), .O(gate55inter10));
  nor2  gate1020(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate1021(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate1022(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate1877(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate1878(.a(gate60inter0), .b(s_190), .O(gate60inter1));
  and2  gate1879(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate1880(.a(s_190), .O(gate60inter3));
  inv1  gate1881(.a(s_191), .O(gate60inter4));
  nand2 gate1882(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate1883(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate1884(.a(G20), .O(gate60inter7));
  inv1  gate1885(.a(G293), .O(gate60inter8));
  nand2 gate1886(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate1887(.a(s_191), .b(gate60inter3), .O(gate60inter10));
  nor2  gate1888(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate1889(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate1890(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate1023(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate1024(.a(gate63inter0), .b(s_68), .O(gate63inter1));
  and2  gate1025(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate1026(.a(s_68), .O(gate63inter3));
  inv1  gate1027(.a(s_69), .O(gate63inter4));
  nand2 gate1028(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate1029(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate1030(.a(G23), .O(gate63inter7));
  inv1  gate1031(.a(G299), .O(gate63inter8));
  nand2 gate1032(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate1033(.a(s_69), .b(gate63inter3), .O(gate63inter10));
  nor2  gate1034(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate1035(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate1036(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate1233(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate1234(.a(gate66inter0), .b(s_98), .O(gate66inter1));
  and2  gate1235(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate1236(.a(s_98), .O(gate66inter3));
  inv1  gate1237(.a(s_99), .O(gate66inter4));
  nand2 gate1238(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate1239(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate1240(.a(G26), .O(gate66inter7));
  inv1  gate1241(.a(G302), .O(gate66inter8));
  nand2 gate1242(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate1243(.a(s_99), .b(gate66inter3), .O(gate66inter10));
  nor2  gate1244(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate1245(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate1246(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate1275(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate1276(.a(gate69inter0), .b(s_104), .O(gate69inter1));
  and2  gate1277(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate1278(.a(s_104), .O(gate69inter3));
  inv1  gate1279(.a(s_105), .O(gate69inter4));
  nand2 gate1280(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate1281(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate1282(.a(G29), .O(gate69inter7));
  inv1  gate1283(.a(G308), .O(gate69inter8));
  nand2 gate1284(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate1285(.a(s_105), .b(gate69inter3), .O(gate69inter10));
  nor2  gate1286(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate1287(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate1288(.a(gate69inter12), .b(gate69inter1), .O(G390));
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate1191(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate1192(.a(gate74inter0), .b(s_92), .O(gate74inter1));
  and2  gate1193(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate1194(.a(s_92), .O(gate74inter3));
  inv1  gate1195(.a(s_93), .O(gate74inter4));
  nand2 gate1196(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate1197(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate1198(.a(G5), .O(gate74inter7));
  inv1  gate1199(.a(G314), .O(gate74inter8));
  nand2 gate1200(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate1201(.a(s_93), .b(gate74inter3), .O(gate74inter10));
  nor2  gate1202(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate1203(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate1204(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate1289(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate1290(.a(gate86inter0), .b(s_106), .O(gate86inter1));
  and2  gate1291(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate1292(.a(s_106), .O(gate86inter3));
  inv1  gate1293(.a(s_107), .O(gate86inter4));
  nand2 gate1294(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate1295(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate1296(.a(G8), .O(gate86inter7));
  inv1  gate1297(.a(G332), .O(gate86inter8));
  nand2 gate1298(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate1299(.a(s_107), .b(gate86inter3), .O(gate86inter10));
  nor2  gate1300(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate1301(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate1302(.a(gate86inter12), .b(gate86inter1), .O(G407));

  xor2  gate1611(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate1612(.a(gate87inter0), .b(s_152), .O(gate87inter1));
  and2  gate1613(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate1614(.a(s_152), .O(gate87inter3));
  inv1  gate1615(.a(s_153), .O(gate87inter4));
  nand2 gate1616(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate1617(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate1618(.a(G12), .O(gate87inter7));
  inv1  gate1619(.a(G335), .O(gate87inter8));
  nand2 gate1620(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate1621(.a(s_153), .b(gate87inter3), .O(gate87inter10));
  nor2  gate1622(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate1623(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate1624(.a(gate87inter12), .b(gate87inter1), .O(G408));

  xor2  gate1849(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate1850(.a(gate88inter0), .b(s_186), .O(gate88inter1));
  and2  gate1851(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate1852(.a(s_186), .O(gate88inter3));
  inv1  gate1853(.a(s_187), .O(gate88inter4));
  nand2 gate1854(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate1855(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate1856(.a(G16), .O(gate88inter7));
  inv1  gate1857(.a(G335), .O(gate88inter8));
  nand2 gate1858(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate1859(.a(s_187), .b(gate88inter3), .O(gate88inter10));
  nor2  gate1860(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate1861(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate1862(.a(gate88inter12), .b(gate88inter1), .O(G409));

  xor2  gate869(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate870(.a(gate89inter0), .b(s_46), .O(gate89inter1));
  and2  gate871(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate872(.a(s_46), .O(gate89inter3));
  inv1  gate873(.a(s_47), .O(gate89inter4));
  nand2 gate874(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate875(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate876(.a(G17), .O(gate89inter7));
  inv1  gate877(.a(G338), .O(gate89inter8));
  nand2 gate878(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate879(.a(s_47), .b(gate89inter3), .O(gate89inter10));
  nor2  gate880(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate881(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate882(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate687(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate688(.a(gate91inter0), .b(s_20), .O(gate91inter1));
  and2  gate689(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate690(.a(s_20), .O(gate91inter3));
  inv1  gate691(.a(s_21), .O(gate91inter4));
  nand2 gate692(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate693(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate694(.a(G25), .O(gate91inter7));
  inv1  gate695(.a(G341), .O(gate91inter8));
  nand2 gate696(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate697(.a(s_21), .b(gate91inter3), .O(gate91inter10));
  nor2  gate698(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate699(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate700(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );

  xor2  gate1933(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate1934(.a(gate93inter0), .b(s_198), .O(gate93inter1));
  and2  gate1935(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate1936(.a(s_198), .O(gate93inter3));
  inv1  gate1937(.a(s_199), .O(gate93inter4));
  nand2 gate1938(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate1939(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate1940(.a(G18), .O(gate93inter7));
  inv1  gate1941(.a(G344), .O(gate93inter8));
  nand2 gate1942(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate1943(.a(s_199), .b(gate93inter3), .O(gate93inter10));
  nor2  gate1944(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate1945(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate1946(.a(gate93inter12), .b(gate93inter1), .O(G414));
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );

  xor2  gate617(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate618(.a(gate97inter0), .b(s_10), .O(gate97inter1));
  and2  gate619(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate620(.a(s_10), .O(gate97inter3));
  inv1  gate621(.a(s_11), .O(gate97inter4));
  nand2 gate622(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate623(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate624(.a(G19), .O(gate97inter7));
  inv1  gate625(.a(G350), .O(gate97inter8));
  nand2 gate626(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate627(.a(s_11), .b(gate97inter3), .O(gate97inter10));
  nor2  gate628(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate629(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate630(.a(gate97inter12), .b(gate97inter1), .O(G418));
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate1695(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate1696(.a(gate99inter0), .b(s_164), .O(gate99inter1));
  and2  gate1697(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate1698(.a(s_164), .O(gate99inter3));
  inv1  gate1699(.a(s_165), .O(gate99inter4));
  nand2 gate1700(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate1701(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate1702(.a(G27), .O(gate99inter7));
  inv1  gate1703(.a(G353), .O(gate99inter8));
  nand2 gate1704(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate1705(.a(s_165), .b(gate99inter3), .O(gate99inter10));
  nor2  gate1706(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate1707(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate1708(.a(gate99inter12), .b(gate99inter1), .O(G420));

  xor2  gate1527(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate1528(.a(gate100inter0), .b(s_140), .O(gate100inter1));
  and2  gate1529(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate1530(.a(s_140), .O(gate100inter3));
  inv1  gate1531(.a(s_141), .O(gate100inter4));
  nand2 gate1532(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate1533(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate1534(.a(G31), .O(gate100inter7));
  inv1  gate1535(.a(G353), .O(gate100inter8));
  nand2 gate1536(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate1537(.a(s_141), .b(gate100inter3), .O(gate100inter10));
  nor2  gate1538(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate1539(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate1540(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate995(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate996(.a(gate102inter0), .b(s_64), .O(gate102inter1));
  and2  gate997(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate998(.a(s_64), .O(gate102inter3));
  inv1  gate999(.a(s_65), .O(gate102inter4));
  nand2 gate1000(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate1001(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate1002(.a(G24), .O(gate102inter7));
  inv1  gate1003(.a(G356), .O(gate102inter8));
  nand2 gate1004(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate1005(.a(s_65), .b(gate102inter3), .O(gate102inter10));
  nor2  gate1006(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate1007(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate1008(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate1317(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate1318(.a(gate104inter0), .b(s_110), .O(gate104inter1));
  and2  gate1319(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate1320(.a(s_110), .O(gate104inter3));
  inv1  gate1321(.a(s_111), .O(gate104inter4));
  nand2 gate1322(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate1323(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate1324(.a(G32), .O(gate104inter7));
  inv1  gate1325(.a(G359), .O(gate104inter8));
  nand2 gate1326(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate1327(.a(s_111), .b(gate104inter3), .O(gate104inter10));
  nor2  gate1328(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate1329(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate1330(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate757(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate758(.a(gate107inter0), .b(s_30), .O(gate107inter1));
  and2  gate759(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate760(.a(s_30), .O(gate107inter3));
  inv1  gate761(.a(s_31), .O(gate107inter4));
  nand2 gate762(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate763(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate764(.a(G366), .O(gate107inter7));
  inv1  gate765(.a(G367), .O(gate107inter8));
  nand2 gate766(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate767(.a(s_31), .b(gate107inter3), .O(gate107inter10));
  nor2  gate768(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate769(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate770(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate1457(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate1458(.a(gate110inter0), .b(s_130), .O(gate110inter1));
  and2  gate1459(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate1460(.a(s_130), .O(gate110inter3));
  inv1  gate1461(.a(s_131), .O(gate110inter4));
  nand2 gate1462(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1463(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1464(.a(G372), .O(gate110inter7));
  inv1  gate1465(.a(G373), .O(gate110inter8));
  nand2 gate1466(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1467(.a(s_131), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1468(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1469(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1470(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate1065(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate1066(.a(gate124inter0), .b(s_74), .O(gate124inter1));
  and2  gate1067(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate1068(.a(s_74), .O(gate124inter3));
  inv1  gate1069(.a(s_75), .O(gate124inter4));
  nand2 gate1070(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate1071(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate1072(.a(G400), .O(gate124inter7));
  inv1  gate1073(.a(G401), .O(gate124inter8));
  nand2 gate1074(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate1075(.a(s_75), .b(gate124inter3), .O(gate124inter10));
  nor2  gate1076(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate1077(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate1078(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );

  xor2  gate1681(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate1682(.a(gate127inter0), .b(s_162), .O(gate127inter1));
  and2  gate1683(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate1684(.a(s_162), .O(gate127inter3));
  inv1  gate1685(.a(s_163), .O(gate127inter4));
  nand2 gate1686(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate1687(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate1688(.a(G406), .O(gate127inter7));
  inv1  gate1689(.a(G407), .O(gate127inter8));
  nand2 gate1690(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate1691(.a(s_163), .b(gate127inter3), .O(gate127inter10));
  nor2  gate1692(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate1693(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate1694(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate1583(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate1584(.a(gate132inter0), .b(s_148), .O(gate132inter1));
  and2  gate1585(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate1586(.a(s_148), .O(gate132inter3));
  inv1  gate1587(.a(s_149), .O(gate132inter4));
  nand2 gate1588(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate1589(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate1590(.a(G416), .O(gate132inter7));
  inv1  gate1591(.a(G417), .O(gate132inter8));
  nand2 gate1592(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate1593(.a(s_149), .b(gate132inter3), .O(gate132inter10));
  nor2  gate1594(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate1595(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate1596(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );

  xor2  gate1779(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate1780(.a(gate145inter0), .b(s_176), .O(gate145inter1));
  and2  gate1781(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate1782(.a(s_176), .O(gate145inter3));
  inv1  gate1783(.a(s_177), .O(gate145inter4));
  nand2 gate1784(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate1785(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate1786(.a(G474), .O(gate145inter7));
  inv1  gate1787(.a(G477), .O(gate145inter8));
  nand2 gate1788(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate1789(.a(s_177), .b(gate145inter3), .O(gate145inter10));
  nor2  gate1790(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate1791(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate1792(.a(gate145inter12), .b(gate145inter1), .O(G546));

  xor2  gate1107(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate1108(.a(gate146inter0), .b(s_80), .O(gate146inter1));
  and2  gate1109(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate1110(.a(s_80), .O(gate146inter3));
  inv1  gate1111(.a(s_81), .O(gate146inter4));
  nand2 gate1112(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate1113(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate1114(.a(G480), .O(gate146inter7));
  inv1  gate1115(.a(G483), .O(gate146inter8));
  nand2 gate1116(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate1117(.a(s_81), .b(gate146inter3), .O(gate146inter10));
  nor2  gate1118(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate1119(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate1120(.a(gate146inter12), .b(gate146inter1), .O(G549));
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate2003(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate2004(.a(gate150inter0), .b(s_208), .O(gate150inter1));
  and2  gate2005(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate2006(.a(s_208), .O(gate150inter3));
  inv1  gate2007(.a(s_209), .O(gate150inter4));
  nand2 gate2008(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate2009(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate2010(.a(G504), .O(gate150inter7));
  inv1  gate2011(.a(G507), .O(gate150inter8));
  nand2 gate2012(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate2013(.a(s_209), .b(gate150inter3), .O(gate150inter10));
  nor2  gate2014(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate2015(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate2016(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate1387(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate1388(.a(gate154inter0), .b(s_120), .O(gate154inter1));
  and2  gate1389(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate1390(.a(s_120), .O(gate154inter3));
  inv1  gate1391(.a(s_121), .O(gate154inter4));
  nand2 gate1392(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate1393(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate1394(.a(G429), .O(gate154inter7));
  inv1  gate1395(.a(G522), .O(gate154inter8));
  nand2 gate1396(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate1397(.a(s_121), .b(gate154inter3), .O(gate154inter10));
  nor2  gate1398(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate1399(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate1400(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate1261(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate1262(.a(gate160inter0), .b(s_102), .O(gate160inter1));
  and2  gate1263(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate1264(.a(s_102), .O(gate160inter3));
  inv1  gate1265(.a(s_103), .O(gate160inter4));
  nand2 gate1266(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate1267(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate1268(.a(G447), .O(gate160inter7));
  inv1  gate1269(.a(G531), .O(gate160inter8));
  nand2 gate1270(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate1271(.a(s_103), .b(gate160inter3), .O(gate160inter10));
  nor2  gate1272(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate1273(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate1274(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate1541(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate1542(.a(gate162inter0), .b(s_142), .O(gate162inter1));
  and2  gate1543(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate1544(.a(s_142), .O(gate162inter3));
  inv1  gate1545(.a(s_143), .O(gate162inter4));
  nand2 gate1546(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate1547(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate1548(.a(G453), .O(gate162inter7));
  inv1  gate1549(.a(G534), .O(gate162inter8));
  nand2 gate1550(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate1551(.a(s_143), .b(gate162inter3), .O(gate162inter10));
  nor2  gate1552(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate1553(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate1554(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate1975(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate1976(.a(gate165inter0), .b(s_204), .O(gate165inter1));
  and2  gate1977(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate1978(.a(s_204), .O(gate165inter3));
  inv1  gate1979(.a(s_205), .O(gate165inter4));
  nand2 gate1980(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate1981(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate1982(.a(G462), .O(gate165inter7));
  inv1  gate1983(.a(G540), .O(gate165inter8));
  nand2 gate1984(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate1985(.a(s_205), .b(gate165inter3), .O(gate165inter10));
  nor2  gate1986(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate1987(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate1988(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );

  xor2  gate1345(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate1346(.a(gate167inter0), .b(s_114), .O(gate167inter1));
  and2  gate1347(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate1348(.a(s_114), .O(gate167inter3));
  inv1  gate1349(.a(s_115), .O(gate167inter4));
  nand2 gate1350(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate1351(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate1352(.a(G468), .O(gate167inter7));
  inv1  gate1353(.a(G543), .O(gate167inter8));
  nand2 gate1354(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate1355(.a(s_115), .b(gate167inter3), .O(gate167inter10));
  nor2  gate1356(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate1357(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate1358(.a(gate167inter12), .b(gate167inter1), .O(G584));

  xor2  gate1513(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate1514(.a(gate168inter0), .b(s_138), .O(gate168inter1));
  and2  gate1515(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate1516(.a(s_138), .O(gate168inter3));
  inv1  gate1517(.a(s_139), .O(gate168inter4));
  nand2 gate1518(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate1519(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate1520(.a(G471), .O(gate168inter7));
  inv1  gate1521(.a(G543), .O(gate168inter8));
  nand2 gate1522(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate1523(.a(s_139), .b(gate168inter3), .O(gate168inter10));
  nor2  gate1524(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate1525(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate1526(.a(gate168inter12), .b(gate168inter1), .O(G585));
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate743(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate744(.a(gate172inter0), .b(s_28), .O(gate172inter1));
  and2  gate745(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate746(.a(s_28), .O(gate172inter3));
  inv1  gate747(.a(s_29), .O(gate172inter4));
  nand2 gate748(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate749(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate750(.a(G483), .O(gate172inter7));
  inv1  gate751(.a(G549), .O(gate172inter8));
  nand2 gate752(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate753(.a(s_29), .b(gate172inter3), .O(gate172inter10));
  nor2  gate754(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate755(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate756(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate1597(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate1598(.a(gate175inter0), .b(s_150), .O(gate175inter1));
  and2  gate1599(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate1600(.a(s_150), .O(gate175inter3));
  inv1  gate1601(.a(s_151), .O(gate175inter4));
  nand2 gate1602(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1603(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1604(.a(G492), .O(gate175inter7));
  inv1  gate1605(.a(G555), .O(gate175inter8));
  nand2 gate1606(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1607(.a(s_151), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1608(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1609(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1610(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate967(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate968(.a(gate185inter0), .b(s_60), .O(gate185inter1));
  and2  gate969(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate970(.a(s_60), .O(gate185inter3));
  inv1  gate971(.a(s_61), .O(gate185inter4));
  nand2 gate972(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate973(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate974(.a(G570), .O(gate185inter7));
  inv1  gate975(.a(G571), .O(gate185inter8));
  nand2 gate976(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate977(.a(s_61), .b(gate185inter3), .O(gate185inter10));
  nor2  gate978(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate979(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate980(.a(gate185inter12), .b(gate185inter1), .O(G602));
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );

  xor2  gate1863(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate1864(.a(gate189inter0), .b(s_188), .O(gate189inter1));
  and2  gate1865(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate1866(.a(s_188), .O(gate189inter3));
  inv1  gate1867(.a(s_189), .O(gate189inter4));
  nand2 gate1868(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate1869(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate1870(.a(G578), .O(gate189inter7));
  inv1  gate1871(.a(G579), .O(gate189inter8));
  nand2 gate1872(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate1873(.a(s_189), .b(gate189inter3), .O(gate189inter10));
  nor2  gate1874(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate1875(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate1876(.a(gate189inter12), .b(gate189inter1), .O(G622));
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate1037(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate1038(.a(gate191inter0), .b(s_70), .O(gate191inter1));
  and2  gate1039(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate1040(.a(s_70), .O(gate191inter3));
  inv1  gate1041(.a(s_71), .O(gate191inter4));
  nand2 gate1042(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate1043(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate1044(.a(G582), .O(gate191inter7));
  inv1  gate1045(.a(G583), .O(gate191inter8));
  nand2 gate1046(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate1047(.a(s_71), .b(gate191inter3), .O(gate191inter10));
  nor2  gate1048(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate1049(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate1050(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate1653(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate1654(.a(gate195inter0), .b(s_158), .O(gate195inter1));
  and2  gate1655(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate1656(.a(s_158), .O(gate195inter3));
  inv1  gate1657(.a(s_159), .O(gate195inter4));
  nand2 gate1658(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate1659(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate1660(.a(G590), .O(gate195inter7));
  inv1  gate1661(.a(G591), .O(gate195inter8));
  nand2 gate1662(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate1663(.a(s_159), .b(gate195inter3), .O(gate195inter10));
  nor2  gate1664(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate1665(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate1666(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );

  xor2  gate981(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate982(.a(gate199inter0), .b(s_62), .O(gate199inter1));
  and2  gate983(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate984(.a(s_62), .O(gate199inter3));
  inv1  gate985(.a(s_63), .O(gate199inter4));
  nand2 gate986(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate987(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate988(.a(G598), .O(gate199inter7));
  inv1  gate989(.a(G599), .O(gate199inter8));
  nand2 gate990(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate991(.a(s_63), .b(gate199inter3), .O(gate199inter10));
  nor2  gate992(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate993(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate994(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate659(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate660(.a(gate201inter0), .b(s_16), .O(gate201inter1));
  and2  gate661(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate662(.a(s_16), .O(gate201inter3));
  inv1  gate663(.a(s_17), .O(gate201inter4));
  nand2 gate664(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate665(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate666(.a(G602), .O(gate201inter7));
  inv1  gate667(.a(G607), .O(gate201inter8));
  nand2 gate668(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate669(.a(s_17), .b(gate201inter3), .O(gate201inter10));
  nor2  gate670(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate671(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate672(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );

  xor2  gate841(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate842(.a(gate209inter0), .b(s_42), .O(gate209inter1));
  and2  gate843(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate844(.a(s_42), .O(gate209inter3));
  inv1  gate845(.a(s_43), .O(gate209inter4));
  nand2 gate846(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate847(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate848(.a(G602), .O(gate209inter7));
  inv1  gate849(.a(G666), .O(gate209inter8));
  nand2 gate850(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate851(.a(s_43), .b(gate209inter3), .O(gate209inter10));
  nor2  gate852(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate853(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate854(.a(gate209inter12), .b(gate209inter1), .O(G690));
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate1765(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate1766(.a(gate216inter0), .b(s_174), .O(gate216inter1));
  and2  gate1767(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate1768(.a(s_174), .O(gate216inter3));
  inv1  gate1769(.a(s_175), .O(gate216inter4));
  nand2 gate1770(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate1771(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate1772(.a(G617), .O(gate216inter7));
  inv1  gate1773(.a(G675), .O(gate216inter8));
  nand2 gate1774(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate1775(.a(s_175), .b(gate216inter3), .O(gate216inter10));
  nor2  gate1776(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate1777(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate1778(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate547(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate548(.a(gate218inter0), .b(s_0), .O(gate218inter1));
  and2  gate549(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate550(.a(s_0), .O(gate218inter3));
  inv1  gate551(.a(s_1), .O(gate218inter4));
  nand2 gate552(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate553(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate554(.a(G627), .O(gate218inter7));
  inv1  gate555(.a(G678), .O(gate218inter8));
  nand2 gate556(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate557(.a(s_1), .b(gate218inter3), .O(gate218inter10));
  nor2  gate558(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate559(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate560(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );

  xor2  gate1569(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate1570(.a(gate222inter0), .b(s_146), .O(gate222inter1));
  and2  gate1571(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate1572(.a(s_146), .O(gate222inter3));
  inv1  gate1573(.a(s_147), .O(gate222inter4));
  nand2 gate1574(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate1575(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate1576(.a(G632), .O(gate222inter7));
  inv1  gate1577(.a(G684), .O(gate222inter8));
  nand2 gate1578(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate1579(.a(s_147), .b(gate222inter3), .O(gate222inter10));
  nor2  gate1580(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate1581(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate1582(.a(gate222inter12), .b(gate222inter1), .O(G703));
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );

  xor2  gate1303(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate1304(.a(gate225inter0), .b(s_108), .O(gate225inter1));
  and2  gate1305(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate1306(.a(s_108), .O(gate225inter3));
  inv1  gate1307(.a(s_109), .O(gate225inter4));
  nand2 gate1308(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate1309(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate1310(.a(G690), .O(gate225inter7));
  inv1  gate1311(.a(G691), .O(gate225inter8));
  nand2 gate1312(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate1313(.a(s_109), .b(gate225inter3), .O(gate225inter10));
  nor2  gate1314(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate1315(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate1316(.a(gate225inter12), .b(gate225inter1), .O(G706));
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate1051(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate1052(.a(gate231inter0), .b(s_72), .O(gate231inter1));
  and2  gate1053(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate1054(.a(s_72), .O(gate231inter3));
  inv1  gate1055(.a(s_73), .O(gate231inter4));
  nand2 gate1056(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate1057(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate1058(.a(G702), .O(gate231inter7));
  inv1  gate1059(.a(G703), .O(gate231inter8));
  nand2 gate1060(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate1061(.a(s_73), .b(gate231inter3), .O(gate231inter10));
  nor2  gate1062(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate1063(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate1064(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate925(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate926(.a(gate236inter0), .b(s_54), .O(gate236inter1));
  and2  gate927(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate928(.a(s_54), .O(gate236inter3));
  inv1  gate929(.a(s_55), .O(gate236inter4));
  nand2 gate930(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate931(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate932(.a(G251), .O(gate236inter7));
  inv1  gate933(.a(G727), .O(gate236inter8));
  nand2 gate934(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate935(.a(s_55), .b(gate236inter3), .O(gate236inter10));
  nor2  gate936(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate937(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate938(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate2017(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate2018(.a(gate240inter0), .b(s_210), .O(gate240inter1));
  and2  gate2019(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate2020(.a(s_210), .O(gate240inter3));
  inv1  gate2021(.a(s_211), .O(gate240inter4));
  nand2 gate2022(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate2023(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate2024(.a(G263), .O(gate240inter7));
  inv1  gate2025(.a(G715), .O(gate240inter8));
  nand2 gate2026(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate2027(.a(s_211), .b(gate240inter3), .O(gate240inter10));
  nor2  gate2028(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate2029(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate2030(.a(gate240inter12), .b(gate240inter1), .O(G751));

  xor2  gate1359(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate1360(.a(gate241inter0), .b(s_116), .O(gate241inter1));
  and2  gate1361(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate1362(.a(s_116), .O(gate241inter3));
  inv1  gate1363(.a(s_117), .O(gate241inter4));
  nand2 gate1364(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate1365(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate1366(.a(G242), .O(gate241inter7));
  inv1  gate1367(.a(G730), .O(gate241inter8));
  nand2 gate1368(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate1369(.a(s_117), .b(gate241inter3), .O(gate241inter10));
  nor2  gate1370(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate1371(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate1372(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate1947(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1948(.a(gate243inter0), .b(s_200), .O(gate243inter1));
  and2  gate1949(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1950(.a(s_200), .O(gate243inter3));
  inv1  gate1951(.a(s_201), .O(gate243inter4));
  nand2 gate1952(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1953(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1954(.a(G245), .O(gate243inter7));
  inv1  gate1955(.a(G733), .O(gate243inter8));
  nand2 gate1956(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1957(.a(s_201), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1958(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1959(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1960(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate1429(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate1430(.a(gate248inter0), .b(s_126), .O(gate248inter1));
  and2  gate1431(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate1432(.a(s_126), .O(gate248inter3));
  inv1  gate1433(.a(s_127), .O(gate248inter4));
  nand2 gate1434(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate1435(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate1436(.a(G727), .O(gate248inter7));
  inv1  gate1437(.a(G739), .O(gate248inter8));
  nand2 gate1438(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate1439(.a(s_127), .b(gate248inter3), .O(gate248inter10));
  nor2  gate1440(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate1441(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate1442(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate1485(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate1486(.a(gate250inter0), .b(s_134), .O(gate250inter1));
  and2  gate1487(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate1488(.a(s_134), .O(gate250inter3));
  inv1  gate1489(.a(s_135), .O(gate250inter4));
  nand2 gate1490(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate1491(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate1492(.a(G706), .O(gate250inter7));
  inv1  gate1493(.a(G742), .O(gate250inter8));
  nand2 gate1494(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate1495(.a(s_135), .b(gate250inter3), .O(gate250inter10));
  nor2  gate1496(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate1497(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate1498(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate1415(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate1416(.a(gate252inter0), .b(s_124), .O(gate252inter1));
  and2  gate1417(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate1418(.a(s_124), .O(gate252inter3));
  inv1  gate1419(.a(s_125), .O(gate252inter4));
  nand2 gate1420(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate1421(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate1422(.a(G709), .O(gate252inter7));
  inv1  gate1423(.a(G745), .O(gate252inter8));
  nand2 gate1424(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate1425(.a(s_125), .b(gate252inter3), .O(gate252inter10));
  nor2  gate1426(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate1427(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate1428(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate855(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate856(.a(gate258inter0), .b(s_44), .O(gate258inter1));
  and2  gate857(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate858(.a(s_44), .O(gate258inter3));
  inv1  gate859(.a(s_45), .O(gate258inter4));
  nand2 gate860(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate861(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate862(.a(G756), .O(gate258inter7));
  inv1  gate863(.a(G757), .O(gate258inter8));
  nand2 gate864(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate865(.a(s_45), .b(gate258inter3), .O(gate258inter10));
  nor2  gate866(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate867(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate868(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate1667(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate1668(.a(gate263inter0), .b(s_160), .O(gate263inter1));
  and2  gate1669(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate1670(.a(s_160), .O(gate263inter3));
  inv1  gate1671(.a(s_161), .O(gate263inter4));
  nand2 gate1672(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate1673(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate1674(.a(G766), .O(gate263inter7));
  inv1  gate1675(.a(G767), .O(gate263inter8));
  nand2 gate1676(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate1677(.a(s_161), .b(gate263inter3), .O(gate263inter10));
  nor2  gate1678(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate1679(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate1680(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate1373(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate1374(.a(gate265inter0), .b(s_118), .O(gate265inter1));
  and2  gate1375(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate1376(.a(s_118), .O(gate265inter3));
  inv1  gate1377(.a(s_119), .O(gate265inter4));
  nand2 gate1378(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate1379(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate1380(.a(G642), .O(gate265inter7));
  inv1  gate1381(.a(G770), .O(gate265inter8));
  nand2 gate1382(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate1383(.a(s_119), .b(gate265inter3), .O(gate265inter10));
  nor2  gate1384(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate1385(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate1386(.a(gate265inter12), .b(gate265inter1), .O(G794));
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate589(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate590(.a(gate270inter0), .b(s_6), .O(gate270inter1));
  and2  gate591(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate592(.a(s_6), .O(gate270inter3));
  inv1  gate593(.a(s_7), .O(gate270inter4));
  nand2 gate594(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate595(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate596(.a(G657), .O(gate270inter7));
  inv1  gate597(.a(G785), .O(gate270inter8));
  nand2 gate598(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate599(.a(s_7), .b(gate270inter3), .O(gate270inter10));
  nor2  gate600(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate601(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate602(.a(gate270inter12), .b(gate270inter1), .O(G809));

  xor2  gate603(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate604(.a(gate271inter0), .b(s_8), .O(gate271inter1));
  and2  gate605(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate606(.a(s_8), .O(gate271inter3));
  inv1  gate607(.a(s_9), .O(gate271inter4));
  nand2 gate608(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate609(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate610(.a(G660), .O(gate271inter7));
  inv1  gate611(.a(G788), .O(gate271inter8));
  nand2 gate612(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate613(.a(s_9), .b(gate271inter3), .O(gate271inter10));
  nor2  gate614(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate615(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate616(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate827(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate828(.a(gate286inter0), .b(s_40), .O(gate286inter1));
  and2  gate829(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate830(.a(s_40), .O(gate286inter3));
  inv1  gate831(.a(s_41), .O(gate286inter4));
  nand2 gate832(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate833(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate834(.a(G788), .O(gate286inter7));
  inv1  gate835(.a(G812), .O(gate286inter8));
  nand2 gate836(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate837(.a(s_41), .b(gate286inter3), .O(gate286inter10));
  nor2  gate838(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate839(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate840(.a(gate286inter12), .b(gate286inter1), .O(G831));
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );

  xor2  gate1079(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate1080(.a(gate289inter0), .b(s_76), .O(gate289inter1));
  and2  gate1081(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate1082(.a(s_76), .O(gate289inter3));
  inv1  gate1083(.a(s_77), .O(gate289inter4));
  nand2 gate1084(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate1085(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate1086(.a(G818), .O(gate289inter7));
  inv1  gate1087(.a(G819), .O(gate289inter8));
  nand2 gate1088(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate1089(.a(s_77), .b(gate289inter3), .O(gate289inter10));
  nor2  gate1090(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate1091(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate1092(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate729(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate730(.a(gate389inter0), .b(s_26), .O(gate389inter1));
  and2  gate731(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate732(.a(s_26), .O(gate389inter3));
  inv1  gate733(.a(s_27), .O(gate389inter4));
  nand2 gate734(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate735(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate736(.a(G3), .O(gate389inter7));
  inv1  gate737(.a(G1042), .O(gate389inter8));
  nand2 gate738(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate739(.a(s_27), .b(gate389inter3), .O(gate389inter10));
  nor2  gate740(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate741(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate742(.a(gate389inter12), .b(gate389inter1), .O(G1138));

  xor2  gate785(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate786(.a(gate390inter0), .b(s_34), .O(gate390inter1));
  and2  gate787(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate788(.a(s_34), .O(gate390inter3));
  inv1  gate789(.a(s_35), .O(gate390inter4));
  nand2 gate790(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate791(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate792(.a(G4), .O(gate390inter7));
  inv1  gate793(.a(G1045), .O(gate390inter8));
  nand2 gate794(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate795(.a(s_35), .b(gate390inter3), .O(gate390inter10));
  nor2  gate796(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate797(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate798(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate1709(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1710(.a(gate395inter0), .b(s_166), .O(gate395inter1));
  and2  gate1711(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1712(.a(s_166), .O(gate395inter3));
  inv1  gate1713(.a(s_167), .O(gate395inter4));
  nand2 gate1714(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1715(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1716(.a(G9), .O(gate395inter7));
  inv1  gate1717(.a(G1060), .O(gate395inter8));
  nand2 gate1718(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1719(.a(s_167), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1720(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1721(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1722(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate813(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate814(.a(gate397inter0), .b(s_38), .O(gate397inter1));
  and2  gate815(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate816(.a(s_38), .O(gate397inter3));
  inv1  gate817(.a(s_39), .O(gate397inter4));
  nand2 gate818(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate819(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate820(.a(G11), .O(gate397inter7));
  inv1  gate821(.a(G1066), .O(gate397inter8));
  nand2 gate822(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate823(.a(s_39), .b(gate397inter3), .O(gate397inter10));
  nor2  gate824(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate825(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate826(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate673(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate674(.a(gate400inter0), .b(s_18), .O(gate400inter1));
  and2  gate675(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate676(.a(s_18), .O(gate400inter3));
  inv1  gate677(.a(s_19), .O(gate400inter4));
  nand2 gate678(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate679(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate680(.a(G14), .O(gate400inter7));
  inv1  gate681(.a(G1075), .O(gate400inter8));
  nand2 gate682(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate683(.a(s_19), .b(gate400inter3), .O(gate400inter10));
  nor2  gate684(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate685(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate686(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );

  xor2  gate1149(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate1150(.a(gate405inter0), .b(s_86), .O(gate405inter1));
  and2  gate1151(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate1152(.a(s_86), .O(gate405inter3));
  inv1  gate1153(.a(s_87), .O(gate405inter4));
  nand2 gate1154(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate1155(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate1156(.a(G19), .O(gate405inter7));
  inv1  gate1157(.a(G1090), .O(gate405inter8));
  nand2 gate1158(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate1159(.a(s_87), .b(gate405inter3), .O(gate405inter10));
  nor2  gate1160(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate1161(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate1162(.a(gate405inter12), .b(gate405inter1), .O(G1186));
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate1471(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate1472(.a(gate409inter0), .b(s_132), .O(gate409inter1));
  and2  gate1473(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate1474(.a(s_132), .O(gate409inter3));
  inv1  gate1475(.a(s_133), .O(gate409inter4));
  nand2 gate1476(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate1477(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate1478(.a(G23), .O(gate409inter7));
  inv1  gate1479(.a(G1102), .O(gate409inter8));
  nand2 gate1480(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate1481(.a(s_133), .b(gate409inter3), .O(gate409inter10));
  nor2  gate1482(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate1483(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate1484(.a(gate409inter12), .b(gate409inter1), .O(G1198));
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate1639(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate1640(.a(gate411inter0), .b(s_156), .O(gate411inter1));
  and2  gate1641(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate1642(.a(s_156), .O(gate411inter3));
  inv1  gate1643(.a(s_157), .O(gate411inter4));
  nand2 gate1644(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate1645(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate1646(.a(G25), .O(gate411inter7));
  inv1  gate1647(.a(G1108), .O(gate411inter8));
  nand2 gate1648(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate1649(.a(s_157), .b(gate411inter3), .O(gate411inter10));
  nor2  gate1650(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate1651(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate1652(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate1555(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1556(.a(gate420inter0), .b(s_144), .O(gate420inter1));
  and2  gate1557(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1558(.a(s_144), .O(gate420inter3));
  inv1  gate1559(.a(s_145), .O(gate420inter4));
  nand2 gate1560(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1561(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1562(.a(G1036), .O(gate420inter7));
  inv1  gate1563(.a(G1132), .O(gate420inter8));
  nand2 gate1564(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1565(.a(s_145), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1566(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1567(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1568(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );

  xor2  gate631(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate632(.a(gate423inter0), .b(s_12), .O(gate423inter1));
  and2  gate633(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate634(.a(s_12), .O(gate423inter3));
  inv1  gate635(.a(s_13), .O(gate423inter4));
  nand2 gate636(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate637(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate638(.a(G3), .O(gate423inter7));
  inv1  gate639(.a(G1138), .O(gate423inter8));
  nand2 gate640(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate641(.a(s_13), .b(gate423inter3), .O(gate423inter10));
  nor2  gate642(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate643(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate644(.a(gate423inter12), .b(gate423inter1), .O(G1232));

  xor2  gate1821(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate1822(.a(gate424inter0), .b(s_182), .O(gate424inter1));
  and2  gate1823(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate1824(.a(s_182), .O(gate424inter3));
  inv1  gate1825(.a(s_183), .O(gate424inter4));
  nand2 gate1826(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate1827(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate1828(.a(G1042), .O(gate424inter7));
  inv1  gate1829(.a(G1138), .O(gate424inter8));
  nand2 gate1830(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate1831(.a(s_183), .b(gate424inter3), .O(gate424inter10));
  nor2  gate1832(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate1833(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate1834(.a(gate424inter12), .b(gate424inter1), .O(G1233));

  xor2  gate1961(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate1962(.a(gate425inter0), .b(s_202), .O(gate425inter1));
  and2  gate1963(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate1964(.a(s_202), .O(gate425inter3));
  inv1  gate1965(.a(s_203), .O(gate425inter4));
  nand2 gate1966(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1967(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1968(.a(G4), .O(gate425inter7));
  inv1  gate1969(.a(G1141), .O(gate425inter8));
  nand2 gate1970(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1971(.a(s_203), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1972(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1973(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1974(.a(gate425inter12), .b(gate425inter1), .O(G1234));

  xor2  gate939(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate940(.a(gate426inter0), .b(s_56), .O(gate426inter1));
  and2  gate941(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate942(.a(s_56), .O(gate426inter3));
  inv1  gate943(.a(s_57), .O(gate426inter4));
  nand2 gate944(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate945(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate946(.a(G1045), .O(gate426inter7));
  inv1  gate947(.a(G1141), .O(gate426inter8));
  nand2 gate948(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate949(.a(s_57), .b(gate426inter3), .O(gate426inter10));
  nor2  gate950(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate951(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate952(.a(gate426inter12), .b(gate426inter1), .O(G1235));

  xor2  gate1163(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate1164(.a(gate427inter0), .b(s_88), .O(gate427inter1));
  and2  gate1165(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate1166(.a(s_88), .O(gate427inter3));
  inv1  gate1167(.a(s_89), .O(gate427inter4));
  nand2 gate1168(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate1169(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate1170(.a(G5), .O(gate427inter7));
  inv1  gate1171(.a(G1144), .O(gate427inter8));
  nand2 gate1172(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate1173(.a(s_89), .b(gate427inter3), .O(gate427inter10));
  nor2  gate1174(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate1175(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate1176(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate883(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate884(.a(gate430inter0), .b(s_48), .O(gate430inter1));
  and2  gate885(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate886(.a(s_48), .O(gate430inter3));
  inv1  gate887(.a(s_49), .O(gate430inter4));
  nand2 gate888(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate889(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate890(.a(G1051), .O(gate430inter7));
  inv1  gate891(.a(G1147), .O(gate430inter8));
  nand2 gate892(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate893(.a(s_49), .b(gate430inter3), .O(gate430inter10));
  nor2  gate894(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate895(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate896(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate645(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate646(.a(gate445inter0), .b(s_14), .O(gate445inter1));
  and2  gate647(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate648(.a(s_14), .O(gate445inter3));
  inv1  gate649(.a(s_15), .O(gate445inter4));
  nand2 gate650(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate651(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate652(.a(G14), .O(gate445inter7));
  inv1  gate653(.a(G1171), .O(gate445inter8));
  nand2 gate654(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate655(.a(s_15), .b(gate445inter3), .O(gate445inter10));
  nor2  gate656(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate657(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate658(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );

  xor2  gate1751(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate1752(.a(gate455inter0), .b(s_172), .O(gate455inter1));
  and2  gate1753(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate1754(.a(s_172), .O(gate455inter3));
  inv1  gate1755(.a(s_173), .O(gate455inter4));
  nand2 gate1756(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate1757(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate1758(.a(G19), .O(gate455inter7));
  inv1  gate1759(.a(G1186), .O(gate455inter8));
  nand2 gate1760(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate1761(.a(s_173), .b(gate455inter3), .O(gate455inter10));
  nor2  gate1762(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate1763(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate1764(.a(gate455inter12), .b(gate455inter1), .O(G1264));

  xor2  gate1443(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate1444(.a(gate456inter0), .b(s_128), .O(gate456inter1));
  and2  gate1445(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate1446(.a(s_128), .O(gate456inter3));
  inv1  gate1447(.a(s_129), .O(gate456inter4));
  nand2 gate1448(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate1449(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate1450(.a(G1090), .O(gate456inter7));
  inv1  gate1451(.a(G1186), .O(gate456inter8));
  nand2 gate1452(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate1453(.a(s_129), .b(gate456inter3), .O(gate456inter10));
  nor2  gate1454(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate1455(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate1456(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );

  xor2  gate1219(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate1220(.a(gate458inter0), .b(s_96), .O(gate458inter1));
  and2  gate1221(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate1222(.a(s_96), .O(gate458inter3));
  inv1  gate1223(.a(s_97), .O(gate458inter4));
  nand2 gate1224(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate1225(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate1226(.a(G1093), .O(gate458inter7));
  inv1  gate1227(.a(G1189), .O(gate458inter8));
  nand2 gate1228(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate1229(.a(s_97), .b(gate458inter3), .O(gate458inter10));
  nor2  gate1230(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate1231(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate1232(.a(gate458inter12), .b(gate458inter1), .O(G1267));

  xor2  gate715(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate716(.a(gate459inter0), .b(s_24), .O(gate459inter1));
  and2  gate717(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate718(.a(s_24), .O(gate459inter3));
  inv1  gate719(.a(s_25), .O(gate459inter4));
  nand2 gate720(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate721(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate722(.a(G21), .O(gate459inter7));
  inv1  gate723(.a(G1192), .O(gate459inter8));
  nand2 gate724(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate725(.a(s_25), .b(gate459inter3), .O(gate459inter10));
  nor2  gate726(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate727(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate728(.a(gate459inter12), .b(gate459inter1), .O(G1268));

  xor2  gate561(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate562(.a(gate460inter0), .b(s_2), .O(gate460inter1));
  and2  gate563(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate564(.a(s_2), .O(gate460inter3));
  inv1  gate565(.a(s_3), .O(gate460inter4));
  nand2 gate566(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate567(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate568(.a(G1096), .O(gate460inter7));
  inv1  gate569(.a(G1192), .O(gate460inter8));
  nand2 gate570(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate571(.a(s_3), .b(gate460inter3), .O(gate460inter10));
  nor2  gate572(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate573(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate574(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate771(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate772(.a(gate465inter0), .b(s_32), .O(gate465inter1));
  and2  gate773(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate774(.a(s_32), .O(gate465inter3));
  inv1  gate775(.a(s_33), .O(gate465inter4));
  nand2 gate776(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate777(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate778(.a(G24), .O(gate465inter7));
  inv1  gate779(.a(G1201), .O(gate465inter8));
  nand2 gate780(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate781(.a(s_33), .b(gate465inter3), .O(gate465inter10));
  nor2  gate782(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate783(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate784(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );

  xor2  gate897(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate898(.a(gate467inter0), .b(s_50), .O(gate467inter1));
  and2  gate899(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate900(.a(s_50), .O(gate467inter3));
  inv1  gate901(.a(s_51), .O(gate467inter4));
  nand2 gate902(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate903(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate904(.a(G25), .O(gate467inter7));
  inv1  gate905(.a(G1204), .O(gate467inter8));
  nand2 gate906(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate907(.a(s_51), .b(gate467inter3), .O(gate467inter10));
  nor2  gate908(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate909(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate910(.a(gate467inter12), .b(gate467inter1), .O(G1276));

  xor2  gate1807(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate1808(.a(gate468inter0), .b(s_180), .O(gate468inter1));
  and2  gate1809(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate1810(.a(s_180), .O(gate468inter3));
  inv1  gate1811(.a(s_181), .O(gate468inter4));
  nand2 gate1812(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate1813(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate1814(.a(G1108), .O(gate468inter7));
  inv1  gate1815(.a(G1204), .O(gate468inter8));
  nand2 gate1816(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate1817(.a(s_181), .b(gate468inter3), .O(gate468inter10));
  nor2  gate1818(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate1819(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate1820(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );

  xor2  gate1135(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate1136(.a(gate470inter0), .b(s_84), .O(gate470inter1));
  and2  gate1137(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate1138(.a(s_84), .O(gate470inter3));
  inv1  gate1139(.a(s_85), .O(gate470inter4));
  nand2 gate1140(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate1141(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate1142(.a(G1111), .O(gate470inter7));
  inv1  gate1143(.a(G1207), .O(gate470inter8));
  nand2 gate1144(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate1145(.a(s_85), .b(gate470inter3), .O(gate470inter10));
  nor2  gate1146(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate1147(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate1148(.a(gate470inter12), .b(gate470inter1), .O(G1279));

  xor2  gate1737(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate1738(.a(gate471inter0), .b(s_170), .O(gate471inter1));
  and2  gate1739(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate1740(.a(s_170), .O(gate471inter3));
  inv1  gate1741(.a(s_171), .O(gate471inter4));
  nand2 gate1742(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate1743(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate1744(.a(G27), .O(gate471inter7));
  inv1  gate1745(.a(G1210), .O(gate471inter8));
  nand2 gate1746(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate1747(.a(s_171), .b(gate471inter3), .O(gate471inter10));
  nor2  gate1748(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate1749(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate1750(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );

  xor2  gate1205(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate1206(.a(gate473inter0), .b(s_94), .O(gate473inter1));
  and2  gate1207(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate1208(.a(s_94), .O(gate473inter3));
  inv1  gate1209(.a(s_95), .O(gate473inter4));
  nand2 gate1210(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate1211(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate1212(.a(G28), .O(gate473inter7));
  inv1  gate1213(.a(G1213), .O(gate473inter8));
  nand2 gate1214(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate1215(.a(s_95), .b(gate473inter3), .O(gate473inter10));
  nor2  gate1216(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate1217(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate1218(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate1177(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate1178(.a(gate475inter0), .b(s_90), .O(gate475inter1));
  and2  gate1179(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate1180(.a(s_90), .O(gate475inter3));
  inv1  gate1181(.a(s_91), .O(gate475inter4));
  nand2 gate1182(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate1183(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate1184(.a(G29), .O(gate475inter7));
  inv1  gate1185(.a(G1216), .O(gate475inter8));
  nand2 gate1186(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate1187(.a(s_91), .b(gate475inter3), .O(gate475inter10));
  nor2  gate1188(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate1189(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate1190(.a(gate475inter12), .b(gate475inter1), .O(G1284));
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );

  xor2  gate1625(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate1626(.a(gate483inter0), .b(s_154), .O(gate483inter1));
  and2  gate1627(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate1628(.a(s_154), .O(gate483inter3));
  inv1  gate1629(.a(s_155), .O(gate483inter4));
  nand2 gate1630(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate1631(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate1632(.a(G1228), .O(gate483inter7));
  inv1  gate1633(.a(G1229), .O(gate483inter8));
  nand2 gate1634(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate1635(.a(s_155), .b(gate483inter3), .O(gate483inter10));
  nor2  gate1636(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate1637(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate1638(.a(gate483inter12), .b(gate483inter1), .O(G1292));

  xor2  gate1905(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate1906(.a(gate484inter0), .b(s_194), .O(gate484inter1));
  and2  gate1907(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate1908(.a(s_194), .O(gate484inter3));
  inv1  gate1909(.a(s_195), .O(gate484inter4));
  nand2 gate1910(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate1911(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate1912(.a(G1230), .O(gate484inter7));
  inv1  gate1913(.a(G1231), .O(gate484inter8));
  nand2 gate1914(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate1915(.a(s_195), .b(gate484inter3), .O(gate484inter10));
  nor2  gate1916(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate1917(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate1918(.a(gate484inter12), .b(gate484inter1), .O(G1293));
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate953(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate954(.a(gate486inter0), .b(s_58), .O(gate486inter1));
  and2  gate955(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate956(.a(s_58), .O(gate486inter3));
  inv1  gate957(.a(s_59), .O(gate486inter4));
  nand2 gate958(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate959(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate960(.a(G1234), .O(gate486inter7));
  inv1  gate961(.a(G1235), .O(gate486inter8));
  nand2 gate962(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate963(.a(s_59), .b(gate486inter3), .O(gate486inter10));
  nor2  gate964(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate965(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate966(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate1093(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate1094(.a(gate493inter0), .b(s_78), .O(gate493inter1));
  and2  gate1095(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate1096(.a(s_78), .O(gate493inter3));
  inv1  gate1097(.a(s_79), .O(gate493inter4));
  nand2 gate1098(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate1099(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate1100(.a(G1248), .O(gate493inter7));
  inv1  gate1101(.a(G1249), .O(gate493inter8));
  nand2 gate1102(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate1103(.a(s_79), .b(gate493inter3), .O(gate493inter10));
  nor2  gate1104(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate1105(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate1106(.a(gate493inter12), .b(gate493inter1), .O(G1302));
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );

  xor2  gate1499(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate1500(.a(gate495inter0), .b(s_136), .O(gate495inter1));
  and2  gate1501(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate1502(.a(s_136), .O(gate495inter3));
  inv1  gate1503(.a(s_137), .O(gate495inter4));
  nand2 gate1504(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate1505(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate1506(.a(G1252), .O(gate495inter7));
  inv1  gate1507(.a(G1253), .O(gate495inter8));
  nand2 gate1508(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate1509(.a(s_137), .b(gate495inter3), .O(gate495inter10));
  nor2  gate1510(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate1511(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate1512(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate1121(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate1122(.a(gate504inter0), .b(s_82), .O(gate504inter1));
  and2  gate1123(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate1124(.a(s_82), .O(gate504inter3));
  inv1  gate1125(.a(s_83), .O(gate504inter4));
  nand2 gate1126(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate1127(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate1128(.a(G1270), .O(gate504inter7));
  inv1  gate1129(.a(G1271), .O(gate504inter8));
  nand2 gate1130(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate1131(.a(s_83), .b(gate504inter3), .O(gate504inter10));
  nor2  gate1132(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate1133(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate1134(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate1793(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate1794(.a(gate511inter0), .b(s_178), .O(gate511inter1));
  and2  gate1795(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate1796(.a(s_178), .O(gate511inter3));
  inv1  gate1797(.a(s_179), .O(gate511inter4));
  nand2 gate1798(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate1799(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate1800(.a(G1284), .O(gate511inter7));
  inv1  gate1801(.a(G1285), .O(gate511inter8));
  nand2 gate1802(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate1803(.a(s_179), .b(gate511inter3), .O(gate511inter10));
  nor2  gate1804(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate1805(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate1806(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule