module c432 (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
             N430,N431,N432);
input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
      N99,N102,N105,N108,N112,N115;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91;
output N223,N329,N370,N421,N430,N431,N432;
wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate123inter0, gate123inter1, gate123inter2, gate123inter3, gate123inter4, gate123inter5, gate123inter6, gate123inter7, gate123inter8, gate123inter9, gate123inter10, gate123inter11, gate123inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12;


inv1 gate1( .a(N1), .O(N118) );
inv1 gate2( .a(N4), .O(N119) );
inv1 gate3( .a(N11), .O(N122) );
inv1 gate4( .a(N17), .O(N123) );
inv1 gate5( .a(N24), .O(N126) );
inv1 gate6( .a(N30), .O(N127) );
inv1 gate7( .a(N37), .O(N130) );
inv1 gate8( .a(N43), .O(N131) );
inv1 gate9( .a(N50), .O(N134) );
inv1 gate10( .a(N56), .O(N135) );
inv1 gate11( .a(N63), .O(N138) );
inv1 gate12( .a(N69), .O(N139) );
inv1 gate13( .a(N76), .O(N142) );
inv1 gate14( .a(N82), .O(N143) );
inv1 gate15( .a(N89), .O(N146) );
inv1 gate16( .a(N95), .O(N147) );
inv1 gate17( .a(N102), .O(N150) );
inv1 gate18( .a(N108), .O(N151) );

  xor2  gate455(.a(N4), .b(N118), .O(gate19inter0));
  nand2 gate456(.a(gate19inter0), .b(s_42), .O(gate19inter1));
  and2  gate457(.a(N4), .b(N118), .O(gate19inter2));
  inv1  gate458(.a(s_42), .O(gate19inter3));
  inv1  gate459(.a(s_43), .O(gate19inter4));
  nand2 gate460(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate461(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate462(.a(N118), .O(gate19inter7));
  inv1  gate463(.a(N4), .O(gate19inter8));
  nand2 gate464(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate465(.a(s_43), .b(gate19inter3), .O(gate19inter10));
  nor2  gate466(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate467(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate468(.a(gate19inter12), .b(gate19inter1), .O(N154));
nor2 gate20( .a(N8), .b(N119), .O(N157) );

  xor2  gate637(.a(N119), .b(N14), .O(gate21inter0));
  nand2 gate638(.a(gate21inter0), .b(s_68), .O(gate21inter1));
  and2  gate639(.a(N119), .b(N14), .O(gate21inter2));
  inv1  gate640(.a(s_68), .O(gate21inter3));
  inv1  gate641(.a(s_69), .O(gate21inter4));
  nand2 gate642(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate643(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate644(.a(N14), .O(gate21inter7));
  inv1  gate645(.a(N119), .O(gate21inter8));
  nand2 gate646(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate647(.a(s_69), .b(gate21inter3), .O(gate21inter10));
  nor2  gate648(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate649(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate650(.a(gate21inter12), .b(gate21inter1), .O(N158));

  xor2  gate189(.a(N17), .b(N122), .O(gate22inter0));
  nand2 gate190(.a(gate22inter0), .b(s_4), .O(gate22inter1));
  and2  gate191(.a(N17), .b(N122), .O(gate22inter2));
  inv1  gate192(.a(s_4), .O(gate22inter3));
  inv1  gate193(.a(s_5), .O(gate22inter4));
  nand2 gate194(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate195(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate196(.a(N122), .O(gate22inter7));
  inv1  gate197(.a(N17), .O(gate22inter8));
  nand2 gate198(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate199(.a(s_5), .b(gate22inter3), .O(gate22inter10));
  nor2  gate200(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate201(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate202(.a(gate22inter12), .b(gate22inter1), .O(N159));
nand2 gate23( .a(N126), .b(N30), .O(N162) );

  xor2  gate273(.a(N43), .b(N130), .O(gate24inter0));
  nand2 gate274(.a(gate24inter0), .b(s_16), .O(gate24inter1));
  and2  gate275(.a(N43), .b(N130), .O(gate24inter2));
  inv1  gate276(.a(s_16), .O(gate24inter3));
  inv1  gate277(.a(s_17), .O(gate24inter4));
  nand2 gate278(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate279(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate280(.a(N130), .O(gate24inter7));
  inv1  gate281(.a(N43), .O(gate24inter8));
  nand2 gate282(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate283(.a(s_17), .b(gate24inter3), .O(gate24inter10));
  nor2  gate284(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate285(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate286(.a(gate24inter12), .b(gate24inter1), .O(N165));
nand2 gate25( .a(N134), .b(N56), .O(N168) );

  xor2  gate707(.a(N69), .b(N138), .O(gate26inter0));
  nand2 gate708(.a(gate26inter0), .b(s_78), .O(gate26inter1));
  and2  gate709(.a(N69), .b(N138), .O(gate26inter2));
  inv1  gate710(.a(s_78), .O(gate26inter3));
  inv1  gate711(.a(s_79), .O(gate26inter4));
  nand2 gate712(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate713(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate714(.a(N138), .O(gate26inter7));
  inv1  gate715(.a(N69), .O(gate26inter8));
  nand2 gate716(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate717(.a(s_79), .b(gate26inter3), .O(gate26inter10));
  nor2  gate718(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate719(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate720(.a(gate26inter12), .b(gate26inter1), .O(N171));
nand2 gate27( .a(N142), .b(N82), .O(N174) );

  xor2  gate301(.a(N95), .b(N146), .O(gate28inter0));
  nand2 gate302(.a(gate28inter0), .b(s_20), .O(gate28inter1));
  and2  gate303(.a(N95), .b(N146), .O(gate28inter2));
  inv1  gate304(.a(s_20), .O(gate28inter3));
  inv1  gate305(.a(s_21), .O(gate28inter4));
  nand2 gate306(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate307(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate308(.a(N146), .O(gate28inter7));
  inv1  gate309(.a(N95), .O(gate28inter8));
  nand2 gate310(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate311(.a(s_21), .b(gate28inter3), .O(gate28inter10));
  nor2  gate312(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate313(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate314(.a(gate28inter12), .b(gate28inter1), .O(N177));

  xor2  gate343(.a(N108), .b(N150), .O(gate29inter0));
  nand2 gate344(.a(gate29inter0), .b(s_26), .O(gate29inter1));
  and2  gate345(.a(N108), .b(N150), .O(gate29inter2));
  inv1  gate346(.a(s_26), .O(gate29inter3));
  inv1  gate347(.a(s_27), .O(gate29inter4));
  nand2 gate348(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate349(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate350(.a(N150), .O(gate29inter7));
  inv1  gate351(.a(N108), .O(gate29inter8));
  nand2 gate352(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate353(.a(s_27), .b(gate29inter3), .O(gate29inter10));
  nor2  gate354(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate355(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate356(.a(gate29inter12), .b(gate29inter1), .O(N180));
nor2 gate30( .a(N21), .b(N123), .O(N183) );
nor2 gate31( .a(N27), .b(N123), .O(N184) );

  xor2  gate399(.a(N127), .b(N34), .O(gate32inter0));
  nand2 gate400(.a(gate32inter0), .b(s_34), .O(gate32inter1));
  and2  gate401(.a(N127), .b(N34), .O(gate32inter2));
  inv1  gate402(.a(s_34), .O(gate32inter3));
  inv1  gate403(.a(s_35), .O(gate32inter4));
  nand2 gate404(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate405(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate406(.a(N34), .O(gate32inter7));
  inv1  gate407(.a(N127), .O(gate32inter8));
  nand2 gate408(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate409(.a(s_35), .b(gate32inter3), .O(gate32inter10));
  nor2  gate410(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate411(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate412(.a(gate32inter12), .b(gate32inter1), .O(N185));
nor2 gate33( .a(N40), .b(N127), .O(N186) );

  xor2  gate525(.a(N131), .b(N47), .O(gate34inter0));
  nand2 gate526(.a(gate34inter0), .b(s_52), .O(gate34inter1));
  and2  gate527(.a(N131), .b(N47), .O(gate34inter2));
  inv1  gate528(.a(s_52), .O(gate34inter3));
  inv1  gate529(.a(s_53), .O(gate34inter4));
  nand2 gate530(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate531(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate532(.a(N47), .O(gate34inter7));
  inv1  gate533(.a(N131), .O(gate34inter8));
  nand2 gate534(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate535(.a(s_53), .b(gate34inter3), .O(gate34inter10));
  nor2  gate536(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate537(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate538(.a(gate34inter12), .b(gate34inter1), .O(N187));
nor2 gate35( .a(N53), .b(N131), .O(N188) );
nor2 gate36( .a(N60), .b(N135), .O(N189) );

  xor2  gate175(.a(N135), .b(N66), .O(gate37inter0));
  nand2 gate176(.a(gate37inter0), .b(s_2), .O(gate37inter1));
  and2  gate177(.a(N135), .b(N66), .O(gate37inter2));
  inv1  gate178(.a(s_2), .O(gate37inter3));
  inv1  gate179(.a(s_3), .O(gate37inter4));
  nand2 gate180(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate181(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate182(.a(N66), .O(gate37inter7));
  inv1  gate183(.a(N135), .O(gate37inter8));
  nand2 gate184(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate185(.a(s_3), .b(gate37inter3), .O(gate37inter10));
  nor2  gate186(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate187(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate188(.a(gate37inter12), .b(gate37inter1), .O(N190));
nor2 gate38( .a(N73), .b(N139), .O(N191) );
nor2 gate39( .a(N79), .b(N139), .O(N192) );

  xor2  gate259(.a(N143), .b(N86), .O(gate40inter0));
  nand2 gate260(.a(gate40inter0), .b(s_14), .O(gate40inter1));
  and2  gate261(.a(N143), .b(N86), .O(gate40inter2));
  inv1  gate262(.a(s_14), .O(gate40inter3));
  inv1  gate263(.a(s_15), .O(gate40inter4));
  nand2 gate264(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate265(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate266(.a(N86), .O(gate40inter7));
  inv1  gate267(.a(N143), .O(gate40inter8));
  nand2 gate268(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate269(.a(s_15), .b(gate40inter3), .O(gate40inter10));
  nor2  gate270(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate271(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate272(.a(gate40inter12), .b(gate40inter1), .O(N193));

  xor2  gate735(.a(N143), .b(N92), .O(gate41inter0));
  nand2 gate736(.a(gate41inter0), .b(s_82), .O(gate41inter1));
  and2  gate737(.a(N143), .b(N92), .O(gate41inter2));
  inv1  gate738(.a(s_82), .O(gate41inter3));
  inv1  gate739(.a(s_83), .O(gate41inter4));
  nand2 gate740(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate741(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate742(.a(N92), .O(gate41inter7));
  inv1  gate743(.a(N143), .O(gate41inter8));
  nand2 gate744(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate745(.a(s_83), .b(gate41inter3), .O(gate41inter10));
  nor2  gate746(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate747(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate748(.a(gate41inter12), .b(gate41inter1), .O(N194));

  xor2  gate315(.a(N147), .b(N99), .O(gate42inter0));
  nand2 gate316(.a(gate42inter0), .b(s_22), .O(gate42inter1));
  and2  gate317(.a(N147), .b(N99), .O(gate42inter2));
  inv1  gate318(.a(s_22), .O(gate42inter3));
  inv1  gate319(.a(s_23), .O(gate42inter4));
  nand2 gate320(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate321(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate322(.a(N99), .O(gate42inter7));
  inv1  gate323(.a(N147), .O(gate42inter8));
  nand2 gate324(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate325(.a(s_23), .b(gate42inter3), .O(gate42inter10));
  nor2  gate326(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate327(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate328(.a(gate42inter12), .b(gate42inter1), .O(N195));
nor2 gate43( .a(N105), .b(N147), .O(N196) );
nor2 gate44( .a(N112), .b(N151), .O(N197) );

  xor2  gate609(.a(N151), .b(N115), .O(gate45inter0));
  nand2 gate610(.a(gate45inter0), .b(s_64), .O(gate45inter1));
  and2  gate611(.a(N151), .b(N115), .O(gate45inter2));
  inv1  gate612(.a(s_64), .O(gate45inter3));
  inv1  gate613(.a(s_65), .O(gate45inter4));
  nand2 gate614(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate615(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate616(.a(N115), .O(gate45inter7));
  inv1  gate617(.a(N151), .O(gate45inter8));
  nand2 gate618(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate619(.a(s_65), .b(gate45inter3), .O(gate45inter10));
  nor2  gate620(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate621(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate622(.a(gate45inter12), .b(gate45inter1), .O(N198));
and9 gate46( .a(N154), .b(N159), .c(N162), .d(N165), .e(N168), .f(N171), .g(N174), .h(N177), .i(N180), .O(N199) );
inv1 gate47( .a(N199), .O(N203) );
inv1 gate48( .a(N199), .O(N213) );
inv1 gate49( .a(N199), .O(N223) );
xor2 gate50( .a(N203), .b(N154), .O(N224) );

  xor2  gate231(.a(N159), .b(N203), .O(gate51inter0));
  nand2 gate232(.a(gate51inter0), .b(s_10), .O(gate51inter1));
  and2  gate233(.a(N159), .b(N203), .O(gate51inter2));
  inv1  gate234(.a(s_10), .O(gate51inter3));
  inv1  gate235(.a(s_11), .O(gate51inter4));
  nand2 gate236(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate237(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate238(.a(N203), .O(gate51inter7));
  inv1  gate239(.a(N159), .O(gate51inter8));
  nand2 gate240(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate241(.a(s_11), .b(gate51inter3), .O(gate51inter10));
  nor2  gate242(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate243(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate244(.a(gate51inter12), .b(gate51inter1), .O(N227));
xor2 gate52( .a(N203), .b(N162), .O(N230) );

  xor2  gate721(.a(N165), .b(N203), .O(gate53inter0));
  nand2 gate722(.a(gate53inter0), .b(s_80), .O(gate53inter1));
  and2  gate723(.a(N165), .b(N203), .O(gate53inter2));
  inv1  gate724(.a(s_80), .O(gate53inter3));
  inv1  gate725(.a(s_81), .O(gate53inter4));
  nand2 gate726(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate727(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate728(.a(N203), .O(gate53inter7));
  inv1  gate729(.a(N165), .O(gate53inter8));
  nand2 gate730(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate731(.a(s_81), .b(gate53inter3), .O(gate53inter10));
  nor2  gate732(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate733(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate734(.a(gate53inter12), .b(gate53inter1), .O(N233));
xor2 gate54( .a(N203), .b(N168), .O(N236) );
xor2 gate55( .a(N203), .b(N171), .O(N239) );

  xor2  gate161(.a(N213), .b(N1), .O(gate56inter0));
  nand2 gate162(.a(gate56inter0), .b(s_0), .O(gate56inter1));
  and2  gate163(.a(N213), .b(N1), .O(gate56inter2));
  inv1  gate164(.a(s_0), .O(gate56inter3));
  inv1  gate165(.a(s_1), .O(gate56inter4));
  nand2 gate166(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate167(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate168(.a(N1), .O(gate56inter7));
  inv1  gate169(.a(N213), .O(gate56inter8));
  nand2 gate170(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate171(.a(s_1), .b(gate56inter3), .O(gate56inter10));
  nor2  gate172(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate173(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate174(.a(gate56inter12), .b(gate56inter1), .O(N242));
xor2 gate57( .a(N203), .b(N174), .O(N243) );
nand2 gate58( .a(N213), .b(N11), .O(N246) );

  xor2  gate763(.a(N177), .b(N203), .O(gate59inter0));
  nand2 gate764(.a(gate59inter0), .b(s_86), .O(gate59inter1));
  and2  gate765(.a(N177), .b(N203), .O(gate59inter2));
  inv1  gate766(.a(s_86), .O(gate59inter3));
  inv1  gate767(.a(s_87), .O(gate59inter4));
  nand2 gate768(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate769(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate770(.a(N203), .O(gate59inter7));
  inv1  gate771(.a(N177), .O(gate59inter8));
  nand2 gate772(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate773(.a(s_87), .b(gate59inter3), .O(gate59inter10));
  nor2  gate774(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate775(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate776(.a(gate59inter12), .b(gate59inter1), .O(N247));

  xor2  gate203(.a(N24), .b(N213), .O(gate60inter0));
  nand2 gate204(.a(gate60inter0), .b(s_6), .O(gate60inter1));
  and2  gate205(.a(N24), .b(N213), .O(gate60inter2));
  inv1  gate206(.a(s_6), .O(gate60inter3));
  inv1  gate207(.a(s_7), .O(gate60inter4));
  nand2 gate208(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate209(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate210(.a(N213), .O(gate60inter7));
  inv1  gate211(.a(N24), .O(gate60inter8));
  nand2 gate212(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate213(.a(s_7), .b(gate60inter3), .O(gate60inter10));
  nor2  gate214(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate215(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate216(.a(gate60inter12), .b(gate60inter1), .O(N250));
xor2 gate61( .a(N203), .b(N180), .O(N251) );
nand2 gate62( .a(N213), .b(N37), .O(N254) );
nand2 gate63( .a(N213), .b(N50), .O(N255) );
nand2 gate64( .a(N213), .b(N63), .O(N256) );

  xor2  gate287(.a(N76), .b(N213), .O(gate65inter0));
  nand2 gate288(.a(gate65inter0), .b(s_18), .O(gate65inter1));
  and2  gate289(.a(N76), .b(N213), .O(gate65inter2));
  inv1  gate290(.a(s_18), .O(gate65inter3));
  inv1  gate291(.a(s_19), .O(gate65inter4));
  nand2 gate292(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate293(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate294(.a(N213), .O(gate65inter7));
  inv1  gate295(.a(N76), .O(gate65inter8));
  nand2 gate296(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate297(.a(s_19), .b(gate65inter3), .O(gate65inter10));
  nor2  gate298(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate299(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate300(.a(gate65inter12), .b(gate65inter1), .O(N257));

  xor2  gate567(.a(N89), .b(N213), .O(gate66inter0));
  nand2 gate568(.a(gate66inter0), .b(s_58), .O(gate66inter1));
  and2  gate569(.a(N89), .b(N213), .O(gate66inter2));
  inv1  gate570(.a(s_58), .O(gate66inter3));
  inv1  gate571(.a(s_59), .O(gate66inter4));
  nand2 gate572(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate573(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate574(.a(N213), .O(gate66inter7));
  inv1  gate575(.a(N89), .O(gate66inter8));
  nand2 gate576(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate577(.a(s_59), .b(gate66inter3), .O(gate66inter10));
  nor2  gate578(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate579(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate580(.a(gate66inter12), .b(gate66inter1), .O(N258));

  xor2  gate539(.a(N102), .b(N213), .O(gate67inter0));
  nand2 gate540(.a(gate67inter0), .b(s_54), .O(gate67inter1));
  and2  gate541(.a(N102), .b(N213), .O(gate67inter2));
  inv1  gate542(.a(s_54), .O(gate67inter3));
  inv1  gate543(.a(s_55), .O(gate67inter4));
  nand2 gate544(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate545(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate546(.a(N213), .O(gate67inter7));
  inv1  gate547(.a(N102), .O(gate67inter8));
  nand2 gate548(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate549(.a(s_55), .b(gate67inter3), .O(gate67inter10));
  nor2  gate550(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate551(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate552(.a(gate67inter12), .b(gate67inter1), .O(N259));

  xor2  gate357(.a(N157), .b(N224), .O(gate68inter0));
  nand2 gate358(.a(gate68inter0), .b(s_28), .O(gate68inter1));
  and2  gate359(.a(N157), .b(N224), .O(gate68inter2));
  inv1  gate360(.a(s_28), .O(gate68inter3));
  inv1  gate361(.a(s_29), .O(gate68inter4));
  nand2 gate362(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate363(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate364(.a(N224), .O(gate68inter7));
  inv1  gate365(.a(N157), .O(gate68inter8));
  nand2 gate366(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate367(.a(s_29), .b(gate68inter3), .O(gate68inter10));
  nor2  gate368(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate369(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate370(.a(gate68inter12), .b(gate68inter1), .O(N260));
nand2 gate69( .a(N224), .b(N158), .O(N263) );
nand2 gate70( .a(N227), .b(N183), .O(N264) );
nand2 gate71( .a(N230), .b(N185), .O(N267) );

  xor2  gate497(.a(N187), .b(N233), .O(gate72inter0));
  nand2 gate498(.a(gate72inter0), .b(s_48), .O(gate72inter1));
  and2  gate499(.a(N187), .b(N233), .O(gate72inter2));
  inv1  gate500(.a(s_48), .O(gate72inter3));
  inv1  gate501(.a(s_49), .O(gate72inter4));
  nand2 gate502(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate503(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate504(.a(N233), .O(gate72inter7));
  inv1  gate505(.a(N187), .O(gate72inter8));
  nand2 gate506(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate507(.a(s_49), .b(gate72inter3), .O(gate72inter10));
  nor2  gate508(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate509(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate510(.a(gate72inter12), .b(gate72inter1), .O(N270));

  xor2  gate791(.a(N189), .b(N236), .O(gate73inter0));
  nand2 gate792(.a(gate73inter0), .b(s_90), .O(gate73inter1));
  and2  gate793(.a(N189), .b(N236), .O(gate73inter2));
  inv1  gate794(.a(s_90), .O(gate73inter3));
  inv1  gate795(.a(s_91), .O(gate73inter4));
  nand2 gate796(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate797(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate798(.a(N236), .O(gate73inter7));
  inv1  gate799(.a(N189), .O(gate73inter8));
  nand2 gate800(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate801(.a(s_91), .b(gate73inter3), .O(gate73inter10));
  nor2  gate802(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate803(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate804(.a(gate73inter12), .b(gate73inter1), .O(N273));

  xor2  gate679(.a(N191), .b(N239), .O(gate74inter0));
  nand2 gate680(.a(gate74inter0), .b(s_74), .O(gate74inter1));
  and2  gate681(.a(N191), .b(N239), .O(gate74inter2));
  inv1  gate682(.a(s_74), .O(gate74inter3));
  inv1  gate683(.a(s_75), .O(gate74inter4));
  nand2 gate684(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate685(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate686(.a(N239), .O(gate74inter7));
  inv1  gate687(.a(N191), .O(gate74inter8));
  nand2 gate688(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate689(.a(s_75), .b(gate74inter3), .O(gate74inter10));
  nor2  gate690(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate691(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate692(.a(gate74inter12), .b(gate74inter1), .O(N276));
nand2 gate75( .a(N243), .b(N193), .O(N279) );
nand2 gate76( .a(N247), .b(N195), .O(N282) );
nand2 gate77( .a(N251), .b(N197), .O(N285) );

  xor2  gate441(.a(N184), .b(N227), .O(gate78inter0));
  nand2 gate442(.a(gate78inter0), .b(s_40), .O(gate78inter1));
  and2  gate443(.a(N184), .b(N227), .O(gate78inter2));
  inv1  gate444(.a(s_40), .O(gate78inter3));
  inv1  gate445(.a(s_41), .O(gate78inter4));
  nand2 gate446(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate447(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate448(.a(N227), .O(gate78inter7));
  inv1  gate449(.a(N184), .O(gate78inter8));
  nand2 gate450(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate451(.a(s_41), .b(gate78inter3), .O(gate78inter10));
  nor2  gate452(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate453(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate454(.a(gate78inter12), .b(gate78inter1), .O(N288));

  xor2  gate665(.a(N186), .b(N230), .O(gate79inter0));
  nand2 gate666(.a(gate79inter0), .b(s_72), .O(gate79inter1));
  and2  gate667(.a(N186), .b(N230), .O(gate79inter2));
  inv1  gate668(.a(s_72), .O(gate79inter3));
  inv1  gate669(.a(s_73), .O(gate79inter4));
  nand2 gate670(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate671(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate672(.a(N230), .O(gate79inter7));
  inv1  gate673(.a(N186), .O(gate79inter8));
  nand2 gate674(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate675(.a(s_73), .b(gate79inter3), .O(gate79inter10));
  nor2  gate676(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate677(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate678(.a(gate79inter12), .b(gate79inter1), .O(N289));

  xor2  gate553(.a(N188), .b(N233), .O(gate80inter0));
  nand2 gate554(.a(gate80inter0), .b(s_56), .O(gate80inter1));
  and2  gate555(.a(N188), .b(N233), .O(gate80inter2));
  inv1  gate556(.a(s_56), .O(gate80inter3));
  inv1  gate557(.a(s_57), .O(gate80inter4));
  nand2 gate558(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate559(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate560(.a(N233), .O(gate80inter7));
  inv1  gate561(.a(N188), .O(gate80inter8));
  nand2 gate562(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate563(.a(s_57), .b(gate80inter3), .O(gate80inter10));
  nor2  gate564(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate565(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate566(.a(gate80inter12), .b(gate80inter1), .O(N290));
nand2 gate81( .a(N236), .b(N190), .O(N291) );
nand2 gate82( .a(N239), .b(N192), .O(N292) );
nand2 gate83( .a(N243), .b(N194), .O(N293) );
nand2 gate84( .a(N247), .b(N196), .O(N294) );
nand2 gate85( .a(N251), .b(N198), .O(N295) );
and9 gate86( .a(N260), .b(N264), .c(N267), .d(N270), .e(N273), .f(N276), .g(N279), .h(N282), .i(N285), .O(N296) );
inv1 gate87( .a(N263), .O(N300) );
inv1 gate88( .a(N288), .O(N301) );
inv1 gate89( .a(N289), .O(N302) );
inv1 gate90( .a(N290), .O(N303) );
inv1 gate91( .a(N291), .O(N304) );
inv1 gate92( .a(N292), .O(N305) );
inv1 gate93( .a(N293), .O(N306) );
inv1 gate94( .a(N294), .O(N307) );
inv1 gate95( .a(N295), .O(N308) );
inv1 gate96( .a(N296), .O(N309) );
inv1 gate97( .a(N296), .O(N319) );
inv1 gate98( .a(N296), .O(N329) );
xor2 gate99( .a(N309), .b(N260), .O(N330) );
xor2 gate100( .a(N309), .b(N264), .O(N331) );

  xor2  gate581(.a(N267), .b(N309), .O(gate101inter0));
  nand2 gate582(.a(gate101inter0), .b(s_60), .O(gate101inter1));
  and2  gate583(.a(N267), .b(N309), .O(gate101inter2));
  inv1  gate584(.a(s_60), .O(gate101inter3));
  inv1  gate585(.a(s_61), .O(gate101inter4));
  nand2 gate586(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate587(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate588(.a(N309), .O(gate101inter7));
  inv1  gate589(.a(N267), .O(gate101inter8));
  nand2 gate590(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate591(.a(s_61), .b(gate101inter3), .O(gate101inter10));
  nor2  gate592(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate593(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate594(.a(gate101inter12), .b(gate101inter1), .O(N332));
xor2 gate102( .a(N309), .b(N270), .O(N333) );
nand2 gate103( .a(N8), .b(N319), .O(N334) );
xor2 gate104( .a(N309), .b(N273), .O(N335) );

  xor2  gate749(.a(N21), .b(N319), .O(gate105inter0));
  nand2 gate750(.a(gate105inter0), .b(s_84), .O(gate105inter1));
  and2  gate751(.a(N21), .b(N319), .O(gate105inter2));
  inv1  gate752(.a(s_84), .O(gate105inter3));
  inv1  gate753(.a(s_85), .O(gate105inter4));
  nand2 gate754(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate755(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate756(.a(N319), .O(gate105inter7));
  inv1  gate757(.a(N21), .O(gate105inter8));
  nand2 gate758(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate759(.a(s_85), .b(gate105inter3), .O(gate105inter10));
  nor2  gate760(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate761(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate762(.a(gate105inter12), .b(gate105inter1), .O(N336));

  xor2  gate623(.a(N276), .b(N309), .O(gate106inter0));
  nand2 gate624(.a(gate106inter0), .b(s_66), .O(gate106inter1));
  and2  gate625(.a(N276), .b(N309), .O(gate106inter2));
  inv1  gate626(.a(s_66), .O(gate106inter3));
  inv1  gate627(.a(s_67), .O(gate106inter4));
  nand2 gate628(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate629(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate630(.a(N309), .O(gate106inter7));
  inv1  gate631(.a(N276), .O(gate106inter8));
  nand2 gate632(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate633(.a(s_67), .b(gate106inter3), .O(gate106inter10));
  nor2  gate634(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate635(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate636(.a(gate106inter12), .b(gate106inter1), .O(N337));
nand2 gate107( .a(N319), .b(N34), .O(N338) );
xor2 gate108( .a(N309), .b(N279), .O(N339) );
nand2 gate109( .a(N319), .b(N47), .O(N340) );

  xor2  gate245(.a(N282), .b(N309), .O(gate110inter0));
  nand2 gate246(.a(gate110inter0), .b(s_12), .O(gate110inter1));
  and2  gate247(.a(N282), .b(N309), .O(gate110inter2));
  inv1  gate248(.a(s_12), .O(gate110inter3));
  inv1  gate249(.a(s_13), .O(gate110inter4));
  nand2 gate250(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate251(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate252(.a(N309), .O(gate110inter7));
  inv1  gate253(.a(N282), .O(gate110inter8));
  nand2 gate254(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate255(.a(s_13), .b(gate110inter3), .O(gate110inter10));
  nor2  gate256(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate257(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate258(.a(gate110inter12), .b(gate110inter1), .O(N341));
nand2 gate111( .a(N319), .b(N60), .O(N342) );

  xor2  gate413(.a(N285), .b(N309), .O(gate112inter0));
  nand2 gate414(.a(gate112inter0), .b(s_36), .O(gate112inter1));
  and2  gate415(.a(N285), .b(N309), .O(gate112inter2));
  inv1  gate416(.a(s_36), .O(gate112inter3));
  inv1  gate417(.a(s_37), .O(gate112inter4));
  nand2 gate418(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate419(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate420(.a(N309), .O(gate112inter7));
  inv1  gate421(.a(N285), .O(gate112inter8));
  nand2 gate422(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate423(.a(s_37), .b(gate112inter3), .O(gate112inter10));
  nor2  gate424(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate425(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate426(.a(gate112inter12), .b(gate112inter1), .O(N343));
nand2 gate113( .a(N319), .b(N73), .O(N344) );
nand2 gate114( .a(N319), .b(N86), .O(N345) );

  xor2  gate217(.a(N99), .b(N319), .O(gate115inter0));
  nand2 gate218(.a(gate115inter0), .b(s_8), .O(gate115inter1));
  and2  gate219(.a(N99), .b(N319), .O(gate115inter2));
  inv1  gate220(.a(s_8), .O(gate115inter3));
  inv1  gate221(.a(s_9), .O(gate115inter4));
  nand2 gate222(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate223(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate224(.a(N319), .O(gate115inter7));
  inv1  gate225(.a(N99), .O(gate115inter8));
  nand2 gate226(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate227(.a(s_9), .b(gate115inter3), .O(gate115inter10));
  nor2  gate228(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate229(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate230(.a(gate115inter12), .b(gate115inter1), .O(N346));

  xor2  gate469(.a(N112), .b(N319), .O(gate116inter0));
  nand2 gate470(.a(gate116inter0), .b(s_44), .O(gate116inter1));
  and2  gate471(.a(N112), .b(N319), .O(gate116inter2));
  inv1  gate472(.a(s_44), .O(gate116inter3));
  inv1  gate473(.a(s_45), .O(gate116inter4));
  nand2 gate474(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate475(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate476(.a(N319), .O(gate116inter7));
  inv1  gate477(.a(N112), .O(gate116inter8));
  nand2 gate478(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate479(.a(s_45), .b(gate116inter3), .O(gate116inter10));
  nor2  gate480(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate481(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate482(.a(gate116inter12), .b(gate116inter1), .O(N347));

  xor2  gate777(.a(N300), .b(N330), .O(gate117inter0));
  nand2 gate778(.a(gate117inter0), .b(s_88), .O(gate117inter1));
  and2  gate779(.a(N300), .b(N330), .O(gate117inter2));
  inv1  gate780(.a(s_88), .O(gate117inter3));
  inv1  gate781(.a(s_89), .O(gate117inter4));
  nand2 gate782(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate783(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate784(.a(N330), .O(gate117inter7));
  inv1  gate785(.a(N300), .O(gate117inter8));
  nand2 gate786(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate787(.a(s_89), .b(gate117inter3), .O(gate117inter10));
  nor2  gate788(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate789(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate790(.a(gate117inter12), .b(gate117inter1), .O(N348));

  xor2  gate427(.a(N301), .b(N331), .O(gate118inter0));
  nand2 gate428(.a(gate118inter0), .b(s_38), .O(gate118inter1));
  and2  gate429(.a(N301), .b(N331), .O(gate118inter2));
  inv1  gate430(.a(s_38), .O(gate118inter3));
  inv1  gate431(.a(s_39), .O(gate118inter4));
  nand2 gate432(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate433(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate434(.a(N331), .O(gate118inter7));
  inv1  gate435(.a(N301), .O(gate118inter8));
  nand2 gate436(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate437(.a(s_39), .b(gate118inter3), .O(gate118inter10));
  nor2  gate438(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate439(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate440(.a(gate118inter12), .b(gate118inter1), .O(N349));
nand2 gate119( .a(N332), .b(N302), .O(N350) );
nand2 gate120( .a(N333), .b(N303), .O(N351) );
nand2 gate121( .a(N335), .b(N304), .O(N352) );
nand2 gate122( .a(N337), .b(N305), .O(N353) );

  xor2  gate483(.a(N306), .b(N339), .O(gate123inter0));
  nand2 gate484(.a(gate123inter0), .b(s_46), .O(gate123inter1));
  and2  gate485(.a(N306), .b(N339), .O(gate123inter2));
  inv1  gate486(.a(s_46), .O(gate123inter3));
  inv1  gate487(.a(s_47), .O(gate123inter4));
  nand2 gate488(.a(gate123inter4), .b(gate123inter3), .O(gate123inter5));
  nor2  gate489(.a(gate123inter5), .b(gate123inter2), .O(gate123inter6));
  inv1  gate490(.a(N339), .O(gate123inter7));
  inv1  gate491(.a(N306), .O(gate123inter8));
  nand2 gate492(.a(gate123inter8), .b(gate123inter7), .O(gate123inter9));
  nand2 gate493(.a(s_47), .b(gate123inter3), .O(gate123inter10));
  nor2  gate494(.a(gate123inter10), .b(gate123inter9), .O(gate123inter11));
  nor2  gate495(.a(gate123inter11), .b(gate123inter6), .O(gate123inter12));
  nand2 gate496(.a(gate123inter12), .b(gate123inter1), .O(N354));

  xor2  gate511(.a(N307), .b(N341), .O(gate124inter0));
  nand2 gate512(.a(gate124inter0), .b(s_50), .O(gate124inter1));
  and2  gate513(.a(N307), .b(N341), .O(gate124inter2));
  inv1  gate514(.a(s_50), .O(gate124inter3));
  inv1  gate515(.a(s_51), .O(gate124inter4));
  nand2 gate516(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate517(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate518(.a(N341), .O(gate124inter7));
  inv1  gate519(.a(N307), .O(gate124inter8));
  nand2 gate520(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate521(.a(s_51), .b(gate124inter3), .O(gate124inter10));
  nor2  gate522(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate523(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate524(.a(gate124inter12), .b(gate124inter1), .O(N355));
nand2 gate125( .a(N343), .b(N308), .O(N356) );
and9 gate126( .a(N348), .b(N349), .c(N350), .d(N351), .e(N352), .f(N353), .g(N354), .h(N355), .i(N356), .O(N357) );
inv1 gate127( .a(N357), .O(N360) );
inv1 gate128( .a(N357), .O(N370) );

  xor2  gate651(.a(N360), .b(N14), .O(gate129inter0));
  nand2 gate652(.a(gate129inter0), .b(s_70), .O(gate129inter1));
  and2  gate653(.a(N360), .b(N14), .O(gate129inter2));
  inv1  gate654(.a(s_70), .O(gate129inter3));
  inv1  gate655(.a(s_71), .O(gate129inter4));
  nand2 gate656(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate657(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate658(.a(N14), .O(gate129inter7));
  inv1  gate659(.a(N360), .O(gate129inter8));
  nand2 gate660(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate661(.a(s_71), .b(gate129inter3), .O(gate129inter10));
  nor2  gate662(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate663(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate664(.a(gate129inter12), .b(gate129inter1), .O(N371));

  xor2  gate595(.a(N27), .b(N360), .O(gate130inter0));
  nand2 gate596(.a(gate130inter0), .b(s_62), .O(gate130inter1));
  and2  gate597(.a(N27), .b(N360), .O(gate130inter2));
  inv1  gate598(.a(s_62), .O(gate130inter3));
  inv1  gate599(.a(s_63), .O(gate130inter4));
  nand2 gate600(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate601(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate602(.a(N360), .O(gate130inter7));
  inv1  gate603(.a(N27), .O(gate130inter8));
  nand2 gate604(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate605(.a(s_63), .b(gate130inter3), .O(gate130inter10));
  nor2  gate606(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate607(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate608(.a(gate130inter12), .b(gate130inter1), .O(N372));
nand2 gate131( .a(N360), .b(N40), .O(N373) );
nand2 gate132( .a(N360), .b(N53), .O(N374) );

  xor2  gate385(.a(N66), .b(N360), .O(gate133inter0));
  nand2 gate386(.a(gate133inter0), .b(s_32), .O(gate133inter1));
  and2  gate387(.a(N66), .b(N360), .O(gate133inter2));
  inv1  gate388(.a(s_32), .O(gate133inter3));
  inv1  gate389(.a(s_33), .O(gate133inter4));
  nand2 gate390(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate391(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate392(.a(N360), .O(gate133inter7));
  inv1  gate393(.a(N66), .O(gate133inter8));
  nand2 gate394(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate395(.a(s_33), .b(gate133inter3), .O(gate133inter10));
  nor2  gate396(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate397(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate398(.a(gate133inter12), .b(gate133inter1), .O(N375));
nand2 gate134( .a(N360), .b(N79), .O(N376) );

  xor2  gate329(.a(N92), .b(N360), .O(gate135inter0));
  nand2 gate330(.a(gate135inter0), .b(s_24), .O(gate135inter1));
  and2  gate331(.a(N92), .b(N360), .O(gate135inter2));
  inv1  gate332(.a(s_24), .O(gate135inter3));
  inv1  gate333(.a(s_25), .O(gate135inter4));
  nand2 gate334(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate335(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate336(.a(N360), .O(gate135inter7));
  inv1  gate337(.a(N92), .O(gate135inter8));
  nand2 gate338(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate339(.a(s_25), .b(gate135inter3), .O(gate135inter10));
  nor2  gate340(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate341(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate342(.a(gate135inter12), .b(gate135inter1), .O(N377));

  xor2  gate371(.a(N105), .b(N360), .O(gate136inter0));
  nand2 gate372(.a(gate136inter0), .b(s_30), .O(gate136inter1));
  and2  gate373(.a(N105), .b(N360), .O(gate136inter2));
  inv1  gate374(.a(s_30), .O(gate136inter3));
  inv1  gate375(.a(s_31), .O(gate136inter4));
  nand2 gate376(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate377(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate378(.a(N360), .O(gate136inter7));
  inv1  gate379(.a(N105), .O(gate136inter8));
  nand2 gate380(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate381(.a(s_31), .b(gate136inter3), .O(gate136inter10));
  nor2  gate382(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate383(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate384(.a(gate136inter12), .b(gate136inter1), .O(N378));
nand2 gate137( .a(N360), .b(N115), .O(N379) );
nand4 gate138( .a(N4), .b(N242), .c(N334), .d(N371), .O(N380) );
nand4 gate139( .a(N246), .b(N336), .c(N372), .d(N17), .O(N381) );
nand4 gate140( .a(N250), .b(N338), .c(N373), .d(N30), .O(N386) );
nand4 gate141( .a(N254), .b(N340), .c(N374), .d(N43), .O(N393) );
nand4 gate142( .a(N255), .b(N342), .c(N375), .d(N56), .O(N399) );
nand4 gate143( .a(N256), .b(N344), .c(N376), .d(N69), .O(N404) );
nand4 gate144( .a(N257), .b(N345), .c(N377), .d(N82), .O(N407) );
nand4 gate145( .a(N258), .b(N346), .c(N378), .d(N95), .O(N411) );
nand4 gate146( .a(N259), .b(N347), .c(N379), .d(N108), .O(N414) );
inv1 gate147( .a(N380), .O(N415) );
and8 gate148( .a(N381), .b(N386), .c(N393), .d(N399), .e(N404), .f(N407), .g(N411), .h(N414), .O(N416) );
inv1 gate149( .a(N393), .O(N417) );
inv1 gate150( .a(N404), .O(N418) );
inv1 gate151( .a(N407), .O(N419) );
inv1 gate152( .a(N411), .O(N420) );
nor2 gate153( .a(N415), .b(N416), .O(N421) );

  xor2  gate693(.a(N417), .b(N386), .O(gate154inter0));
  nand2 gate694(.a(gate154inter0), .b(s_76), .O(gate154inter1));
  and2  gate695(.a(N417), .b(N386), .O(gate154inter2));
  inv1  gate696(.a(s_76), .O(gate154inter3));
  inv1  gate697(.a(s_77), .O(gate154inter4));
  nand2 gate698(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate699(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate700(.a(N386), .O(gate154inter7));
  inv1  gate701(.a(N417), .O(gate154inter8));
  nand2 gate702(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate703(.a(s_77), .b(gate154inter3), .O(gate154inter10));
  nor2  gate704(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate705(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate706(.a(gate154inter12), .b(gate154inter1), .O(N422));
nand4 gate155( .a(N386), .b(N393), .c(N418), .d(N399), .O(N425) );
nand3 gate156( .a(N399), .b(N393), .c(N419), .O(N428) );
nand4 gate157( .a(N386), .b(N393), .c(N407), .d(N420), .O(N429) );
nand4 gate158( .a(N381), .b(N386), .c(N422), .d(N399), .O(N430) );
nand4 gate159( .a(N381), .b(N386), .c(N425), .d(N428), .O(N431) );
nand4 gate160( .a(N381), .b(N422), .c(N425), .d(N429), .O(N432) );

endmodule