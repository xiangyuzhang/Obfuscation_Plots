module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate631(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate632(.a(gate9inter0), .b(s_12), .O(gate9inter1));
  and2  gate633(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate634(.a(s_12), .O(gate9inter3));
  inv1  gate635(.a(s_13), .O(gate9inter4));
  nand2 gate636(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate637(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate638(.a(G1), .O(gate9inter7));
  inv1  gate639(.a(G2), .O(gate9inter8));
  nand2 gate640(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate641(.a(s_13), .b(gate9inter3), .O(gate9inter10));
  nor2  gate642(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate643(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate644(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate1275(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate1276(.a(gate12inter0), .b(s_104), .O(gate12inter1));
  and2  gate1277(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate1278(.a(s_104), .O(gate12inter3));
  inv1  gate1279(.a(s_105), .O(gate12inter4));
  nand2 gate1280(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate1281(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate1282(.a(G7), .O(gate12inter7));
  inv1  gate1283(.a(G8), .O(gate12inter8));
  nand2 gate1284(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate1285(.a(s_105), .b(gate12inter3), .O(gate12inter10));
  nor2  gate1286(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate1287(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate1288(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate855(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate856(.a(gate17inter0), .b(s_44), .O(gate17inter1));
  and2  gate857(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate858(.a(s_44), .O(gate17inter3));
  inv1  gate859(.a(s_45), .O(gate17inter4));
  nand2 gate860(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate861(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate862(.a(G17), .O(gate17inter7));
  inv1  gate863(.a(G18), .O(gate17inter8));
  nand2 gate864(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate865(.a(s_45), .b(gate17inter3), .O(gate17inter10));
  nor2  gate866(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate867(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate868(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate827(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate828(.a(gate19inter0), .b(s_40), .O(gate19inter1));
  and2  gate829(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate830(.a(s_40), .O(gate19inter3));
  inv1  gate831(.a(s_41), .O(gate19inter4));
  nand2 gate832(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate833(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate834(.a(G21), .O(gate19inter7));
  inv1  gate835(.a(G22), .O(gate19inter8));
  nand2 gate836(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate837(.a(s_41), .b(gate19inter3), .O(gate19inter10));
  nor2  gate838(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate839(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate840(.a(gate19inter12), .b(gate19inter1), .O(G296));

  xor2  gate645(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate646(.a(gate20inter0), .b(s_14), .O(gate20inter1));
  and2  gate647(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate648(.a(s_14), .O(gate20inter3));
  inv1  gate649(.a(s_15), .O(gate20inter4));
  nand2 gate650(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate651(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate652(.a(G23), .O(gate20inter7));
  inv1  gate653(.a(G24), .O(gate20inter8));
  nand2 gate654(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate655(.a(s_15), .b(gate20inter3), .O(gate20inter10));
  nor2  gate656(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate657(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate658(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate743(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate744(.a(gate29inter0), .b(s_28), .O(gate29inter1));
  and2  gate745(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate746(.a(s_28), .O(gate29inter3));
  inv1  gate747(.a(s_29), .O(gate29inter4));
  nand2 gate748(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate749(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate750(.a(G3), .O(gate29inter7));
  inv1  gate751(.a(G7), .O(gate29inter8));
  nand2 gate752(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate753(.a(s_29), .b(gate29inter3), .O(gate29inter10));
  nor2  gate754(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate755(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate756(.a(gate29inter12), .b(gate29inter1), .O(G326));

  xor2  gate799(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate800(.a(gate30inter0), .b(s_36), .O(gate30inter1));
  and2  gate801(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate802(.a(s_36), .O(gate30inter3));
  inv1  gate803(.a(s_37), .O(gate30inter4));
  nand2 gate804(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate805(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate806(.a(G11), .O(gate30inter7));
  inv1  gate807(.a(G15), .O(gate30inter8));
  nand2 gate808(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate809(.a(s_37), .b(gate30inter3), .O(gate30inter10));
  nor2  gate810(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate811(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate812(.a(gate30inter12), .b(gate30inter1), .O(G329));
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate1331(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate1332(.a(gate36inter0), .b(s_112), .O(gate36inter1));
  and2  gate1333(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate1334(.a(s_112), .O(gate36inter3));
  inv1  gate1335(.a(s_113), .O(gate36inter4));
  nand2 gate1336(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate1337(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate1338(.a(G26), .O(gate36inter7));
  inv1  gate1339(.a(G30), .O(gate36inter8));
  nand2 gate1340(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate1341(.a(s_113), .b(gate36inter3), .O(gate36inter10));
  nor2  gate1342(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate1343(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate1344(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate1415(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate1416(.a(gate41inter0), .b(s_124), .O(gate41inter1));
  and2  gate1417(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate1418(.a(s_124), .O(gate41inter3));
  inv1  gate1419(.a(s_125), .O(gate41inter4));
  nand2 gate1420(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate1421(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate1422(.a(G1), .O(gate41inter7));
  inv1  gate1423(.a(G266), .O(gate41inter8));
  nand2 gate1424(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate1425(.a(s_125), .b(gate41inter3), .O(gate41inter10));
  nor2  gate1426(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate1427(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate1428(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );

  xor2  gate1247(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate1248(.a(gate45inter0), .b(s_100), .O(gate45inter1));
  and2  gate1249(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate1250(.a(s_100), .O(gate45inter3));
  inv1  gate1251(.a(s_101), .O(gate45inter4));
  nand2 gate1252(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate1253(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate1254(.a(G5), .O(gate45inter7));
  inv1  gate1255(.a(G272), .O(gate45inter8));
  nand2 gate1256(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate1257(.a(s_101), .b(gate45inter3), .O(gate45inter10));
  nor2  gate1258(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate1259(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate1260(.a(gate45inter12), .b(gate45inter1), .O(G366));
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate659(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate660(.a(gate54inter0), .b(s_16), .O(gate54inter1));
  and2  gate661(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate662(.a(s_16), .O(gate54inter3));
  inv1  gate663(.a(s_17), .O(gate54inter4));
  nand2 gate664(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate665(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate666(.a(G14), .O(gate54inter7));
  inv1  gate667(.a(G284), .O(gate54inter8));
  nand2 gate668(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate669(.a(s_17), .b(gate54inter3), .O(gate54inter10));
  nor2  gate670(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate671(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate672(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );

  xor2  gate1177(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate1178(.a(gate56inter0), .b(s_90), .O(gate56inter1));
  and2  gate1179(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate1180(.a(s_90), .O(gate56inter3));
  inv1  gate1181(.a(s_91), .O(gate56inter4));
  nand2 gate1182(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate1183(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate1184(.a(G16), .O(gate56inter7));
  inv1  gate1185(.a(G287), .O(gate56inter8));
  nand2 gate1186(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate1187(.a(s_91), .b(gate56inter3), .O(gate56inter10));
  nor2  gate1188(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate1189(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate1190(.a(gate56inter12), .b(gate56inter1), .O(G377));

  xor2  gate1373(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate1374(.a(gate57inter0), .b(s_118), .O(gate57inter1));
  and2  gate1375(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate1376(.a(s_118), .O(gate57inter3));
  inv1  gate1377(.a(s_119), .O(gate57inter4));
  nand2 gate1378(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate1379(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate1380(.a(G17), .O(gate57inter7));
  inv1  gate1381(.a(G290), .O(gate57inter8));
  nand2 gate1382(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate1383(.a(s_119), .b(gate57inter3), .O(gate57inter10));
  nor2  gate1384(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate1385(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate1386(.a(gate57inter12), .b(gate57inter1), .O(G378));
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate1443(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate1444(.a(gate66inter0), .b(s_128), .O(gate66inter1));
  and2  gate1445(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate1446(.a(s_128), .O(gate66inter3));
  inv1  gate1447(.a(s_129), .O(gate66inter4));
  nand2 gate1448(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate1449(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate1450(.a(G26), .O(gate66inter7));
  inv1  gate1451(.a(G302), .O(gate66inter8));
  nand2 gate1452(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate1453(.a(s_129), .b(gate66inter3), .O(gate66inter10));
  nor2  gate1454(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate1455(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate1456(.a(gate66inter12), .b(gate66inter1), .O(G387));

  xor2  gate1359(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate1360(.a(gate67inter0), .b(s_116), .O(gate67inter1));
  and2  gate1361(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate1362(.a(s_116), .O(gate67inter3));
  inv1  gate1363(.a(s_117), .O(gate67inter4));
  nand2 gate1364(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate1365(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate1366(.a(G27), .O(gate67inter7));
  inv1  gate1367(.a(G305), .O(gate67inter8));
  nand2 gate1368(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate1369(.a(s_117), .b(gate67inter3), .O(gate67inter10));
  nor2  gate1370(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate1371(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate1372(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate729(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate730(.a(gate70inter0), .b(s_26), .O(gate70inter1));
  and2  gate731(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate732(.a(s_26), .O(gate70inter3));
  inv1  gate733(.a(s_27), .O(gate70inter4));
  nand2 gate734(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate735(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate736(.a(G30), .O(gate70inter7));
  inv1  gate737(.a(G308), .O(gate70inter8));
  nand2 gate738(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate739(.a(s_27), .b(gate70inter3), .O(gate70inter10));
  nor2  gate740(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate741(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate742(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );

  xor2  gate785(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate786(.a(gate84inter0), .b(s_34), .O(gate84inter1));
  and2  gate787(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate788(.a(s_34), .O(gate84inter3));
  inv1  gate789(.a(s_35), .O(gate84inter4));
  nand2 gate790(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate791(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate792(.a(G15), .O(gate84inter7));
  inv1  gate793(.a(G329), .O(gate84inter8));
  nand2 gate794(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate795(.a(s_35), .b(gate84inter3), .O(gate84inter10));
  nor2  gate796(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate797(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate798(.a(gate84inter12), .b(gate84inter1), .O(G405));
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );

  xor2  gate841(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate842(.a(gate89inter0), .b(s_42), .O(gate89inter1));
  and2  gate843(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate844(.a(s_42), .O(gate89inter3));
  inv1  gate845(.a(s_43), .O(gate89inter4));
  nand2 gate846(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate847(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate848(.a(G17), .O(gate89inter7));
  inv1  gate849(.a(G338), .O(gate89inter8));
  nand2 gate850(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate851(.a(s_43), .b(gate89inter3), .O(gate89inter10));
  nor2  gate852(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate853(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate854(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );

  xor2  gate925(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate926(.a(gate97inter0), .b(s_54), .O(gate97inter1));
  and2  gate927(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate928(.a(s_54), .O(gate97inter3));
  inv1  gate929(.a(s_55), .O(gate97inter4));
  nand2 gate930(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate931(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate932(.a(G19), .O(gate97inter7));
  inv1  gate933(.a(G350), .O(gate97inter8));
  nand2 gate934(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate935(.a(s_55), .b(gate97inter3), .O(gate97inter10));
  nor2  gate936(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate937(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate938(.a(gate97inter12), .b(gate97inter1), .O(G418));
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate1135(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate1136(.a(gate102inter0), .b(s_84), .O(gate102inter1));
  and2  gate1137(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate1138(.a(s_84), .O(gate102inter3));
  inv1  gate1139(.a(s_85), .O(gate102inter4));
  nand2 gate1140(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate1141(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate1142(.a(G24), .O(gate102inter7));
  inv1  gate1143(.a(G356), .O(gate102inter8));
  nand2 gate1144(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate1145(.a(s_85), .b(gate102inter3), .O(gate102inter10));
  nor2  gate1146(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate1147(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate1148(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate1457(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate1458(.a(gate104inter0), .b(s_130), .O(gate104inter1));
  and2  gate1459(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate1460(.a(s_130), .O(gate104inter3));
  inv1  gate1461(.a(s_131), .O(gate104inter4));
  nand2 gate1462(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate1463(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate1464(.a(G32), .O(gate104inter7));
  inv1  gate1465(.a(G359), .O(gate104inter8));
  nand2 gate1466(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate1467(.a(s_131), .b(gate104inter3), .O(gate104inter10));
  nor2  gate1468(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate1469(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate1470(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate1429(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate1430(.a(gate124inter0), .b(s_126), .O(gate124inter1));
  and2  gate1431(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate1432(.a(s_126), .O(gate124inter3));
  inv1  gate1433(.a(s_127), .O(gate124inter4));
  nand2 gate1434(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate1435(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate1436(.a(G400), .O(gate124inter7));
  inv1  gate1437(.a(G401), .O(gate124inter8));
  nand2 gate1438(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate1439(.a(s_127), .b(gate124inter3), .O(gate124inter10));
  nor2  gate1440(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate1441(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate1442(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate1205(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate1206(.a(gate135inter0), .b(s_94), .O(gate135inter1));
  and2  gate1207(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate1208(.a(s_94), .O(gate135inter3));
  inv1  gate1209(.a(s_95), .O(gate135inter4));
  nand2 gate1210(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate1211(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate1212(.a(G422), .O(gate135inter7));
  inv1  gate1213(.a(G423), .O(gate135inter8));
  nand2 gate1214(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate1215(.a(s_95), .b(gate135inter3), .O(gate135inter10));
  nor2  gate1216(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate1217(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate1218(.a(gate135inter12), .b(gate135inter1), .O(G516));

  xor2  gate911(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate912(.a(gate136inter0), .b(s_52), .O(gate136inter1));
  and2  gate913(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate914(.a(s_52), .O(gate136inter3));
  inv1  gate915(.a(s_53), .O(gate136inter4));
  nand2 gate916(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate917(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate918(.a(G424), .O(gate136inter7));
  inv1  gate919(.a(G425), .O(gate136inter8));
  nand2 gate920(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate921(.a(s_53), .b(gate136inter3), .O(gate136inter10));
  nor2  gate922(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate923(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate924(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate1121(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate1122(.a(gate154inter0), .b(s_82), .O(gate154inter1));
  and2  gate1123(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate1124(.a(s_82), .O(gate154inter3));
  inv1  gate1125(.a(s_83), .O(gate154inter4));
  nand2 gate1126(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate1127(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate1128(.a(G429), .O(gate154inter7));
  inv1  gate1129(.a(G522), .O(gate154inter8));
  nand2 gate1130(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate1131(.a(s_83), .b(gate154inter3), .O(gate154inter10));
  nor2  gate1132(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate1133(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate1134(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate939(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate940(.a(gate157inter0), .b(s_56), .O(gate157inter1));
  and2  gate941(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate942(.a(s_56), .O(gate157inter3));
  inv1  gate943(.a(s_57), .O(gate157inter4));
  nand2 gate944(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate945(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate946(.a(G438), .O(gate157inter7));
  inv1  gate947(.a(G528), .O(gate157inter8));
  nand2 gate948(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate949(.a(s_57), .b(gate157inter3), .O(gate157inter10));
  nor2  gate950(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate951(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate952(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate1107(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate1108(.a(gate159inter0), .b(s_80), .O(gate159inter1));
  and2  gate1109(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate1110(.a(s_80), .O(gate159inter3));
  inv1  gate1111(.a(s_81), .O(gate159inter4));
  nand2 gate1112(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate1113(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate1114(.a(G444), .O(gate159inter7));
  inv1  gate1115(.a(G531), .O(gate159inter8));
  nand2 gate1116(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate1117(.a(s_81), .b(gate159inter3), .O(gate159inter10));
  nor2  gate1118(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate1119(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate1120(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate1093(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate1094(.a(gate162inter0), .b(s_78), .O(gate162inter1));
  and2  gate1095(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate1096(.a(s_78), .O(gate162inter3));
  inv1  gate1097(.a(s_79), .O(gate162inter4));
  nand2 gate1098(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate1099(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate1100(.a(G453), .O(gate162inter7));
  inv1  gate1101(.a(G534), .O(gate162inter8));
  nand2 gate1102(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate1103(.a(s_79), .b(gate162inter3), .O(gate162inter10));
  nor2  gate1104(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate1105(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate1106(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate1079(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate1080(.a(gate164inter0), .b(s_76), .O(gate164inter1));
  and2  gate1081(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate1082(.a(s_76), .O(gate164inter3));
  inv1  gate1083(.a(s_77), .O(gate164inter4));
  nand2 gate1084(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate1085(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate1086(.a(G459), .O(gate164inter7));
  inv1  gate1087(.a(G537), .O(gate164inter8));
  nand2 gate1088(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate1089(.a(s_77), .b(gate164inter3), .O(gate164inter10));
  nor2  gate1090(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate1091(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate1092(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );

  xor2  gate561(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate562(.a(gate166inter0), .b(s_2), .O(gate166inter1));
  and2  gate563(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate564(.a(s_2), .O(gate166inter3));
  inv1  gate565(.a(s_3), .O(gate166inter4));
  nand2 gate566(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate567(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate568(.a(G465), .O(gate166inter7));
  inv1  gate569(.a(G540), .O(gate166inter8));
  nand2 gate570(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate571(.a(s_3), .b(gate166inter3), .O(gate166inter10));
  nor2  gate572(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate573(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate574(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate715(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate716(.a(gate183inter0), .b(s_24), .O(gate183inter1));
  and2  gate717(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate718(.a(s_24), .O(gate183inter3));
  inv1  gate719(.a(s_25), .O(gate183inter4));
  nand2 gate720(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate721(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate722(.a(G516), .O(gate183inter7));
  inv1  gate723(.a(G567), .O(gate183inter8));
  nand2 gate724(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate725(.a(s_25), .b(gate183inter3), .O(gate183inter10));
  nor2  gate726(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate727(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate728(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate1345(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate1346(.a(gate198inter0), .b(s_114), .O(gate198inter1));
  and2  gate1347(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate1348(.a(s_114), .O(gate198inter3));
  inv1  gate1349(.a(s_115), .O(gate198inter4));
  nand2 gate1350(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate1351(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate1352(.a(G596), .O(gate198inter7));
  inv1  gate1353(.a(G597), .O(gate198inter8));
  nand2 gate1354(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate1355(.a(s_115), .b(gate198inter3), .O(gate198inter10));
  nor2  gate1356(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate1357(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate1358(.a(gate198inter12), .b(gate198inter1), .O(G657));
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate673(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate674(.a(gate200inter0), .b(s_18), .O(gate200inter1));
  and2  gate675(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate676(.a(s_18), .O(gate200inter3));
  inv1  gate677(.a(s_19), .O(gate200inter4));
  nand2 gate678(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate679(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate680(.a(G600), .O(gate200inter7));
  inv1  gate681(.a(G601), .O(gate200inter8));
  nand2 gate682(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate683(.a(s_19), .b(gate200inter3), .O(gate200inter10));
  nor2  gate684(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate685(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate686(.a(gate200inter12), .b(gate200inter1), .O(G663));
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate981(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate982(.a(gate203inter0), .b(s_62), .O(gate203inter1));
  and2  gate983(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate984(.a(s_62), .O(gate203inter3));
  inv1  gate985(.a(s_63), .O(gate203inter4));
  nand2 gate986(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate987(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate988(.a(G602), .O(gate203inter7));
  inv1  gate989(.a(G612), .O(gate203inter8));
  nand2 gate990(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate991(.a(s_63), .b(gate203inter3), .O(gate203inter10));
  nor2  gate992(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate993(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate994(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );

  xor2  gate1303(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate1304(.a(gate225inter0), .b(s_108), .O(gate225inter1));
  and2  gate1305(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate1306(.a(s_108), .O(gate225inter3));
  inv1  gate1307(.a(s_109), .O(gate225inter4));
  nand2 gate1308(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate1309(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate1310(.a(G690), .O(gate225inter7));
  inv1  gate1311(.a(G691), .O(gate225inter8));
  nand2 gate1312(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate1313(.a(s_109), .b(gate225inter3), .O(gate225inter10));
  nor2  gate1314(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate1315(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate1316(.a(gate225inter12), .b(gate225inter1), .O(G706));
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );

  xor2  gate967(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate968(.a(gate230inter0), .b(s_60), .O(gate230inter1));
  and2  gate969(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate970(.a(s_60), .O(gate230inter3));
  inv1  gate971(.a(s_61), .O(gate230inter4));
  nand2 gate972(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate973(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate974(.a(G700), .O(gate230inter7));
  inv1  gate975(.a(G701), .O(gate230inter8));
  nand2 gate976(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate977(.a(s_61), .b(gate230inter3), .O(gate230inter10));
  nor2  gate978(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate979(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate980(.a(gate230inter12), .b(gate230inter1), .O(G721));
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );

  xor2  gate1163(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate1164(.a(gate244inter0), .b(s_88), .O(gate244inter1));
  and2  gate1165(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate1166(.a(s_88), .O(gate244inter3));
  inv1  gate1167(.a(s_89), .O(gate244inter4));
  nand2 gate1168(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate1169(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate1170(.a(G721), .O(gate244inter7));
  inv1  gate1171(.a(G733), .O(gate244inter8));
  nand2 gate1172(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate1173(.a(s_89), .b(gate244inter3), .O(gate244inter10));
  nor2  gate1174(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate1175(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate1176(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate1051(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate1052(.a(gate248inter0), .b(s_72), .O(gate248inter1));
  and2  gate1053(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate1054(.a(s_72), .O(gate248inter3));
  inv1  gate1055(.a(s_73), .O(gate248inter4));
  nand2 gate1056(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate1057(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate1058(.a(G727), .O(gate248inter7));
  inv1  gate1059(.a(G739), .O(gate248inter8));
  nand2 gate1060(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate1061(.a(s_73), .b(gate248inter3), .O(gate248inter10));
  nor2  gate1062(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate1063(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate1064(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );

  xor2  gate1289(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate1290(.a(gate250inter0), .b(s_106), .O(gate250inter1));
  and2  gate1291(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate1292(.a(s_106), .O(gate250inter3));
  inv1  gate1293(.a(s_107), .O(gate250inter4));
  nand2 gate1294(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate1295(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate1296(.a(G706), .O(gate250inter7));
  inv1  gate1297(.a(G742), .O(gate250inter8));
  nand2 gate1298(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate1299(.a(s_107), .b(gate250inter3), .O(gate250inter10));
  nor2  gate1300(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate1301(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate1302(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate575(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate576(.a(gate263inter0), .b(s_4), .O(gate263inter1));
  and2  gate577(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate578(.a(s_4), .O(gate263inter3));
  inv1  gate579(.a(s_5), .O(gate263inter4));
  nand2 gate580(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate581(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate582(.a(G766), .O(gate263inter7));
  inv1  gate583(.a(G767), .O(gate263inter8));
  nand2 gate584(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate585(.a(s_5), .b(gate263inter3), .O(gate263inter10));
  nor2  gate586(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate587(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate588(.a(gate263inter12), .b(gate263inter1), .O(G788));

  xor2  gate1009(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate1010(.a(gate264inter0), .b(s_66), .O(gate264inter1));
  and2  gate1011(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate1012(.a(s_66), .O(gate264inter3));
  inv1  gate1013(.a(s_67), .O(gate264inter4));
  nand2 gate1014(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate1015(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate1016(.a(G768), .O(gate264inter7));
  inv1  gate1017(.a(G769), .O(gate264inter8));
  nand2 gate1018(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate1019(.a(s_67), .b(gate264inter3), .O(gate264inter10));
  nor2  gate1020(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate1021(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate1022(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate897(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate898(.a(gate268inter0), .b(s_50), .O(gate268inter1));
  and2  gate899(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate900(.a(s_50), .O(gate268inter3));
  inv1  gate901(.a(s_51), .O(gate268inter4));
  nand2 gate902(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate903(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate904(.a(G651), .O(gate268inter7));
  inv1  gate905(.a(G779), .O(gate268inter8));
  nand2 gate906(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate907(.a(s_51), .b(gate268inter3), .O(gate268inter10));
  nor2  gate908(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate909(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate910(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate1261(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate1262(.a(gate272inter0), .b(s_102), .O(gate272inter1));
  and2  gate1263(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate1264(.a(s_102), .O(gate272inter3));
  inv1  gate1265(.a(s_103), .O(gate272inter4));
  nand2 gate1266(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate1267(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate1268(.a(G663), .O(gate272inter7));
  inv1  gate1269(.a(G791), .O(gate272inter8));
  nand2 gate1270(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate1271(.a(s_103), .b(gate272inter3), .O(gate272inter10));
  nor2  gate1272(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate1273(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate1274(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate1065(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate1066(.a(gate280inter0), .b(s_74), .O(gate280inter1));
  and2  gate1067(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate1068(.a(s_74), .O(gate280inter3));
  inv1  gate1069(.a(s_75), .O(gate280inter4));
  nand2 gate1070(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate1071(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate1072(.a(G779), .O(gate280inter7));
  inv1  gate1073(.a(G803), .O(gate280inter8));
  nand2 gate1074(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate1075(.a(s_75), .b(gate280inter3), .O(gate280inter10));
  nor2  gate1076(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate1077(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate1078(.a(gate280inter12), .b(gate280inter1), .O(G825));
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate1191(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate1192(.a(gate287inter0), .b(s_92), .O(gate287inter1));
  and2  gate1193(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate1194(.a(s_92), .O(gate287inter3));
  inv1  gate1195(.a(s_93), .O(gate287inter4));
  nand2 gate1196(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate1197(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate1198(.a(G663), .O(gate287inter7));
  inv1  gate1199(.a(G815), .O(gate287inter8));
  nand2 gate1200(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate1201(.a(s_93), .b(gate287inter3), .O(gate287inter10));
  nor2  gate1202(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate1203(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate1204(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate617(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate618(.a(gate387inter0), .b(s_10), .O(gate387inter1));
  and2  gate619(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate620(.a(s_10), .O(gate387inter3));
  inv1  gate621(.a(s_11), .O(gate387inter4));
  nand2 gate622(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate623(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate624(.a(G1), .O(gate387inter7));
  inv1  gate625(.a(G1036), .O(gate387inter8));
  nand2 gate626(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate627(.a(s_11), .b(gate387inter3), .O(gate387inter10));
  nor2  gate628(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate629(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate630(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate995(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate996(.a(gate394inter0), .b(s_64), .O(gate394inter1));
  and2  gate997(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate998(.a(s_64), .O(gate394inter3));
  inv1  gate999(.a(s_65), .O(gate394inter4));
  nand2 gate1000(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate1001(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate1002(.a(G8), .O(gate394inter7));
  inv1  gate1003(.a(G1057), .O(gate394inter8));
  nand2 gate1004(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate1005(.a(s_65), .b(gate394inter3), .O(gate394inter10));
  nor2  gate1006(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate1007(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate1008(.a(gate394inter12), .b(gate394inter1), .O(G1153));

  xor2  gate1149(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate1150(.a(gate395inter0), .b(s_86), .O(gate395inter1));
  and2  gate1151(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate1152(.a(s_86), .O(gate395inter3));
  inv1  gate1153(.a(s_87), .O(gate395inter4));
  nand2 gate1154(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate1155(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate1156(.a(G9), .O(gate395inter7));
  inv1  gate1157(.a(G1060), .O(gate395inter8));
  nand2 gate1158(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate1159(.a(s_87), .b(gate395inter3), .O(gate395inter10));
  nor2  gate1160(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate1161(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate1162(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );

  xor2  gate757(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate758(.a(gate401inter0), .b(s_30), .O(gate401inter1));
  and2  gate759(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate760(.a(s_30), .O(gate401inter3));
  inv1  gate761(.a(s_31), .O(gate401inter4));
  nand2 gate762(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate763(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate764(.a(G15), .O(gate401inter7));
  inv1  gate765(.a(G1078), .O(gate401inter8));
  nand2 gate766(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate767(.a(s_31), .b(gate401inter3), .O(gate401inter10));
  nor2  gate768(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate769(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate770(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate1233(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate1234(.a(gate403inter0), .b(s_98), .O(gate403inter1));
  and2  gate1235(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate1236(.a(s_98), .O(gate403inter3));
  inv1  gate1237(.a(s_99), .O(gate403inter4));
  nand2 gate1238(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate1239(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate1240(.a(G17), .O(gate403inter7));
  inv1  gate1241(.a(G1084), .O(gate403inter8));
  nand2 gate1242(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate1243(.a(s_99), .b(gate403inter3), .O(gate403inter10));
  nor2  gate1244(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate1245(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate1246(.a(gate403inter12), .b(gate403inter1), .O(G1180));
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );

  xor2  gate1401(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate1402(.a(gate405inter0), .b(s_122), .O(gate405inter1));
  and2  gate1403(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate1404(.a(s_122), .O(gate405inter3));
  inv1  gate1405(.a(s_123), .O(gate405inter4));
  nand2 gate1406(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate1407(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate1408(.a(G19), .O(gate405inter7));
  inv1  gate1409(.a(G1090), .O(gate405inter8));
  nand2 gate1410(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate1411(.a(s_123), .b(gate405inter3), .O(gate405inter10));
  nor2  gate1412(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate1413(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate1414(.a(gate405inter12), .b(gate405inter1), .O(G1186));
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate701(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate702(.a(gate407inter0), .b(s_22), .O(gate407inter1));
  and2  gate703(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate704(.a(s_22), .O(gate407inter3));
  inv1  gate705(.a(s_23), .O(gate407inter4));
  nand2 gate706(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate707(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate708(.a(G21), .O(gate407inter7));
  inv1  gate709(.a(G1096), .O(gate407inter8));
  nand2 gate710(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate711(.a(s_23), .b(gate407inter3), .O(gate407inter10));
  nor2  gate712(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate713(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate714(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );

  xor2  gate1037(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate1038(.a(gate409inter0), .b(s_70), .O(gate409inter1));
  and2  gate1039(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate1040(.a(s_70), .O(gate409inter3));
  inv1  gate1041(.a(s_71), .O(gate409inter4));
  nand2 gate1042(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate1043(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate1044(.a(G23), .O(gate409inter7));
  inv1  gate1045(.a(G1102), .O(gate409inter8));
  nand2 gate1046(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate1047(.a(s_71), .b(gate409inter3), .O(gate409inter10));
  nor2  gate1048(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate1049(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate1050(.a(gate409inter12), .b(gate409inter1), .O(G1198));
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );

  xor2  gate813(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate814(.a(gate412inter0), .b(s_38), .O(gate412inter1));
  and2  gate815(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate816(.a(s_38), .O(gate412inter3));
  inv1  gate817(.a(s_39), .O(gate412inter4));
  nand2 gate818(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate819(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate820(.a(G26), .O(gate412inter7));
  inv1  gate821(.a(G1111), .O(gate412inter8));
  nand2 gate822(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate823(.a(s_39), .b(gate412inter3), .O(gate412inter10));
  nor2  gate824(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate825(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate826(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );

  xor2  gate1023(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate1024(.a(gate416inter0), .b(s_68), .O(gate416inter1));
  and2  gate1025(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate1026(.a(s_68), .O(gate416inter3));
  inv1  gate1027(.a(s_69), .O(gate416inter4));
  nand2 gate1028(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate1029(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate1030(.a(G30), .O(gate416inter7));
  inv1  gate1031(.a(G1123), .O(gate416inter8));
  nand2 gate1032(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate1033(.a(s_69), .b(gate416inter3), .O(gate416inter10));
  nor2  gate1034(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate1035(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate1036(.a(gate416inter12), .b(gate416inter1), .O(G1219));

  xor2  gate953(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate954(.a(gate417inter0), .b(s_58), .O(gate417inter1));
  and2  gate955(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate956(.a(s_58), .O(gate417inter3));
  inv1  gate957(.a(s_59), .O(gate417inter4));
  nand2 gate958(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate959(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate960(.a(G31), .O(gate417inter7));
  inv1  gate961(.a(G1126), .O(gate417inter8));
  nand2 gate962(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate963(.a(s_59), .b(gate417inter3), .O(gate417inter10));
  nor2  gate964(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate965(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate966(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate771(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate772(.a(gate419inter0), .b(s_32), .O(gate419inter1));
  and2  gate773(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate774(.a(s_32), .O(gate419inter3));
  inv1  gate775(.a(s_33), .O(gate419inter4));
  nand2 gate776(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate777(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate778(.a(G1), .O(gate419inter7));
  inv1  gate779(.a(G1132), .O(gate419inter8));
  nand2 gate780(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate781(.a(s_33), .b(gate419inter3), .O(gate419inter10));
  nor2  gate782(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate783(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate784(.a(gate419inter12), .b(gate419inter1), .O(G1228));
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate603(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate604(.a(gate431inter0), .b(s_8), .O(gate431inter1));
  and2  gate605(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate606(.a(s_8), .O(gate431inter3));
  inv1  gate607(.a(s_9), .O(gate431inter4));
  nand2 gate608(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate609(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate610(.a(G7), .O(gate431inter7));
  inv1  gate611(.a(G1150), .O(gate431inter8));
  nand2 gate612(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate613(.a(s_9), .b(gate431inter3), .O(gate431inter10));
  nor2  gate614(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate615(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate616(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate883(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate884(.a(gate435inter0), .b(s_48), .O(gate435inter1));
  and2  gate885(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate886(.a(s_48), .O(gate435inter3));
  inv1  gate887(.a(s_49), .O(gate435inter4));
  nand2 gate888(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate889(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate890(.a(G9), .O(gate435inter7));
  inv1  gate891(.a(G1156), .O(gate435inter8));
  nand2 gate892(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate893(.a(s_49), .b(gate435inter3), .O(gate435inter10));
  nor2  gate894(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate895(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate896(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate1317(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate1318(.a(gate441inter0), .b(s_110), .O(gate441inter1));
  and2  gate1319(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate1320(.a(s_110), .O(gate441inter3));
  inv1  gate1321(.a(s_111), .O(gate441inter4));
  nand2 gate1322(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate1323(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate1324(.a(G12), .O(gate441inter7));
  inv1  gate1325(.a(G1165), .O(gate441inter8));
  nand2 gate1326(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate1327(.a(s_111), .b(gate441inter3), .O(gate441inter10));
  nor2  gate1328(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate1329(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate1330(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );

  xor2  gate589(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate590(.a(gate449inter0), .b(s_6), .O(gate449inter1));
  and2  gate591(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate592(.a(s_6), .O(gate449inter3));
  inv1  gate593(.a(s_7), .O(gate449inter4));
  nand2 gate594(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate595(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate596(.a(G16), .O(gate449inter7));
  inv1  gate597(.a(G1177), .O(gate449inter8));
  nand2 gate598(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate599(.a(s_7), .b(gate449inter3), .O(gate449inter10));
  nor2  gate600(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate601(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate602(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate687(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate688(.a(gate453inter0), .b(s_20), .O(gate453inter1));
  and2  gate689(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate690(.a(s_20), .O(gate453inter3));
  inv1  gate691(.a(s_21), .O(gate453inter4));
  nand2 gate692(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate693(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate694(.a(G18), .O(gate453inter7));
  inv1  gate695(.a(G1183), .O(gate453inter8));
  nand2 gate696(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate697(.a(s_21), .b(gate453inter3), .O(gate453inter10));
  nor2  gate698(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate699(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate700(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate1387(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate1388(.a(gate459inter0), .b(s_120), .O(gate459inter1));
  and2  gate1389(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate1390(.a(s_120), .O(gate459inter3));
  inv1  gate1391(.a(s_121), .O(gate459inter4));
  nand2 gate1392(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate1393(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate1394(.a(G21), .O(gate459inter7));
  inv1  gate1395(.a(G1192), .O(gate459inter8));
  nand2 gate1396(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate1397(.a(s_121), .b(gate459inter3), .O(gate459inter10));
  nor2  gate1398(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate1399(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate1400(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate869(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate870(.a(gate492inter0), .b(s_46), .O(gate492inter1));
  and2  gate871(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate872(.a(s_46), .O(gate492inter3));
  inv1  gate873(.a(s_47), .O(gate492inter4));
  nand2 gate874(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate875(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate876(.a(G1246), .O(gate492inter7));
  inv1  gate877(.a(G1247), .O(gate492inter8));
  nand2 gate878(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate879(.a(s_47), .b(gate492inter3), .O(gate492inter10));
  nor2  gate880(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate881(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate882(.a(gate492inter12), .b(gate492inter1), .O(G1301));
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate1219(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1220(.a(gate494inter0), .b(s_96), .O(gate494inter1));
  and2  gate1221(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1222(.a(s_96), .O(gate494inter3));
  inv1  gate1223(.a(s_97), .O(gate494inter4));
  nand2 gate1224(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1225(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1226(.a(G1250), .O(gate494inter7));
  inv1  gate1227(.a(G1251), .O(gate494inter8));
  nand2 gate1228(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1229(.a(s_97), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1230(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1231(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1232(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate547(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate548(.a(gate500inter0), .b(s_0), .O(gate500inter1));
  and2  gate549(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate550(.a(s_0), .O(gate500inter3));
  inv1  gate551(.a(s_1), .O(gate500inter4));
  nand2 gate552(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate553(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate554(.a(G1262), .O(gate500inter7));
  inv1  gate555(.a(G1263), .O(gate500inter8));
  nand2 gate556(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate557(.a(s_1), .b(gate500inter3), .O(gate500inter10));
  nor2  gate558(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate559(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate560(.a(gate500inter12), .b(gate500inter1), .O(G1309));
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule