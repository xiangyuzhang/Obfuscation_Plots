module c432 (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
             N430,N431,N432);
input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
      N99,N102,N105,N108,N112,N115;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61;
output N223,N329,N370,N421,N430,N431,N432;
wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12;


inv1 gate1( .a(N1), .O(N118) );
inv1 gate2( .a(N4), .O(N119) );
inv1 gate3( .a(N11), .O(N122) );
inv1 gate4( .a(N17), .O(N123) );
inv1 gate5( .a(N24), .O(N126) );
inv1 gate6( .a(N30), .O(N127) );
inv1 gate7( .a(N37), .O(N130) );
inv1 gate8( .a(N43), .O(N131) );
inv1 gate9( .a(N50), .O(N134) );
inv1 gate10( .a(N56), .O(N135) );
inv1 gate11( .a(N63), .O(N138) );
inv1 gate12( .a(N69), .O(N139) );
inv1 gate13( .a(N76), .O(N142) );
inv1 gate14( .a(N82), .O(N143) );
inv1 gate15( .a(N89), .O(N146) );
inv1 gate16( .a(N95), .O(N147) );
inv1 gate17( .a(N102), .O(N150) );
inv1 gate18( .a(N108), .O(N151) );

  xor2  gate511(.a(N4), .b(N118), .O(gate19inter0));
  nand2 gate512(.a(gate19inter0), .b(s_50), .O(gate19inter1));
  and2  gate513(.a(N4), .b(N118), .O(gate19inter2));
  inv1  gate514(.a(s_50), .O(gate19inter3));
  inv1  gate515(.a(s_51), .O(gate19inter4));
  nand2 gate516(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate517(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate518(.a(N118), .O(gate19inter7));
  inv1  gate519(.a(N4), .O(gate19inter8));
  nand2 gate520(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate521(.a(s_51), .b(gate19inter3), .O(gate19inter10));
  nor2  gate522(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate523(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate524(.a(gate19inter12), .b(gate19inter1), .O(N154));

  xor2  gate525(.a(N119), .b(N8), .O(gate20inter0));
  nand2 gate526(.a(gate20inter0), .b(s_52), .O(gate20inter1));
  and2  gate527(.a(N119), .b(N8), .O(gate20inter2));
  inv1  gate528(.a(s_52), .O(gate20inter3));
  inv1  gate529(.a(s_53), .O(gate20inter4));
  nand2 gate530(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate531(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate532(.a(N8), .O(gate20inter7));
  inv1  gate533(.a(N119), .O(gate20inter8));
  nand2 gate534(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate535(.a(s_53), .b(gate20inter3), .O(gate20inter10));
  nor2  gate536(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate537(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate538(.a(gate20inter12), .b(gate20inter1), .O(N157));
nor2 gate21( .a(N14), .b(N119), .O(N158) );
nand2 gate22( .a(N122), .b(N17), .O(N159) );

  xor2  gate231(.a(N30), .b(N126), .O(gate23inter0));
  nand2 gate232(.a(gate23inter0), .b(s_10), .O(gate23inter1));
  and2  gate233(.a(N30), .b(N126), .O(gate23inter2));
  inv1  gate234(.a(s_10), .O(gate23inter3));
  inv1  gate235(.a(s_11), .O(gate23inter4));
  nand2 gate236(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate237(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate238(.a(N126), .O(gate23inter7));
  inv1  gate239(.a(N30), .O(gate23inter8));
  nand2 gate240(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate241(.a(s_11), .b(gate23inter3), .O(gate23inter10));
  nor2  gate242(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate243(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate244(.a(gate23inter12), .b(gate23inter1), .O(N162));
nand2 gate24( .a(N130), .b(N43), .O(N165) );
nand2 gate25( .a(N134), .b(N56), .O(N168) );
nand2 gate26( .a(N138), .b(N69), .O(N171) );
nand2 gate27( .a(N142), .b(N82), .O(N174) );
nand2 gate28( .a(N146), .b(N95), .O(N177) );

  xor2  gate441(.a(N108), .b(N150), .O(gate29inter0));
  nand2 gate442(.a(gate29inter0), .b(s_40), .O(gate29inter1));
  and2  gate443(.a(N108), .b(N150), .O(gate29inter2));
  inv1  gate444(.a(s_40), .O(gate29inter3));
  inv1  gate445(.a(s_41), .O(gate29inter4));
  nand2 gate446(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate447(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate448(.a(N150), .O(gate29inter7));
  inv1  gate449(.a(N108), .O(gate29inter8));
  nand2 gate450(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate451(.a(s_41), .b(gate29inter3), .O(gate29inter10));
  nor2  gate452(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate453(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate454(.a(gate29inter12), .b(gate29inter1), .O(N180));

  xor2  gate581(.a(N123), .b(N21), .O(gate30inter0));
  nand2 gate582(.a(gate30inter0), .b(s_60), .O(gate30inter1));
  and2  gate583(.a(N123), .b(N21), .O(gate30inter2));
  inv1  gate584(.a(s_60), .O(gate30inter3));
  inv1  gate585(.a(s_61), .O(gate30inter4));
  nand2 gate586(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate587(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate588(.a(N21), .O(gate30inter7));
  inv1  gate589(.a(N123), .O(gate30inter8));
  nand2 gate590(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate591(.a(s_61), .b(gate30inter3), .O(gate30inter10));
  nor2  gate592(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate593(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate594(.a(gate30inter12), .b(gate30inter1), .O(N183));
nor2 gate31( .a(N27), .b(N123), .O(N184) );

  xor2  gate483(.a(N127), .b(N34), .O(gate32inter0));
  nand2 gate484(.a(gate32inter0), .b(s_46), .O(gate32inter1));
  and2  gate485(.a(N127), .b(N34), .O(gate32inter2));
  inv1  gate486(.a(s_46), .O(gate32inter3));
  inv1  gate487(.a(s_47), .O(gate32inter4));
  nand2 gate488(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate489(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate490(.a(N34), .O(gate32inter7));
  inv1  gate491(.a(N127), .O(gate32inter8));
  nand2 gate492(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate493(.a(s_47), .b(gate32inter3), .O(gate32inter10));
  nor2  gate494(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate495(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate496(.a(gate32inter12), .b(gate32inter1), .O(N185));
nor2 gate33( .a(N40), .b(N127), .O(N186) );

  xor2  gate385(.a(N131), .b(N47), .O(gate34inter0));
  nand2 gate386(.a(gate34inter0), .b(s_32), .O(gate34inter1));
  and2  gate387(.a(N131), .b(N47), .O(gate34inter2));
  inv1  gate388(.a(s_32), .O(gate34inter3));
  inv1  gate389(.a(s_33), .O(gate34inter4));
  nand2 gate390(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate391(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate392(.a(N47), .O(gate34inter7));
  inv1  gate393(.a(N131), .O(gate34inter8));
  nand2 gate394(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate395(.a(s_33), .b(gate34inter3), .O(gate34inter10));
  nor2  gate396(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate397(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate398(.a(gate34inter12), .b(gate34inter1), .O(N187));
nor2 gate35( .a(N53), .b(N131), .O(N188) );
nor2 gate36( .a(N60), .b(N135), .O(N189) );

  xor2  gate217(.a(N135), .b(N66), .O(gate37inter0));
  nand2 gate218(.a(gate37inter0), .b(s_8), .O(gate37inter1));
  and2  gate219(.a(N135), .b(N66), .O(gate37inter2));
  inv1  gate220(.a(s_8), .O(gate37inter3));
  inv1  gate221(.a(s_9), .O(gate37inter4));
  nand2 gate222(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate223(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate224(.a(N66), .O(gate37inter7));
  inv1  gate225(.a(N135), .O(gate37inter8));
  nand2 gate226(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate227(.a(s_9), .b(gate37inter3), .O(gate37inter10));
  nor2  gate228(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate229(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate230(.a(gate37inter12), .b(gate37inter1), .O(N190));
nor2 gate38( .a(N73), .b(N139), .O(N191) );
nor2 gate39( .a(N79), .b(N139), .O(N192) );
nor2 gate40( .a(N86), .b(N143), .O(N193) );
nor2 gate41( .a(N92), .b(N143), .O(N194) );

  xor2  gate301(.a(N147), .b(N99), .O(gate42inter0));
  nand2 gate302(.a(gate42inter0), .b(s_20), .O(gate42inter1));
  and2  gate303(.a(N147), .b(N99), .O(gate42inter2));
  inv1  gate304(.a(s_20), .O(gate42inter3));
  inv1  gate305(.a(s_21), .O(gate42inter4));
  nand2 gate306(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate307(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate308(.a(N99), .O(gate42inter7));
  inv1  gate309(.a(N147), .O(gate42inter8));
  nand2 gate310(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate311(.a(s_21), .b(gate42inter3), .O(gate42inter10));
  nor2  gate312(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate313(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate314(.a(gate42inter12), .b(gate42inter1), .O(N195));
nor2 gate43( .a(N105), .b(N147), .O(N196) );
nor2 gate44( .a(N112), .b(N151), .O(N197) );

  xor2  gate315(.a(N151), .b(N115), .O(gate45inter0));
  nand2 gate316(.a(gate45inter0), .b(s_22), .O(gate45inter1));
  and2  gate317(.a(N151), .b(N115), .O(gate45inter2));
  inv1  gate318(.a(s_22), .O(gate45inter3));
  inv1  gate319(.a(s_23), .O(gate45inter4));
  nand2 gate320(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate321(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate322(.a(N115), .O(gate45inter7));
  inv1  gate323(.a(N151), .O(gate45inter8));
  nand2 gate324(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate325(.a(s_23), .b(gate45inter3), .O(gate45inter10));
  nor2  gate326(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate327(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate328(.a(gate45inter12), .b(gate45inter1), .O(N198));
and9 gate46( .a(N154), .b(N159), .c(N162), .d(N165), .e(N168), .f(N171), .g(N174), .h(N177), .i(N180), .O(N199) );
inv1 gate47( .a(N199), .O(N203) );
inv1 gate48( .a(N199), .O(N213) );
inv1 gate49( .a(N199), .O(N223) );
xor2 gate50( .a(N203), .b(N154), .O(N224) );

  xor2  gate469(.a(N159), .b(N203), .O(gate51inter0));
  nand2 gate470(.a(gate51inter0), .b(s_44), .O(gate51inter1));
  and2  gate471(.a(N159), .b(N203), .O(gate51inter2));
  inv1  gate472(.a(s_44), .O(gate51inter3));
  inv1  gate473(.a(s_45), .O(gate51inter4));
  nand2 gate474(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate475(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate476(.a(N203), .O(gate51inter7));
  inv1  gate477(.a(N159), .O(gate51inter8));
  nand2 gate478(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate479(.a(s_45), .b(gate51inter3), .O(gate51inter10));
  nor2  gate480(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate481(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate482(.a(gate51inter12), .b(gate51inter1), .O(N227));

  xor2  gate329(.a(N162), .b(N203), .O(gate52inter0));
  nand2 gate330(.a(gate52inter0), .b(s_24), .O(gate52inter1));
  and2  gate331(.a(N162), .b(N203), .O(gate52inter2));
  inv1  gate332(.a(s_24), .O(gate52inter3));
  inv1  gate333(.a(s_25), .O(gate52inter4));
  nand2 gate334(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate335(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate336(.a(N203), .O(gate52inter7));
  inv1  gate337(.a(N162), .O(gate52inter8));
  nand2 gate338(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate339(.a(s_25), .b(gate52inter3), .O(gate52inter10));
  nor2  gate340(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate341(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate342(.a(gate52inter12), .b(gate52inter1), .O(N230));
xor2 gate53( .a(N203), .b(N165), .O(N233) );

  xor2  gate371(.a(N168), .b(N203), .O(gate54inter0));
  nand2 gate372(.a(gate54inter0), .b(s_30), .O(gate54inter1));
  and2  gate373(.a(N168), .b(N203), .O(gate54inter2));
  inv1  gate374(.a(s_30), .O(gate54inter3));
  inv1  gate375(.a(s_31), .O(gate54inter4));
  nand2 gate376(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate377(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate378(.a(N203), .O(gate54inter7));
  inv1  gate379(.a(N168), .O(gate54inter8));
  nand2 gate380(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate381(.a(s_31), .b(gate54inter3), .O(gate54inter10));
  nor2  gate382(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate383(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate384(.a(gate54inter12), .b(gate54inter1), .O(N236));
xor2 gate55( .a(N203), .b(N171), .O(N239) );
nand2 gate56( .a(N1), .b(N213), .O(N242) );
xor2 gate57( .a(N203), .b(N174), .O(N243) );
nand2 gate58( .a(N213), .b(N11), .O(N246) );
xor2 gate59( .a(N203), .b(N177), .O(N247) );
nand2 gate60( .a(N213), .b(N24), .O(N250) );
xor2 gate61( .a(N203), .b(N180), .O(N251) );
nand2 gate62( .a(N213), .b(N37), .O(N254) );
nand2 gate63( .a(N213), .b(N50), .O(N255) );
nand2 gate64( .a(N213), .b(N63), .O(N256) );
nand2 gate65( .a(N213), .b(N76), .O(N257) );
nand2 gate66( .a(N213), .b(N89), .O(N258) );
nand2 gate67( .a(N213), .b(N102), .O(N259) );

  xor2  gate455(.a(N157), .b(N224), .O(gate68inter0));
  nand2 gate456(.a(gate68inter0), .b(s_42), .O(gate68inter1));
  and2  gate457(.a(N157), .b(N224), .O(gate68inter2));
  inv1  gate458(.a(s_42), .O(gate68inter3));
  inv1  gate459(.a(s_43), .O(gate68inter4));
  nand2 gate460(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate461(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate462(.a(N224), .O(gate68inter7));
  inv1  gate463(.a(N157), .O(gate68inter8));
  nand2 gate464(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate465(.a(s_43), .b(gate68inter3), .O(gate68inter10));
  nor2  gate466(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate467(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate468(.a(gate68inter12), .b(gate68inter1), .O(N260));
nand2 gate69( .a(N224), .b(N158), .O(N263) );
nand2 gate70( .a(N227), .b(N183), .O(N264) );

  xor2  gate273(.a(N185), .b(N230), .O(gate71inter0));
  nand2 gate274(.a(gate71inter0), .b(s_16), .O(gate71inter1));
  and2  gate275(.a(N185), .b(N230), .O(gate71inter2));
  inv1  gate276(.a(s_16), .O(gate71inter3));
  inv1  gate277(.a(s_17), .O(gate71inter4));
  nand2 gate278(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate279(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate280(.a(N230), .O(gate71inter7));
  inv1  gate281(.a(N185), .O(gate71inter8));
  nand2 gate282(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate283(.a(s_17), .b(gate71inter3), .O(gate71inter10));
  nor2  gate284(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate285(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate286(.a(gate71inter12), .b(gate71inter1), .O(N267));
nand2 gate72( .a(N233), .b(N187), .O(N270) );
nand2 gate73( .a(N236), .b(N189), .O(N273) );
nand2 gate74( .a(N239), .b(N191), .O(N276) );

  xor2  gate539(.a(N193), .b(N243), .O(gate75inter0));
  nand2 gate540(.a(gate75inter0), .b(s_54), .O(gate75inter1));
  and2  gate541(.a(N193), .b(N243), .O(gate75inter2));
  inv1  gate542(.a(s_54), .O(gate75inter3));
  inv1  gate543(.a(s_55), .O(gate75inter4));
  nand2 gate544(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate545(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate546(.a(N243), .O(gate75inter7));
  inv1  gate547(.a(N193), .O(gate75inter8));
  nand2 gate548(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate549(.a(s_55), .b(gate75inter3), .O(gate75inter10));
  nor2  gate550(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate551(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate552(.a(gate75inter12), .b(gate75inter1), .O(N279));

  xor2  gate567(.a(N195), .b(N247), .O(gate76inter0));
  nand2 gate568(.a(gate76inter0), .b(s_58), .O(gate76inter1));
  and2  gate569(.a(N195), .b(N247), .O(gate76inter2));
  inv1  gate570(.a(s_58), .O(gate76inter3));
  inv1  gate571(.a(s_59), .O(gate76inter4));
  nand2 gate572(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate573(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate574(.a(N247), .O(gate76inter7));
  inv1  gate575(.a(N195), .O(gate76inter8));
  nand2 gate576(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate577(.a(s_59), .b(gate76inter3), .O(gate76inter10));
  nor2  gate578(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate579(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate580(.a(gate76inter12), .b(gate76inter1), .O(N282));
nand2 gate77( .a(N251), .b(N197), .O(N285) );

  xor2  gate357(.a(N184), .b(N227), .O(gate78inter0));
  nand2 gate358(.a(gate78inter0), .b(s_28), .O(gate78inter1));
  and2  gate359(.a(N184), .b(N227), .O(gate78inter2));
  inv1  gate360(.a(s_28), .O(gate78inter3));
  inv1  gate361(.a(s_29), .O(gate78inter4));
  nand2 gate362(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate363(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate364(.a(N227), .O(gate78inter7));
  inv1  gate365(.a(N184), .O(gate78inter8));
  nand2 gate366(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate367(.a(s_29), .b(gate78inter3), .O(gate78inter10));
  nor2  gate368(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate369(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate370(.a(gate78inter12), .b(gate78inter1), .O(N288));
nand2 gate79( .a(N230), .b(N186), .O(N289) );
nand2 gate80( .a(N233), .b(N188), .O(N290) );
nand2 gate81( .a(N236), .b(N190), .O(N291) );
nand2 gate82( .a(N239), .b(N192), .O(N292) );
nand2 gate83( .a(N243), .b(N194), .O(N293) );

  xor2  gate553(.a(N196), .b(N247), .O(gate84inter0));
  nand2 gate554(.a(gate84inter0), .b(s_56), .O(gate84inter1));
  and2  gate555(.a(N196), .b(N247), .O(gate84inter2));
  inv1  gate556(.a(s_56), .O(gate84inter3));
  inv1  gate557(.a(s_57), .O(gate84inter4));
  nand2 gate558(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate559(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate560(.a(N247), .O(gate84inter7));
  inv1  gate561(.a(N196), .O(gate84inter8));
  nand2 gate562(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate563(.a(s_57), .b(gate84inter3), .O(gate84inter10));
  nor2  gate564(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate565(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate566(.a(gate84inter12), .b(gate84inter1), .O(N294));

  xor2  gate203(.a(N198), .b(N251), .O(gate85inter0));
  nand2 gate204(.a(gate85inter0), .b(s_6), .O(gate85inter1));
  and2  gate205(.a(N198), .b(N251), .O(gate85inter2));
  inv1  gate206(.a(s_6), .O(gate85inter3));
  inv1  gate207(.a(s_7), .O(gate85inter4));
  nand2 gate208(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate209(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate210(.a(N251), .O(gate85inter7));
  inv1  gate211(.a(N198), .O(gate85inter8));
  nand2 gate212(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate213(.a(s_7), .b(gate85inter3), .O(gate85inter10));
  nor2  gate214(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate215(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate216(.a(gate85inter12), .b(gate85inter1), .O(N295));
and9 gate86( .a(N260), .b(N264), .c(N267), .d(N270), .e(N273), .f(N276), .g(N279), .h(N282), .i(N285), .O(N296) );
inv1 gate87( .a(N263), .O(N300) );
inv1 gate88( .a(N288), .O(N301) );
inv1 gate89( .a(N289), .O(N302) );
inv1 gate90( .a(N290), .O(N303) );
inv1 gate91( .a(N291), .O(N304) );
inv1 gate92( .a(N292), .O(N305) );
inv1 gate93( .a(N293), .O(N306) );
inv1 gate94( .a(N294), .O(N307) );
inv1 gate95( .a(N295), .O(N308) );
inv1 gate96( .a(N296), .O(N309) );
inv1 gate97( .a(N296), .O(N319) );
inv1 gate98( .a(N296), .O(N329) );
xor2 gate99( .a(N309), .b(N260), .O(N330) );

  xor2  gate497(.a(N264), .b(N309), .O(gate100inter0));
  nand2 gate498(.a(gate100inter0), .b(s_48), .O(gate100inter1));
  and2  gate499(.a(N264), .b(N309), .O(gate100inter2));
  inv1  gate500(.a(s_48), .O(gate100inter3));
  inv1  gate501(.a(s_49), .O(gate100inter4));
  nand2 gate502(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate503(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate504(.a(N309), .O(gate100inter7));
  inv1  gate505(.a(N264), .O(gate100inter8));
  nand2 gate506(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate507(.a(s_49), .b(gate100inter3), .O(gate100inter10));
  nor2  gate508(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate509(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate510(.a(gate100inter12), .b(gate100inter1), .O(N331));

  xor2  gate161(.a(N267), .b(N309), .O(gate101inter0));
  nand2 gate162(.a(gate101inter0), .b(s_0), .O(gate101inter1));
  and2  gate163(.a(N267), .b(N309), .O(gate101inter2));
  inv1  gate164(.a(s_0), .O(gate101inter3));
  inv1  gate165(.a(s_1), .O(gate101inter4));
  nand2 gate166(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate167(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate168(.a(N309), .O(gate101inter7));
  inv1  gate169(.a(N267), .O(gate101inter8));
  nand2 gate170(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate171(.a(s_1), .b(gate101inter3), .O(gate101inter10));
  nor2  gate172(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate173(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate174(.a(gate101inter12), .b(gate101inter1), .O(N332));
xor2 gate102( .a(N309), .b(N270), .O(N333) );
nand2 gate103( .a(N8), .b(N319), .O(N334) );
xor2 gate104( .a(N309), .b(N273), .O(N335) );
nand2 gate105( .a(N319), .b(N21), .O(N336) );
xor2 gate106( .a(N309), .b(N276), .O(N337) );

  xor2  gate413(.a(N34), .b(N319), .O(gate107inter0));
  nand2 gate414(.a(gate107inter0), .b(s_36), .O(gate107inter1));
  and2  gate415(.a(N34), .b(N319), .O(gate107inter2));
  inv1  gate416(.a(s_36), .O(gate107inter3));
  inv1  gate417(.a(s_37), .O(gate107inter4));
  nand2 gate418(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate419(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate420(.a(N319), .O(gate107inter7));
  inv1  gate421(.a(N34), .O(gate107inter8));
  nand2 gate422(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate423(.a(s_37), .b(gate107inter3), .O(gate107inter10));
  nor2  gate424(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate425(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate426(.a(gate107inter12), .b(gate107inter1), .O(N338));
xor2 gate108( .a(N309), .b(N279), .O(N339) );
nand2 gate109( .a(N319), .b(N47), .O(N340) );
xor2 gate110( .a(N309), .b(N282), .O(N341) );
nand2 gate111( .a(N319), .b(N60), .O(N342) );
xor2 gate112( .a(N309), .b(N285), .O(N343) );
nand2 gate113( .a(N319), .b(N73), .O(N344) );
nand2 gate114( .a(N319), .b(N86), .O(N345) );
nand2 gate115( .a(N319), .b(N99), .O(N346) );
nand2 gate116( .a(N319), .b(N112), .O(N347) );

  xor2  gate189(.a(N300), .b(N330), .O(gate117inter0));
  nand2 gate190(.a(gate117inter0), .b(s_4), .O(gate117inter1));
  and2  gate191(.a(N300), .b(N330), .O(gate117inter2));
  inv1  gate192(.a(s_4), .O(gate117inter3));
  inv1  gate193(.a(s_5), .O(gate117inter4));
  nand2 gate194(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate195(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate196(.a(N330), .O(gate117inter7));
  inv1  gate197(.a(N300), .O(gate117inter8));
  nand2 gate198(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate199(.a(s_5), .b(gate117inter3), .O(gate117inter10));
  nor2  gate200(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate201(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate202(.a(gate117inter12), .b(gate117inter1), .O(N348));
nand2 gate118( .a(N331), .b(N301), .O(N349) );
nand2 gate119( .a(N332), .b(N302), .O(N350) );

  xor2  gate343(.a(N303), .b(N333), .O(gate120inter0));
  nand2 gate344(.a(gate120inter0), .b(s_26), .O(gate120inter1));
  and2  gate345(.a(N303), .b(N333), .O(gate120inter2));
  inv1  gate346(.a(s_26), .O(gate120inter3));
  inv1  gate347(.a(s_27), .O(gate120inter4));
  nand2 gate348(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate349(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate350(.a(N333), .O(gate120inter7));
  inv1  gate351(.a(N303), .O(gate120inter8));
  nand2 gate352(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate353(.a(s_27), .b(gate120inter3), .O(gate120inter10));
  nor2  gate354(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate355(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate356(.a(gate120inter12), .b(gate120inter1), .O(N351));

  xor2  gate245(.a(N304), .b(N335), .O(gate121inter0));
  nand2 gate246(.a(gate121inter0), .b(s_12), .O(gate121inter1));
  and2  gate247(.a(N304), .b(N335), .O(gate121inter2));
  inv1  gate248(.a(s_12), .O(gate121inter3));
  inv1  gate249(.a(s_13), .O(gate121inter4));
  nand2 gate250(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate251(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate252(.a(N335), .O(gate121inter7));
  inv1  gate253(.a(N304), .O(gate121inter8));
  nand2 gate254(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate255(.a(s_13), .b(gate121inter3), .O(gate121inter10));
  nor2  gate256(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate257(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate258(.a(gate121inter12), .b(gate121inter1), .O(N352));
nand2 gate122( .a(N337), .b(N305), .O(N353) );
nand2 gate123( .a(N339), .b(N306), .O(N354) );
nand2 gate124( .a(N341), .b(N307), .O(N355) );
nand2 gate125( .a(N343), .b(N308), .O(N356) );
and9 gate126( .a(N348), .b(N349), .c(N350), .d(N351), .e(N352), .f(N353), .g(N354), .h(N355), .i(N356), .O(N357) );
inv1 gate127( .a(N357), .O(N360) );
inv1 gate128( .a(N357), .O(N370) );

  xor2  gate427(.a(N360), .b(N14), .O(gate129inter0));
  nand2 gate428(.a(gate129inter0), .b(s_38), .O(gate129inter1));
  and2  gate429(.a(N360), .b(N14), .O(gate129inter2));
  inv1  gate430(.a(s_38), .O(gate129inter3));
  inv1  gate431(.a(s_39), .O(gate129inter4));
  nand2 gate432(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate433(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate434(.a(N14), .O(gate129inter7));
  inv1  gate435(.a(N360), .O(gate129inter8));
  nand2 gate436(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate437(.a(s_39), .b(gate129inter3), .O(gate129inter10));
  nor2  gate438(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate439(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate440(.a(gate129inter12), .b(gate129inter1), .O(N371));
nand2 gate130( .a(N360), .b(N27), .O(N372) );
nand2 gate131( .a(N360), .b(N40), .O(N373) );
nand2 gate132( .a(N360), .b(N53), .O(N374) );

  xor2  gate399(.a(N66), .b(N360), .O(gate133inter0));
  nand2 gate400(.a(gate133inter0), .b(s_34), .O(gate133inter1));
  and2  gate401(.a(N66), .b(N360), .O(gate133inter2));
  inv1  gate402(.a(s_34), .O(gate133inter3));
  inv1  gate403(.a(s_35), .O(gate133inter4));
  nand2 gate404(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate405(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate406(.a(N360), .O(gate133inter7));
  inv1  gate407(.a(N66), .O(gate133inter8));
  nand2 gate408(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate409(.a(s_35), .b(gate133inter3), .O(gate133inter10));
  nor2  gate410(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate411(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate412(.a(gate133inter12), .b(gate133inter1), .O(N375));
nand2 gate134( .a(N360), .b(N79), .O(N376) );

  xor2  gate259(.a(N92), .b(N360), .O(gate135inter0));
  nand2 gate260(.a(gate135inter0), .b(s_14), .O(gate135inter1));
  and2  gate261(.a(N92), .b(N360), .O(gate135inter2));
  inv1  gate262(.a(s_14), .O(gate135inter3));
  inv1  gate263(.a(s_15), .O(gate135inter4));
  nand2 gate264(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate265(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate266(.a(N360), .O(gate135inter7));
  inv1  gate267(.a(N92), .O(gate135inter8));
  nand2 gate268(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate269(.a(s_15), .b(gate135inter3), .O(gate135inter10));
  nor2  gate270(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate271(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate272(.a(gate135inter12), .b(gate135inter1), .O(N377));
nand2 gate136( .a(N360), .b(N105), .O(N378) );
nand2 gate137( .a(N360), .b(N115), .O(N379) );
nand4 gate138( .a(N4), .b(N242), .c(N334), .d(N371), .O(N380) );
nand4 gate139( .a(N246), .b(N336), .c(N372), .d(N17), .O(N381) );
nand4 gate140( .a(N250), .b(N338), .c(N373), .d(N30), .O(N386) );
nand4 gate141( .a(N254), .b(N340), .c(N374), .d(N43), .O(N393) );
nand4 gate142( .a(N255), .b(N342), .c(N375), .d(N56), .O(N399) );
nand4 gate143( .a(N256), .b(N344), .c(N376), .d(N69), .O(N404) );
nand4 gate144( .a(N257), .b(N345), .c(N377), .d(N82), .O(N407) );
nand4 gate145( .a(N258), .b(N346), .c(N378), .d(N95), .O(N411) );
nand4 gate146( .a(N259), .b(N347), .c(N379), .d(N108), .O(N414) );
inv1 gate147( .a(N380), .O(N415) );
and8 gate148( .a(N381), .b(N386), .c(N393), .d(N399), .e(N404), .f(N407), .g(N411), .h(N414), .O(N416) );
inv1 gate149( .a(N393), .O(N417) );
inv1 gate150( .a(N404), .O(N418) );
inv1 gate151( .a(N407), .O(N419) );
inv1 gate152( .a(N411), .O(N420) );

  xor2  gate287(.a(N416), .b(N415), .O(gate153inter0));
  nand2 gate288(.a(gate153inter0), .b(s_18), .O(gate153inter1));
  and2  gate289(.a(N416), .b(N415), .O(gate153inter2));
  inv1  gate290(.a(s_18), .O(gate153inter3));
  inv1  gate291(.a(s_19), .O(gate153inter4));
  nand2 gate292(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate293(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate294(.a(N415), .O(gate153inter7));
  inv1  gate295(.a(N416), .O(gate153inter8));
  nand2 gate296(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate297(.a(s_19), .b(gate153inter3), .O(gate153inter10));
  nor2  gate298(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate299(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate300(.a(gate153inter12), .b(gate153inter1), .O(N421));

  xor2  gate175(.a(N417), .b(N386), .O(gate154inter0));
  nand2 gate176(.a(gate154inter0), .b(s_2), .O(gate154inter1));
  and2  gate177(.a(N417), .b(N386), .O(gate154inter2));
  inv1  gate178(.a(s_2), .O(gate154inter3));
  inv1  gate179(.a(s_3), .O(gate154inter4));
  nand2 gate180(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate181(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate182(.a(N386), .O(gate154inter7));
  inv1  gate183(.a(N417), .O(gate154inter8));
  nand2 gate184(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate185(.a(s_3), .b(gate154inter3), .O(gate154inter10));
  nor2  gate186(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate187(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate188(.a(gate154inter12), .b(gate154inter1), .O(N422));
nand4 gate155( .a(N386), .b(N393), .c(N418), .d(N399), .O(N425) );
nand3 gate156( .a(N399), .b(N393), .c(N419), .O(N428) );
nand4 gate157( .a(N386), .b(N393), .c(N407), .d(N420), .O(N429) );
nand4 gate158( .a(N381), .b(N386), .c(N422), .d(N399), .O(N430) );
nand4 gate159( .a(N381), .b(N386), .c(N425), .d(N428), .O(N431) );
nand4 gate160( .a(N381), .b(N422), .c(N425), .d(N429), .O(N432) );

endmodule