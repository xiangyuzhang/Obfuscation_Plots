module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate497inter0, gate497inter1, gate497inter2, gate497inter3, gate497inter4, gate497inter5, gate497inter6, gate497inter7, gate497inter8, gate497inter9, gate497inter10, gate497inter11, gate497inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate1289(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate1290(.a(gate16inter0), .b(s_106), .O(gate16inter1));
  and2  gate1291(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate1292(.a(s_106), .O(gate16inter3));
  inv1  gate1293(.a(s_107), .O(gate16inter4));
  nand2 gate1294(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate1295(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate1296(.a(G15), .O(gate16inter7));
  inv1  gate1297(.a(G16), .O(gate16inter8));
  nand2 gate1298(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate1299(.a(s_107), .b(gate16inter3), .O(gate16inter10));
  nor2  gate1300(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate1301(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate1302(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate771(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate772(.a(gate21inter0), .b(s_32), .O(gate21inter1));
  and2  gate773(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate774(.a(s_32), .O(gate21inter3));
  inv1  gate775(.a(s_33), .O(gate21inter4));
  nand2 gate776(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate777(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate778(.a(G25), .O(gate21inter7));
  inv1  gate779(.a(G26), .O(gate21inter8));
  nand2 gate780(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate781(.a(s_33), .b(gate21inter3), .O(gate21inter10));
  nor2  gate782(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate783(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate784(.a(gate21inter12), .b(gate21inter1), .O(G302));

  xor2  gate799(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate800(.a(gate22inter0), .b(s_36), .O(gate22inter1));
  and2  gate801(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate802(.a(s_36), .O(gate22inter3));
  inv1  gate803(.a(s_37), .O(gate22inter4));
  nand2 gate804(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate805(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate806(.a(G27), .O(gate22inter7));
  inv1  gate807(.a(G28), .O(gate22inter8));
  nand2 gate808(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate809(.a(s_37), .b(gate22inter3), .O(gate22inter10));
  nor2  gate810(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate811(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate812(.a(gate22inter12), .b(gate22inter1), .O(G305));
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate1191(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate1192(.a(gate29inter0), .b(s_92), .O(gate29inter1));
  and2  gate1193(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate1194(.a(s_92), .O(gate29inter3));
  inv1  gate1195(.a(s_93), .O(gate29inter4));
  nand2 gate1196(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate1197(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate1198(.a(G3), .O(gate29inter7));
  inv1  gate1199(.a(G7), .O(gate29inter8));
  nand2 gate1200(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate1201(.a(s_93), .b(gate29inter3), .O(gate29inter10));
  nor2  gate1202(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate1203(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate1204(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate1163(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate1164(.a(gate34inter0), .b(s_88), .O(gate34inter1));
  and2  gate1165(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate1166(.a(s_88), .O(gate34inter3));
  inv1  gate1167(.a(s_89), .O(gate34inter4));
  nand2 gate1168(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate1169(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate1170(.a(G25), .O(gate34inter7));
  inv1  gate1171(.a(G29), .O(gate34inter8));
  nand2 gate1172(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate1173(.a(s_89), .b(gate34inter3), .O(gate34inter10));
  nor2  gate1174(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate1175(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate1176(.a(gate34inter12), .b(gate34inter1), .O(G341));

  xor2  gate2087(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate2088(.a(gate35inter0), .b(s_220), .O(gate35inter1));
  and2  gate2089(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate2090(.a(s_220), .O(gate35inter3));
  inv1  gate2091(.a(s_221), .O(gate35inter4));
  nand2 gate2092(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate2093(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate2094(.a(G18), .O(gate35inter7));
  inv1  gate2095(.a(G22), .O(gate35inter8));
  nand2 gate2096(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate2097(.a(s_221), .b(gate35inter3), .O(gate35inter10));
  nor2  gate2098(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate2099(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate2100(.a(gate35inter12), .b(gate35inter1), .O(G344));

  xor2  gate603(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate604(.a(gate36inter0), .b(s_8), .O(gate36inter1));
  and2  gate605(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate606(.a(s_8), .O(gate36inter3));
  inv1  gate607(.a(s_9), .O(gate36inter4));
  nand2 gate608(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate609(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate610(.a(G26), .O(gate36inter7));
  inv1  gate611(.a(G30), .O(gate36inter8));
  nand2 gate612(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate613(.a(s_9), .b(gate36inter3), .O(gate36inter10));
  nor2  gate614(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate615(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate616(.a(gate36inter12), .b(gate36inter1), .O(G347));

  xor2  gate939(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate940(.a(gate37inter0), .b(s_56), .O(gate37inter1));
  and2  gate941(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate942(.a(s_56), .O(gate37inter3));
  inv1  gate943(.a(s_57), .O(gate37inter4));
  nand2 gate944(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate945(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate946(.a(G19), .O(gate37inter7));
  inv1  gate947(.a(G23), .O(gate37inter8));
  nand2 gate948(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate949(.a(s_57), .b(gate37inter3), .O(gate37inter10));
  nor2  gate950(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate951(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate952(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate869(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate870(.a(gate39inter0), .b(s_46), .O(gate39inter1));
  and2  gate871(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate872(.a(s_46), .O(gate39inter3));
  inv1  gate873(.a(s_47), .O(gate39inter4));
  nand2 gate874(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate875(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate876(.a(G20), .O(gate39inter7));
  inv1  gate877(.a(G24), .O(gate39inter8));
  nand2 gate878(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate879(.a(s_47), .b(gate39inter3), .O(gate39inter10));
  nor2  gate880(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate881(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate882(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate1709(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate1710(.a(gate41inter0), .b(s_166), .O(gate41inter1));
  and2  gate1711(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate1712(.a(s_166), .O(gate41inter3));
  inv1  gate1713(.a(s_167), .O(gate41inter4));
  nand2 gate1714(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate1715(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate1716(.a(G1), .O(gate41inter7));
  inv1  gate1717(.a(G266), .O(gate41inter8));
  nand2 gate1718(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate1719(.a(s_167), .b(gate41inter3), .O(gate41inter10));
  nor2  gate1720(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate1721(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate1722(.a(gate41inter12), .b(gate41inter1), .O(G362));

  xor2  gate1849(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate1850(.a(gate42inter0), .b(s_186), .O(gate42inter1));
  and2  gate1851(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate1852(.a(s_186), .O(gate42inter3));
  inv1  gate1853(.a(s_187), .O(gate42inter4));
  nand2 gate1854(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate1855(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate1856(.a(G2), .O(gate42inter7));
  inv1  gate1857(.a(G266), .O(gate42inter8));
  nand2 gate1858(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate1859(.a(s_187), .b(gate42inter3), .O(gate42inter10));
  nor2  gate1860(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate1861(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate1862(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );

  xor2  gate1415(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate1416(.a(gate47inter0), .b(s_124), .O(gate47inter1));
  and2  gate1417(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate1418(.a(s_124), .O(gate47inter3));
  inv1  gate1419(.a(s_125), .O(gate47inter4));
  nand2 gate1420(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate1421(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate1422(.a(G7), .O(gate47inter7));
  inv1  gate1423(.a(G275), .O(gate47inter8));
  nand2 gate1424(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate1425(.a(s_125), .b(gate47inter3), .O(gate47inter10));
  nor2  gate1426(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate1427(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate1428(.a(gate47inter12), .b(gate47inter1), .O(G368));
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate1009(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate1010(.a(gate51inter0), .b(s_66), .O(gate51inter1));
  and2  gate1011(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate1012(.a(s_66), .O(gate51inter3));
  inv1  gate1013(.a(s_67), .O(gate51inter4));
  nand2 gate1014(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate1015(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate1016(.a(G11), .O(gate51inter7));
  inv1  gate1017(.a(G281), .O(gate51inter8));
  nand2 gate1018(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate1019(.a(s_67), .b(gate51inter3), .O(gate51inter10));
  nor2  gate1020(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate1021(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate1022(.a(gate51inter12), .b(gate51inter1), .O(G372));

  xor2  gate1975(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate1976(.a(gate52inter0), .b(s_204), .O(gate52inter1));
  and2  gate1977(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate1978(.a(s_204), .O(gate52inter3));
  inv1  gate1979(.a(s_205), .O(gate52inter4));
  nand2 gate1980(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate1981(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate1982(.a(G12), .O(gate52inter7));
  inv1  gate1983(.a(G281), .O(gate52inter8));
  nand2 gate1984(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate1985(.a(s_205), .b(gate52inter3), .O(gate52inter10));
  nor2  gate1986(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate1987(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate1988(.a(gate52inter12), .b(gate52inter1), .O(G373));

  xor2  gate2045(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate2046(.a(gate53inter0), .b(s_214), .O(gate53inter1));
  and2  gate2047(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate2048(.a(s_214), .O(gate53inter3));
  inv1  gate2049(.a(s_215), .O(gate53inter4));
  nand2 gate2050(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate2051(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate2052(.a(G13), .O(gate53inter7));
  inv1  gate2053(.a(G284), .O(gate53inter8));
  nand2 gate2054(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate2055(.a(s_215), .b(gate53inter3), .O(gate53inter10));
  nor2  gate2056(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate2057(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate2058(.a(gate53inter12), .b(gate53inter1), .O(G374));

  xor2  gate1807(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate1808(.a(gate54inter0), .b(s_180), .O(gate54inter1));
  and2  gate1809(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate1810(.a(s_180), .O(gate54inter3));
  inv1  gate1811(.a(s_181), .O(gate54inter4));
  nand2 gate1812(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate1813(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate1814(.a(G14), .O(gate54inter7));
  inv1  gate1815(.a(G284), .O(gate54inter8));
  nand2 gate1816(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate1817(.a(s_181), .b(gate54inter3), .O(gate54inter10));
  nor2  gate1818(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate1819(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate1820(.a(gate54inter12), .b(gate54inter1), .O(G375));

  xor2  gate757(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate758(.a(gate55inter0), .b(s_30), .O(gate55inter1));
  and2  gate759(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate760(.a(s_30), .O(gate55inter3));
  inv1  gate761(.a(s_31), .O(gate55inter4));
  nand2 gate762(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate763(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate764(.a(G15), .O(gate55inter7));
  inv1  gate765(.a(G287), .O(gate55inter8));
  nand2 gate766(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate767(.a(s_31), .b(gate55inter3), .O(gate55inter10));
  nor2  gate768(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate769(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate770(.a(gate55inter12), .b(gate55inter1), .O(G376));
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate1051(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate1052(.a(gate59inter0), .b(s_72), .O(gate59inter1));
  and2  gate1053(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate1054(.a(s_72), .O(gate59inter3));
  inv1  gate1055(.a(s_73), .O(gate59inter4));
  nand2 gate1056(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate1057(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate1058(.a(G19), .O(gate59inter7));
  inv1  gate1059(.a(G293), .O(gate59inter8));
  nand2 gate1060(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate1061(.a(s_73), .b(gate59inter3), .O(gate59inter10));
  nor2  gate1062(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate1063(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate1064(.a(gate59inter12), .b(gate59inter1), .O(G380));

  xor2  gate967(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate968(.a(gate60inter0), .b(s_60), .O(gate60inter1));
  and2  gate969(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate970(.a(s_60), .O(gate60inter3));
  inv1  gate971(.a(s_61), .O(gate60inter4));
  nand2 gate972(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate973(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate974(.a(G20), .O(gate60inter7));
  inv1  gate975(.a(G293), .O(gate60inter8));
  nand2 gate976(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate977(.a(s_61), .b(gate60inter3), .O(gate60inter10));
  nor2  gate978(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate979(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate980(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate2115(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate2116(.a(gate67inter0), .b(s_224), .O(gate67inter1));
  and2  gate2117(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate2118(.a(s_224), .O(gate67inter3));
  inv1  gate2119(.a(s_225), .O(gate67inter4));
  nand2 gate2120(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate2121(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate2122(.a(G27), .O(gate67inter7));
  inv1  gate2123(.a(G305), .O(gate67inter8));
  nand2 gate2124(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate2125(.a(s_225), .b(gate67inter3), .O(gate67inter10));
  nor2  gate2126(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate2127(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate2128(.a(gate67inter12), .b(gate67inter1), .O(G388));

  xor2  gate1205(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate1206(.a(gate68inter0), .b(s_94), .O(gate68inter1));
  and2  gate1207(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate1208(.a(s_94), .O(gate68inter3));
  inv1  gate1209(.a(s_95), .O(gate68inter4));
  nand2 gate1210(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate1211(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate1212(.a(G28), .O(gate68inter7));
  inv1  gate1213(.a(G305), .O(gate68inter8));
  nand2 gate1214(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate1215(.a(s_95), .b(gate68inter3), .O(gate68inter10));
  nor2  gate1216(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate1217(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate1218(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate2157(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate2158(.a(gate70inter0), .b(s_230), .O(gate70inter1));
  and2  gate2159(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate2160(.a(s_230), .O(gate70inter3));
  inv1  gate2161(.a(s_231), .O(gate70inter4));
  nand2 gate2162(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate2163(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate2164(.a(G30), .O(gate70inter7));
  inv1  gate2165(.a(G308), .O(gate70inter8));
  nand2 gate2166(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate2167(.a(s_231), .b(gate70inter3), .O(gate70inter10));
  nor2  gate2168(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate2169(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate2170(.a(gate70inter12), .b(gate70inter1), .O(G391));

  xor2  gate1037(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate1038(.a(gate71inter0), .b(s_70), .O(gate71inter1));
  and2  gate1039(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate1040(.a(s_70), .O(gate71inter3));
  inv1  gate1041(.a(s_71), .O(gate71inter4));
  nand2 gate1042(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate1043(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate1044(.a(G31), .O(gate71inter7));
  inv1  gate1045(.a(G311), .O(gate71inter8));
  nand2 gate1046(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate1047(.a(s_71), .b(gate71inter3), .O(gate71inter10));
  nor2  gate1048(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate1049(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate1050(.a(gate71inter12), .b(gate71inter1), .O(G392));

  xor2  gate1247(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate1248(.a(gate72inter0), .b(s_100), .O(gate72inter1));
  and2  gate1249(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate1250(.a(s_100), .O(gate72inter3));
  inv1  gate1251(.a(s_101), .O(gate72inter4));
  nand2 gate1252(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate1253(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate1254(.a(G32), .O(gate72inter7));
  inv1  gate1255(.a(G311), .O(gate72inter8));
  nand2 gate1256(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate1257(.a(s_101), .b(gate72inter3), .O(gate72inter10));
  nor2  gate1258(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate1259(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate1260(.a(gate72inter12), .b(gate72inter1), .O(G393));
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate841(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate842(.a(gate74inter0), .b(s_42), .O(gate74inter1));
  and2  gate843(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate844(.a(s_42), .O(gate74inter3));
  inv1  gate845(.a(s_43), .O(gate74inter4));
  nand2 gate846(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate847(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate848(.a(G5), .O(gate74inter7));
  inv1  gate849(.a(G314), .O(gate74inter8));
  nand2 gate850(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate851(.a(s_43), .b(gate74inter3), .O(gate74inter10));
  nor2  gate852(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate853(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate854(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate855(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate856(.a(gate77inter0), .b(s_44), .O(gate77inter1));
  and2  gate857(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate858(.a(s_44), .O(gate77inter3));
  inv1  gate859(.a(s_45), .O(gate77inter4));
  nand2 gate860(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate861(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate862(.a(G2), .O(gate77inter7));
  inv1  gate863(.a(G320), .O(gate77inter8));
  nand2 gate864(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate865(.a(s_45), .b(gate77inter3), .O(gate77inter10));
  nor2  gate866(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate867(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate868(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );

  xor2  gate2059(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate2060(.a(gate79inter0), .b(s_216), .O(gate79inter1));
  and2  gate2061(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate2062(.a(s_216), .O(gate79inter3));
  inv1  gate2063(.a(s_217), .O(gate79inter4));
  nand2 gate2064(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate2065(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate2066(.a(G10), .O(gate79inter7));
  inv1  gate2067(.a(G323), .O(gate79inter8));
  nand2 gate2068(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate2069(.a(s_217), .b(gate79inter3), .O(gate79inter10));
  nor2  gate2070(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate2071(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate2072(.a(gate79inter12), .b(gate79inter1), .O(G400));
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate701(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate702(.a(gate81inter0), .b(s_22), .O(gate81inter1));
  and2  gate703(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate704(.a(s_22), .O(gate81inter3));
  inv1  gate705(.a(s_23), .O(gate81inter4));
  nand2 gate706(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate707(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate708(.a(G3), .O(gate81inter7));
  inv1  gate709(.a(G326), .O(gate81inter8));
  nand2 gate710(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate711(.a(s_23), .b(gate81inter3), .O(gate81inter10));
  nor2  gate712(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate713(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate714(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate1723(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate1724(.a(gate94inter0), .b(s_168), .O(gate94inter1));
  and2  gate1725(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate1726(.a(s_168), .O(gate94inter3));
  inv1  gate1727(.a(s_169), .O(gate94inter4));
  nand2 gate1728(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate1729(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate1730(.a(G22), .O(gate94inter7));
  inv1  gate1731(.a(G344), .O(gate94inter8));
  nand2 gate1732(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate1733(.a(s_169), .b(gate94inter3), .O(gate94inter10));
  nor2  gate1734(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate1735(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate1736(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );

  xor2  gate1737(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate1738(.a(gate96inter0), .b(s_170), .O(gate96inter1));
  and2  gate1739(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate1740(.a(s_170), .O(gate96inter3));
  inv1  gate1741(.a(s_171), .O(gate96inter4));
  nand2 gate1742(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate1743(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate1744(.a(G30), .O(gate96inter7));
  inv1  gate1745(.a(G347), .O(gate96inter8));
  nand2 gate1746(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate1747(.a(s_171), .b(gate96inter3), .O(gate96inter10));
  nor2  gate1748(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate1749(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate1750(.a(gate96inter12), .b(gate96inter1), .O(G417));
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate1779(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate1780(.a(gate98inter0), .b(s_176), .O(gate98inter1));
  and2  gate1781(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate1782(.a(s_176), .O(gate98inter3));
  inv1  gate1783(.a(s_177), .O(gate98inter4));
  nand2 gate1784(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1785(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1786(.a(G23), .O(gate98inter7));
  inv1  gate1787(.a(G350), .O(gate98inter8));
  nand2 gate1788(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1789(.a(s_177), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1790(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1791(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1792(.a(gate98inter12), .b(gate98inter1), .O(G419));

  xor2  gate631(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate632(.a(gate99inter0), .b(s_12), .O(gate99inter1));
  and2  gate633(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate634(.a(s_12), .O(gate99inter3));
  inv1  gate635(.a(s_13), .O(gate99inter4));
  nand2 gate636(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate637(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate638(.a(G27), .O(gate99inter7));
  inv1  gate639(.a(G353), .O(gate99inter8));
  nand2 gate640(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate641(.a(s_13), .b(gate99inter3), .O(gate99inter10));
  nor2  gate642(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate643(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate644(.a(gate99inter12), .b(gate99inter1), .O(G420));

  xor2  gate1443(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate1444(.a(gate100inter0), .b(s_128), .O(gate100inter1));
  and2  gate1445(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate1446(.a(s_128), .O(gate100inter3));
  inv1  gate1447(.a(s_129), .O(gate100inter4));
  nand2 gate1448(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate1449(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate1450(.a(G31), .O(gate100inter7));
  inv1  gate1451(.a(G353), .O(gate100inter8));
  nand2 gate1452(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate1453(.a(s_129), .b(gate100inter3), .O(gate100inter10));
  nor2  gate1454(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate1455(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate1456(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );

  xor2  gate1359(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate1360(.a(gate103inter0), .b(s_116), .O(gate103inter1));
  and2  gate1361(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate1362(.a(s_116), .O(gate103inter3));
  inv1  gate1363(.a(s_117), .O(gate103inter4));
  nand2 gate1364(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate1365(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate1366(.a(G28), .O(gate103inter7));
  inv1  gate1367(.a(G359), .O(gate103inter8));
  nand2 gate1368(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate1369(.a(s_117), .b(gate103inter3), .O(gate103inter10));
  nor2  gate1370(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate1371(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate1372(.a(gate103inter12), .b(gate103inter1), .O(G424));
nand2 gate104( .a(G32), .b(G359), .O(G425) );

  xor2  gate1303(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate1304(.a(gate105inter0), .b(s_108), .O(gate105inter1));
  and2  gate1305(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate1306(.a(s_108), .O(gate105inter3));
  inv1  gate1307(.a(s_109), .O(gate105inter4));
  nand2 gate1308(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate1309(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate1310(.a(G362), .O(gate105inter7));
  inv1  gate1311(.a(G363), .O(gate105inter8));
  nand2 gate1312(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate1313(.a(s_109), .b(gate105inter3), .O(gate105inter10));
  nor2  gate1314(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate1315(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate1316(.a(gate105inter12), .b(gate105inter1), .O(G426));

  xor2  gate1485(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate1486(.a(gate106inter0), .b(s_134), .O(gate106inter1));
  and2  gate1487(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate1488(.a(s_134), .O(gate106inter3));
  inv1  gate1489(.a(s_135), .O(gate106inter4));
  nand2 gate1490(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate1491(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate1492(.a(G364), .O(gate106inter7));
  inv1  gate1493(.a(G365), .O(gate106inter8));
  nand2 gate1494(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate1495(.a(s_135), .b(gate106inter3), .O(gate106inter10));
  nor2  gate1496(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate1497(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate1498(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );

  xor2  gate1429(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate1430(.a(gate112inter0), .b(s_126), .O(gate112inter1));
  and2  gate1431(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate1432(.a(s_126), .O(gate112inter3));
  inv1  gate1433(.a(s_127), .O(gate112inter4));
  nand2 gate1434(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate1435(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate1436(.a(G376), .O(gate112inter7));
  inv1  gate1437(.a(G377), .O(gate112inter8));
  nand2 gate1438(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate1439(.a(s_127), .b(gate112inter3), .O(gate112inter10));
  nor2  gate1440(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate1441(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate1442(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );

  xor2  gate1149(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate1150(.a(gate114inter0), .b(s_86), .O(gate114inter1));
  and2  gate1151(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate1152(.a(s_86), .O(gate114inter3));
  inv1  gate1153(.a(s_87), .O(gate114inter4));
  nand2 gate1154(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate1155(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate1156(.a(G380), .O(gate114inter7));
  inv1  gate1157(.a(G381), .O(gate114inter8));
  nand2 gate1158(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate1159(.a(s_87), .b(gate114inter3), .O(gate114inter10));
  nor2  gate1160(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate1161(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate1162(.a(gate114inter12), .b(gate114inter1), .O(G453));

  xor2  gate1569(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate1570(.a(gate115inter0), .b(s_146), .O(gate115inter1));
  and2  gate1571(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate1572(.a(s_146), .O(gate115inter3));
  inv1  gate1573(.a(s_147), .O(gate115inter4));
  nand2 gate1574(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate1575(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate1576(.a(G382), .O(gate115inter7));
  inv1  gate1577(.a(G383), .O(gate115inter8));
  nand2 gate1578(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate1579(.a(s_147), .b(gate115inter3), .O(gate115inter10));
  nor2  gate1580(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate1581(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate1582(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );

  xor2  gate2073(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate2074(.a(gate122inter0), .b(s_218), .O(gate122inter1));
  and2  gate2075(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate2076(.a(s_218), .O(gate122inter3));
  inv1  gate2077(.a(s_219), .O(gate122inter4));
  nand2 gate2078(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate2079(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate2080(.a(G396), .O(gate122inter7));
  inv1  gate2081(.a(G397), .O(gate122inter8));
  nand2 gate2082(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate2083(.a(s_219), .b(gate122inter3), .O(gate122inter10));
  nor2  gate2084(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate2085(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate2086(.a(gate122inter12), .b(gate122inter1), .O(G477));
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );

  xor2  gate673(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate674(.a(gate127inter0), .b(s_18), .O(gate127inter1));
  and2  gate675(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate676(.a(s_18), .O(gate127inter3));
  inv1  gate677(.a(s_19), .O(gate127inter4));
  nand2 gate678(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate679(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate680(.a(G406), .O(gate127inter7));
  inv1  gate681(.a(G407), .O(gate127inter8));
  nand2 gate682(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate683(.a(s_19), .b(gate127inter3), .O(gate127inter10));
  nor2  gate684(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate685(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate686(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate1793(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate1794(.a(gate132inter0), .b(s_178), .O(gate132inter1));
  and2  gate1795(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate1796(.a(s_178), .O(gate132inter3));
  inv1  gate1797(.a(s_179), .O(gate132inter4));
  nand2 gate1798(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate1799(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate1800(.a(G416), .O(gate132inter7));
  inv1  gate1801(.a(G417), .O(gate132inter8));
  nand2 gate1802(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate1803(.a(s_179), .b(gate132inter3), .O(gate132inter10));
  nor2  gate1804(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate1805(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate1806(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );

  xor2  gate1261(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate1262(.a(gate139inter0), .b(s_102), .O(gate139inter1));
  and2  gate1263(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate1264(.a(s_102), .O(gate139inter3));
  inv1  gate1265(.a(s_103), .O(gate139inter4));
  nand2 gate1266(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate1267(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate1268(.a(G438), .O(gate139inter7));
  inv1  gate1269(.a(G441), .O(gate139inter8));
  nand2 gate1270(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate1271(.a(s_103), .b(gate139inter3), .O(gate139inter10));
  nor2  gate1272(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate1273(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate1274(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );

  xor2  gate1513(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate1514(.a(gate145inter0), .b(s_138), .O(gate145inter1));
  and2  gate1515(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate1516(.a(s_138), .O(gate145inter3));
  inv1  gate1517(.a(s_139), .O(gate145inter4));
  nand2 gate1518(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate1519(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate1520(.a(G474), .O(gate145inter7));
  inv1  gate1521(.a(G477), .O(gate145inter8));
  nand2 gate1522(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate1523(.a(s_139), .b(gate145inter3), .O(gate145inter10));
  nor2  gate1524(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate1525(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate1526(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate2101(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate2102(.a(gate157inter0), .b(s_222), .O(gate157inter1));
  and2  gate2103(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate2104(.a(s_222), .O(gate157inter3));
  inv1  gate2105(.a(s_223), .O(gate157inter4));
  nand2 gate2106(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate2107(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate2108(.a(G438), .O(gate157inter7));
  inv1  gate2109(.a(G528), .O(gate157inter8));
  nand2 gate2110(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate2111(.a(s_223), .b(gate157inter3), .O(gate157inter10));
  nor2  gate2112(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate2113(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate2114(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate729(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate730(.a(gate159inter0), .b(s_26), .O(gate159inter1));
  and2  gate731(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate732(.a(s_26), .O(gate159inter3));
  inv1  gate733(.a(s_27), .O(gate159inter4));
  nand2 gate734(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate735(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate736(.a(G444), .O(gate159inter7));
  inv1  gate737(.a(G531), .O(gate159inter8));
  nand2 gate738(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate739(.a(s_27), .b(gate159inter3), .O(gate159inter10));
  nor2  gate740(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate741(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate742(.a(gate159inter12), .b(gate159inter1), .O(G576));

  xor2  gate1905(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate1906(.a(gate160inter0), .b(s_194), .O(gate160inter1));
  and2  gate1907(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate1908(.a(s_194), .O(gate160inter3));
  inv1  gate1909(.a(s_195), .O(gate160inter4));
  nand2 gate1910(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate1911(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate1912(.a(G447), .O(gate160inter7));
  inv1  gate1913(.a(G531), .O(gate160inter8));
  nand2 gate1914(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate1915(.a(s_195), .b(gate160inter3), .O(gate160inter10));
  nor2  gate1916(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate1917(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate1918(.a(gate160inter12), .b(gate160inter1), .O(G577));

  xor2  gate1919(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate1920(.a(gate161inter0), .b(s_196), .O(gate161inter1));
  and2  gate1921(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate1922(.a(s_196), .O(gate161inter3));
  inv1  gate1923(.a(s_197), .O(gate161inter4));
  nand2 gate1924(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate1925(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate1926(.a(G450), .O(gate161inter7));
  inv1  gate1927(.a(G534), .O(gate161inter8));
  nand2 gate1928(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate1929(.a(s_197), .b(gate161inter3), .O(gate161inter10));
  nor2  gate1930(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate1931(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate1932(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate1555(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate1556(.a(gate170inter0), .b(s_144), .O(gate170inter1));
  and2  gate1557(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate1558(.a(s_144), .O(gate170inter3));
  inv1  gate1559(.a(s_145), .O(gate170inter4));
  nand2 gate1560(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate1561(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate1562(.a(G477), .O(gate170inter7));
  inv1  gate1563(.a(G546), .O(gate170inter8));
  nand2 gate1564(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate1565(.a(s_145), .b(gate170inter3), .O(gate170inter10));
  nor2  gate1566(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate1567(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate1568(.a(gate170inter12), .b(gate170inter1), .O(G587));

  xor2  gate2185(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate2186(.a(gate171inter0), .b(s_234), .O(gate171inter1));
  and2  gate2187(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate2188(.a(s_234), .O(gate171inter3));
  inv1  gate2189(.a(s_235), .O(gate171inter4));
  nand2 gate2190(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate2191(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate2192(.a(G480), .O(gate171inter7));
  inv1  gate2193(.a(G549), .O(gate171inter8));
  nand2 gate2194(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate2195(.a(s_235), .b(gate171inter3), .O(gate171inter10));
  nor2  gate2196(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate2197(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate2198(.a(gate171inter12), .b(gate171inter1), .O(G588));
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate1345(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate1346(.a(gate175inter0), .b(s_114), .O(gate175inter1));
  and2  gate1347(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate1348(.a(s_114), .O(gate175inter3));
  inv1  gate1349(.a(s_115), .O(gate175inter4));
  nand2 gate1350(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1351(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1352(.a(G492), .O(gate175inter7));
  inv1  gate1353(.a(G555), .O(gate175inter8));
  nand2 gate1354(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1355(.a(s_115), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1356(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1357(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1358(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );

  xor2  gate1331(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate1332(.a(gate177inter0), .b(s_112), .O(gate177inter1));
  and2  gate1333(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate1334(.a(s_112), .O(gate177inter3));
  inv1  gate1335(.a(s_113), .O(gate177inter4));
  nand2 gate1336(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate1337(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate1338(.a(G498), .O(gate177inter7));
  inv1  gate1339(.a(G558), .O(gate177inter8));
  nand2 gate1340(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate1341(.a(s_113), .b(gate177inter3), .O(gate177inter10));
  nor2  gate1342(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate1343(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate1344(.a(gate177inter12), .b(gate177inter1), .O(G594));
nand2 gate178( .a(G501), .b(G558), .O(G595) );

  xor2  gate561(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate562(.a(gate179inter0), .b(s_2), .O(gate179inter1));
  and2  gate563(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate564(.a(s_2), .O(gate179inter3));
  inv1  gate565(.a(s_3), .O(gate179inter4));
  nand2 gate566(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate567(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate568(.a(G504), .O(gate179inter7));
  inv1  gate569(.a(G561), .O(gate179inter8));
  nand2 gate570(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate571(.a(s_3), .b(gate179inter3), .O(gate179inter10));
  nor2  gate572(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate573(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate574(.a(gate179inter12), .b(gate179inter1), .O(G596));
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate1079(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate1080(.a(gate191inter0), .b(s_76), .O(gate191inter1));
  and2  gate1081(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate1082(.a(s_76), .O(gate191inter3));
  inv1  gate1083(.a(s_77), .O(gate191inter4));
  nand2 gate1084(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate1085(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate1086(.a(G582), .O(gate191inter7));
  inv1  gate1087(.a(G583), .O(gate191inter8));
  nand2 gate1088(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate1089(.a(s_77), .b(gate191inter3), .O(gate191inter10));
  nor2  gate1090(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate1091(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate1092(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate617(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate618(.a(gate196inter0), .b(s_10), .O(gate196inter1));
  and2  gate619(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate620(.a(s_10), .O(gate196inter3));
  inv1  gate621(.a(s_11), .O(gate196inter4));
  nand2 gate622(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate623(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate624(.a(G592), .O(gate196inter7));
  inv1  gate625(.a(G593), .O(gate196inter8));
  nand2 gate626(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate627(.a(s_11), .b(gate196inter3), .O(gate196inter10));
  nor2  gate628(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate629(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate630(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate2129(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate2130(.a(gate200inter0), .b(s_226), .O(gate200inter1));
  and2  gate2131(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate2132(.a(s_226), .O(gate200inter3));
  inv1  gate2133(.a(s_227), .O(gate200inter4));
  nand2 gate2134(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate2135(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate2136(.a(G600), .O(gate200inter7));
  inv1  gate2137(.a(G601), .O(gate200inter8));
  nand2 gate2138(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate2139(.a(s_227), .b(gate200inter3), .O(gate200inter10));
  nor2  gate2140(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate2141(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate2142(.a(gate200inter12), .b(gate200inter1), .O(G663));
nand2 gate201( .a(G602), .b(G607), .O(G666) );

  xor2  gate1471(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate1472(.a(gate202inter0), .b(s_132), .O(gate202inter1));
  and2  gate1473(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate1474(.a(s_132), .O(gate202inter3));
  inv1  gate1475(.a(s_133), .O(gate202inter4));
  nand2 gate1476(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate1477(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate1478(.a(G612), .O(gate202inter7));
  inv1  gate1479(.a(G617), .O(gate202inter8));
  nand2 gate1480(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate1481(.a(s_133), .b(gate202inter3), .O(gate202inter10));
  nor2  gate1482(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate1483(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate1484(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );

  xor2  gate715(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate716(.a(gate207inter0), .b(s_24), .O(gate207inter1));
  and2  gate717(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate718(.a(s_24), .O(gate207inter3));
  inv1  gate719(.a(s_25), .O(gate207inter4));
  nand2 gate720(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate721(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate722(.a(G622), .O(gate207inter7));
  inv1  gate723(.a(G632), .O(gate207inter8));
  nand2 gate724(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate725(.a(s_25), .b(gate207inter3), .O(gate207inter10));
  nor2  gate726(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate727(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate728(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );

  xor2  gate1751(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate1752(.a(gate212inter0), .b(s_172), .O(gate212inter1));
  and2  gate1753(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate1754(.a(s_172), .O(gate212inter3));
  inv1  gate1755(.a(s_173), .O(gate212inter4));
  nand2 gate1756(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate1757(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate1758(.a(G617), .O(gate212inter7));
  inv1  gate1759(.a(G669), .O(gate212inter8));
  nand2 gate1760(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate1761(.a(s_173), .b(gate212inter3), .O(gate212inter10));
  nor2  gate1762(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate1763(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate1764(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate1317(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate1318(.a(gate215inter0), .b(s_110), .O(gate215inter1));
  and2  gate1319(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate1320(.a(s_110), .O(gate215inter3));
  inv1  gate1321(.a(s_111), .O(gate215inter4));
  nand2 gate1322(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate1323(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate1324(.a(G607), .O(gate215inter7));
  inv1  gate1325(.a(G675), .O(gate215inter8));
  nand2 gate1326(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate1327(.a(s_111), .b(gate215inter3), .O(gate215inter10));
  nor2  gate1328(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate1329(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate1330(.a(gate215inter12), .b(gate215inter1), .O(G696));

  xor2  gate1625(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate1626(.a(gate216inter0), .b(s_154), .O(gate216inter1));
  and2  gate1627(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate1628(.a(s_154), .O(gate216inter3));
  inv1  gate1629(.a(s_155), .O(gate216inter4));
  nand2 gate1630(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate1631(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate1632(.a(G617), .O(gate216inter7));
  inv1  gate1633(.a(G675), .O(gate216inter8));
  nand2 gate1634(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate1635(.a(s_155), .b(gate216inter3), .O(gate216inter10));
  nor2  gate1636(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate1637(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate1638(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate1695(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate1696(.a(gate220inter0), .b(s_164), .O(gate220inter1));
  and2  gate1697(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate1698(.a(s_164), .O(gate220inter3));
  inv1  gate1699(.a(s_165), .O(gate220inter4));
  nand2 gate1700(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate1701(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate1702(.a(G637), .O(gate220inter7));
  inv1  gate1703(.a(G681), .O(gate220inter8));
  nand2 gate1704(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate1705(.a(s_165), .b(gate220inter3), .O(gate220inter10));
  nor2  gate1706(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate1707(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate1708(.a(gate220inter12), .b(gate220inter1), .O(G701));
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate827(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate828(.a(gate223inter0), .b(s_40), .O(gate223inter1));
  and2  gate829(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate830(.a(s_40), .O(gate223inter3));
  inv1  gate831(.a(s_41), .O(gate223inter4));
  nand2 gate832(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate833(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate834(.a(G627), .O(gate223inter7));
  inv1  gate835(.a(G687), .O(gate223inter8));
  nand2 gate836(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate837(.a(s_41), .b(gate223inter3), .O(gate223inter10));
  nor2  gate838(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate839(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate840(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );

  xor2  gate1821(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate1822(.a(gate225inter0), .b(s_182), .O(gate225inter1));
  and2  gate1823(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate1824(.a(s_182), .O(gate225inter3));
  inv1  gate1825(.a(s_183), .O(gate225inter4));
  nand2 gate1826(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate1827(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate1828(.a(G690), .O(gate225inter7));
  inv1  gate1829(.a(G691), .O(gate225inter8));
  nand2 gate1830(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate1831(.a(s_183), .b(gate225inter3), .O(gate225inter10));
  nor2  gate1832(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate1833(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate1834(.a(gate225inter12), .b(gate225inter1), .O(G706));
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate589(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate590(.a(gate228inter0), .b(s_6), .O(gate228inter1));
  and2  gate591(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate592(.a(s_6), .O(gate228inter3));
  inv1  gate593(.a(s_7), .O(gate228inter4));
  nand2 gate594(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate595(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate596(.a(G696), .O(gate228inter7));
  inv1  gate597(.a(G697), .O(gate228inter8));
  nand2 gate598(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate599(.a(s_7), .b(gate228inter3), .O(gate228inter10));
  nor2  gate600(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate601(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate602(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate1597(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate1598(.a(gate233inter0), .b(s_150), .O(gate233inter1));
  and2  gate1599(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate1600(.a(s_150), .O(gate233inter3));
  inv1  gate1601(.a(s_151), .O(gate233inter4));
  nand2 gate1602(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1603(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1604(.a(G242), .O(gate233inter7));
  inv1  gate1605(.a(G718), .O(gate233inter8));
  nand2 gate1606(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1607(.a(s_151), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1608(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1609(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1610(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );

  xor2  gate1863(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate1864(.a(gate239inter0), .b(s_188), .O(gate239inter1));
  and2  gate1865(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate1866(.a(s_188), .O(gate239inter3));
  inv1  gate1867(.a(s_189), .O(gate239inter4));
  nand2 gate1868(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate1869(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate1870(.a(G260), .O(gate239inter7));
  inv1  gate1871(.a(G712), .O(gate239inter8));
  nand2 gate1872(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate1873(.a(s_189), .b(gate239inter3), .O(gate239inter10));
  nor2  gate1874(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate1875(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate1876(.a(gate239inter12), .b(gate239inter1), .O(G748));
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate1065(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate1066(.a(gate241inter0), .b(s_74), .O(gate241inter1));
  and2  gate1067(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate1068(.a(s_74), .O(gate241inter3));
  inv1  gate1069(.a(s_75), .O(gate241inter4));
  nand2 gate1070(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate1071(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate1072(.a(G242), .O(gate241inter7));
  inv1  gate1073(.a(G730), .O(gate241inter8));
  nand2 gate1074(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate1075(.a(s_75), .b(gate241inter3), .O(gate241inter10));
  nor2  gate1076(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate1077(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate1078(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate1639(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1640(.a(gate243inter0), .b(s_156), .O(gate243inter1));
  and2  gate1641(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1642(.a(s_156), .O(gate243inter3));
  inv1  gate1643(.a(s_157), .O(gate243inter4));
  nand2 gate1644(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1645(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1646(.a(G245), .O(gate243inter7));
  inv1  gate1647(.a(G733), .O(gate243inter8));
  nand2 gate1648(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1649(.a(s_157), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1650(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1651(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1652(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );

  xor2  gate1765(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate1766(.a(gate248inter0), .b(s_174), .O(gate248inter1));
  and2  gate1767(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate1768(.a(s_174), .O(gate248inter3));
  inv1  gate1769(.a(s_175), .O(gate248inter4));
  nand2 gate1770(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate1771(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate1772(.a(G727), .O(gate248inter7));
  inv1  gate1773(.a(G739), .O(gate248inter8));
  nand2 gate1774(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate1775(.a(s_175), .b(gate248inter3), .O(gate248inter10));
  nor2  gate1776(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate1777(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate1778(.a(gate248inter12), .b(gate248inter1), .O(G761));

  xor2  gate953(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate954(.a(gate249inter0), .b(s_58), .O(gate249inter1));
  and2  gate955(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate956(.a(s_58), .O(gate249inter3));
  inv1  gate957(.a(s_59), .O(gate249inter4));
  nand2 gate958(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate959(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate960(.a(G254), .O(gate249inter7));
  inv1  gate961(.a(G742), .O(gate249inter8));
  nand2 gate962(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate963(.a(s_59), .b(gate249inter3), .O(gate249inter10));
  nor2  gate964(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate965(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate966(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );

  xor2  gate995(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate996(.a(gate251inter0), .b(s_64), .O(gate251inter1));
  and2  gate997(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate998(.a(s_64), .O(gate251inter3));
  inv1  gate999(.a(s_65), .O(gate251inter4));
  nand2 gate1000(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate1001(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate1002(.a(G257), .O(gate251inter7));
  inv1  gate1003(.a(G745), .O(gate251inter8));
  nand2 gate1004(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate1005(.a(s_65), .b(gate251inter3), .O(gate251inter10));
  nor2  gate1006(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate1007(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate1008(.a(gate251inter12), .b(gate251inter1), .O(G764));
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );

  xor2  gate1387(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate1388(.a(gate259inter0), .b(s_120), .O(gate259inter1));
  and2  gate1389(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate1390(.a(s_120), .O(gate259inter3));
  inv1  gate1391(.a(s_121), .O(gate259inter4));
  nand2 gate1392(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate1393(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate1394(.a(G758), .O(gate259inter7));
  inv1  gate1395(.a(G759), .O(gate259inter8));
  nand2 gate1396(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate1397(.a(s_121), .b(gate259inter3), .O(gate259inter10));
  nor2  gate1398(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate1399(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate1400(.a(gate259inter12), .b(gate259inter1), .O(G776));

  xor2  gate1233(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate1234(.a(gate260inter0), .b(s_98), .O(gate260inter1));
  and2  gate1235(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate1236(.a(s_98), .O(gate260inter3));
  inv1  gate1237(.a(s_99), .O(gate260inter4));
  nand2 gate1238(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate1239(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate1240(.a(G760), .O(gate260inter7));
  inv1  gate1241(.a(G761), .O(gate260inter8));
  nand2 gate1242(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate1243(.a(s_99), .b(gate260inter3), .O(gate260inter10));
  nor2  gate1244(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate1245(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate1246(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate1947(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate1948(.a(gate262inter0), .b(s_200), .O(gate262inter1));
  and2  gate1949(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate1950(.a(s_200), .O(gate262inter3));
  inv1  gate1951(.a(s_201), .O(gate262inter4));
  nand2 gate1952(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate1953(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate1954(.a(G764), .O(gate262inter7));
  inv1  gate1955(.a(G765), .O(gate262inter8));
  nand2 gate1956(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate1957(.a(s_201), .b(gate262inter3), .O(gate262inter10));
  nor2  gate1958(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate1959(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate1960(.a(gate262inter12), .b(gate262inter1), .O(G785));

  xor2  gate659(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate660(.a(gate263inter0), .b(s_16), .O(gate263inter1));
  and2  gate661(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate662(.a(s_16), .O(gate263inter3));
  inv1  gate663(.a(s_17), .O(gate263inter4));
  nand2 gate664(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate665(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate666(.a(G766), .O(gate263inter7));
  inv1  gate667(.a(G767), .O(gate263inter8));
  nand2 gate668(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate669(.a(s_17), .b(gate263inter3), .O(gate263inter10));
  nor2  gate670(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate671(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate672(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate1093(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate1094(.a(gate266inter0), .b(s_78), .O(gate266inter1));
  and2  gate1095(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate1096(.a(s_78), .O(gate266inter3));
  inv1  gate1097(.a(s_79), .O(gate266inter4));
  nand2 gate1098(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate1099(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate1100(.a(G645), .O(gate266inter7));
  inv1  gate1101(.a(G773), .O(gate266inter8));
  nand2 gate1102(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate1103(.a(s_79), .b(gate266inter3), .O(gate266inter10));
  nor2  gate1104(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate1105(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate1106(.a(gate266inter12), .b(gate266inter1), .O(G797));

  xor2  gate1135(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate1136(.a(gate267inter0), .b(s_84), .O(gate267inter1));
  and2  gate1137(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate1138(.a(s_84), .O(gate267inter3));
  inv1  gate1139(.a(s_85), .O(gate267inter4));
  nand2 gate1140(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate1141(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate1142(.a(G648), .O(gate267inter7));
  inv1  gate1143(.a(G776), .O(gate267inter8));
  nand2 gate1144(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate1145(.a(s_85), .b(gate267inter3), .O(gate267inter10));
  nor2  gate1146(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate1147(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate1148(.a(gate267inter12), .b(gate267inter1), .O(G800));

  xor2  gate1527(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate1528(.a(gate268inter0), .b(s_140), .O(gate268inter1));
  and2  gate1529(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate1530(.a(s_140), .O(gate268inter3));
  inv1  gate1531(.a(s_141), .O(gate268inter4));
  nand2 gate1532(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1533(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1534(.a(G651), .O(gate268inter7));
  inv1  gate1535(.a(G779), .O(gate268inter8));
  nand2 gate1536(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1537(.a(s_141), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1538(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1539(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1540(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate743(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate744(.a(gate272inter0), .b(s_28), .O(gate272inter1));
  and2  gate745(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate746(.a(s_28), .O(gate272inter3));
  inv1  gate747(.a(s_29), .O(gate272inter4));
  nand2 gate748(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate749(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate750(.a(G663), .O(gate272inter7));
  inv1  gate751(.a(G791), .O(gate272inter8));
  nand2 gate752(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate753(.a(s_29), .b(gate272inter3), .O(gate272inter10));
  nor2  gate754(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate755(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate756(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate1107(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate1108(.a(gate274inter0), .b(s_80), .O(gate274inter1));
  and2  gate1109(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate1110(.a(s_80), .O(gate274inter3));
  inv1  gate1111(.a(s_81), .O(gate274inter4));
  nand2 gate1112(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate1113(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate1114(.a(G770), .O(gate274inter7));
  inv1  gate1115(.a(G794), .O(gate274inter8));
  nand2 gate1116(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate1117(.a(s_81), .b(gate274inter3), .O(gate274inter10));
  nor2  gate1118(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate1119(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate1120(.a(gate274inter12), .b(gate274inter1), .O(G819));

  xor2  gate575(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate576(.a(gate275inter0), .b(s_4), .O(gate275inter1));
  and2  gate577(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate578(.a(s_4), .O(gate275inter3));
  inv1  gate579(.a(s_5), .O(gate275inter4));
  nand2 gate580(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate581(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate582(.a(G645), .O(gate275inter7));
  inv1  gate583(.a(G797), .O(gate275inter8));
  nand2 gate584(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate585(.a(s_5), .b(gate275inter3), .O(gate275inter10));
  nor2  gate586(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate587(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate588(.a(gate275inter12), .b(gate275inter1), .O(G820));
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate2227(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate2228(.a(gate278inter0), .b(s_240), .O(gate278inter1));
  and2  gate2229(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate2230(.a(s_240), .O(gate278inter3));
  inv1  gate2231(.a(s_241), .O(gate278inter4));
  nand2 gate2232(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate2233(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate2234(.a(G776), .O(gate278inter7));
  inv1  gate2235(.a(G800), .O(gate278inter8));
  nand2 gate2236(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate2237(.a(s_241), .b(gate278inter3), .O(gate278inter10));
  nor2  gate2238(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate2239(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate2240(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate1457(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate1458(.a(gate293inter0), .b(s_130), .O(gate293inter1));
  and2  gate1459(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate1460(.a(s_130), .O(gate293inter3));
  inv1  gate1461(.a(s_131), .O(gate293inter4));
  nand2 gate1462(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate1463(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate1464(.a(G828), .O(gate293inter7));
  inv1  gate1465(.a(G829), .O(gate293inter8));
  nand2 gate1466(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate1467(.a(s_131), .b(gate293inter3), .O(gate293inter10));
  nor2  gate1468(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate1469(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate1470(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate645(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate646(.a(gate388inter0), .b(s_14), .O(gate388inter1));
  and2  gate647(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate648(.a(s_14), .O(gate388inter3));
  inv1  gate649(.a(s_15), .O(gate388inter4));
  nand2 gate650(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate651(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate652(.a(G2), .O(gate388inter7));
  inv1  gate653(.a(G1039), .O(gate388inter8));
  nand2 gate654(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate655(.a(s_15), .b(gate388inter3), .O(gate388inter10));
  nor2  gate656(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate657(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate658(.a(gate388inter12), .b(gate388inter1), .O(G1135));

  xor2  gate1275(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate1276(.a(gate389inter0), .b(s_104), .O(gate389inter1));
  and2  gate1277(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate1278(.a(s_104), .O(gate389inter3));
  inv1  gate1279(.a(s_105), .O(gate389inter4));
  nand2 gate1280(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate1281(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate1282(.a(G3), .O(gate389inter7));
  inv1  gate1283(.a(G1042), .O(gate389inter8));
  nand2 gate1284(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate1285(.a(s_105), .b(gate389inter3), .O(gate389inter10));
  nor2  gate1286(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate1287(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate1288(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );

  xor2  gate1583(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate1584(.a(gate392inter0), .b(s_148), .O(gate392inter1));
  and2  gate1585(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate1586(.a(s_148), .O(gate392inter3));
  inv1  gate1587(.a(s_149), .O(gate392inter4));
  nand2 gate1588(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate1589(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate1590(.a(G6), .O(gate392inter7));
  inv1  gate1591(.a(G1051), .O(gate392inter8));
  nand2 gate1592(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate1593(.a(s_149), .b(gate392inter3), .O(gate392inter10));
  nor2  gate1594(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate1595(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate1596(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate1023(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate1024(.a(gate394inter0), .b(s_68), .O(gate394inter1));
  and2  gate1025(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate1026(.a(s_68), .O(gate394inter3));
  inv1  gate1027(.a(s_69), .O(gate394inter4));
  nand2 gate1028(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate1029(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate1030(.a(G8), .O(gate394inter7));
  inv1  gate1031(.a(G1057), .O(gate394inter8));
  nand2 gate1032(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate1033(.a(s_69), .b(gate394inter3), .O(gate394inter10));
  nor2  gate1034(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate1035(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate1036(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );

  xor2  gate2017(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate2018(.a(gate401inter0), .b(s_210), .O(gate401inter1));
  and2  gate2019(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate2020(.a(s_210), .O(gate401inter3));
  inv1  gate2021(.a(s_211), .O(gate401inter4));
  nand2 gate2022(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate2023(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate2024(.a(G15), .O(gate401inter7));
  inv1  gate2025(.a(G1078), .O(gate401inter8));
  nand2 gate2026(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate2027(.a(s_211), .b(gate401inter3), .O(gate401inter10));
  nor2  gate2028(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate2029(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate2030(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );

  xor2  gate1933(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate1934(.a(gate408inter0), .b(s_198), .O(gate408inter1));
  and2  gate1935(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate1936(.a(s_198), .O(gate408inter3));
  inv1  gate1937(.a(s_199), .O(gate408inter4));
  nand2 gate1938(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate1939(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate1940(.a(G22), .O(gate408inter7));
  inv1  gate1941(.a(G1099), .O(gate408inter8));
  nand2 gate1942(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate1943(.a(s_199), .b(gate408inter3), .O(gate408inter10));
  nor2  gate1944(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate1945(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate1946(.a(gate408inter12), .b(gate408inter1), .O(G1195));
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate1681(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate1682(.a(gate413inter0), .b(s_162), .O(gate413inter1));
  and2  gate1683(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate1684(.a(s_162), .O(gate413inter3));
  inv1  gate1685(.a(s_163), .O(gate413inter4));
  nand2 gate1686(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1687(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1688(.a(G27), .O(gate413inter7));
  inv1  gate1689(.a(G1114), .O(gate413inter8));
  nand2 gate1690(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1691(.a(s_163), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1692(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1693(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1694(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate2031(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate2032(.a(gate415inter0), .b(s_212), .O(gate415inter1));
  and2  gate2033(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate2034(.a(s_212), .O(gate415inter3));
  inv1  gate2035(.a(s_213), .O(gate415inter4));
  nand2 gate2036(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate2037(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate2038(.a(G29), .O(gate415inter7));
  inv1  gate2039(.a(G1120), .O(gate415inter8));
  nand2 gate2040(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate2041(.a(s_213), .b(gate415inter3), .O(gate415inter10));
  nor2  gate2042(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate2043(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate2044(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate1541(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate1542(.a(gate417inter0), .b(s_142), .O(gate417inter1));
  and2  gate1543(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate1544(.a(s_142), .O(gate417inter3));
  inv1  gate1545(.a(s_143), .O(gate417inter4));
  nand2 gate1546(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate1547(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate1548(.a(G31), .O(gate417inter7));
  inv1  gate1549(.a(G1126), .O(gate417inter8));
  nand2 gate1550(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate1551(.a(s_143), .b(gate417inter3), .O(gate417inter10));
  nor2  gate1552(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate1553(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate1554(.a(gate417inter12), .b(gate417inter1), .O(G1222));
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate1835(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate1836(.a(gate425inter0), .b(s_184), .O(gate425inter1));
  and2  gate1837(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate1838(.a(s_184), .O(gate425inter3));
  inv1  gate1839(.a(s_185), .O(gate425inter4));
  nand2 gate1840(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1841(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1842(.a(G4), .O(gate425inter7));
  inv1  gate1843(.a(G1141), .O(gate425inter8));
  nand2 gate1844(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1845(.a(s_185), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1846(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1847(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1848(.a(gate425inter12), .b(gate425inter1), .O(G1234));
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate1611(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate1612(.a(gate430inter0), .b(s_152), .O(gate430inter1));
  and2  gate1613(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate1614(.a(s_152), .O(gate430inter3));
  inv1  gate1615(.a(s_153), .O(gate430inter4));
  nand2 gate1616(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate1617(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate1618(.a(G1051), .O(gate430inter7));
  inv1  gate1619(.a(G1147), .O(gate430inter8));
  nand2 gate1620(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate1621(.a(s_153), .b(gate430inter3), .O(gate430inter10));
  nor2  gate1622(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate1623(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate1624(.a(gate430inter12), .b(gate430inter1), .O(G1239));

  xor2  gate2003(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate2004(.a(gate431inter0), .b(s_208), .O(gate431inter1));
  and2  gate2005(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate2006(.a(s_208), .O(gate431inter3));
  inv1  gate2007(.a(s_209), .O(gate431inter4));
  nand2 gate2008(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate2009(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate2010(.a(G7), .O(gate431inter7));
  inv1  gate2011(.a(G1150), .O(gate431inter8));
  nand2 gate2012(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate2013(.a(s_209), .b(gate431inter3), .O(gate431inter10));
  nor2  gate2014(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate2015(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate2016(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate897(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate898(.a(gate434inter0), .b(s_50), .O(gate434inter1));
  and2  gate899(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate900(.a(s_50), .O(gate434inter3));
  inv1  gate901(.a(s_51), .O(gate434inter4));
  nand2 gate902(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate903(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate904(.a(G1057), .O(gate434inter7));
  inv1  gate905(.a(G1153), .O(gate434inter8));
  nand2 gate906(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate907(.a(s_51), .b(gate434inter3), .O(gate434inter10));
  nor2  gate908(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate909(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate910(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );

  xor2  gate547(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate548(.a(gate436inter0), .b(s_0), .O(gate436inter1));
  and2  gate549(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate550(.a(s_0), .O(gate436inter3));
  inv1  gate551(.a(s_1), .O(gate436inter4));
  nand2 gate552(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate553(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate554(.a(G1060), .O(gate436inter7));
  inv1  gate555(.a(G1156), .O(gate436inter8));
  nand2 gate556(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate557(.a(s_1), .b(gate436inter3), .O(gate436inter10));
  nor2  gate558(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate559(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate560(.a(gate436inter12), .b(gate436inter1), .O(G1245));

  xor2  gate883(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate884(.a(gate437inter0), .b(s_48), .O(gate437inter1));
  and2  gate885(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate886(.a(s_48), .O(gate437inter3));
  inv1  gate887(.a(s_49), .O(gate437inter4));
  nand2 gate888(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate889(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate890(.a(G10), .O(gate437inter7));
  inv1  gate891(.a(G1159), .O(gate437inter8));
  nand2 gate892(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate893(.a(s_49), .b(gate437inter3), .O(gate437inter10));
  nor2  gate894(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate895(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate896(.a(gate437inter12), .b(gate437inter1), .O(G1246));
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate2143(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate2144(.a(gate443inter0), .b(s_228), .O(gate443inter1));
  and2  gate2145(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate2146(.a(s_228), .O(gate443inter3));
  inv1  gate2147(.a(s_229), .O(gate443inter4));
  nand2 gate2148(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate2149(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate2150(.a(G13), .O(gate443inter7));
  inv1  gate2151(.a(G1168), .O(gate443inter8));
  nand2 gate2152(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate2153(.a(s_229), .b(gate443inter3), .O(gate443inter10));
  nor2  gate2154(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate2155(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate2156(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate1121(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate1122(.a(gate445inter0), .b(s_82), .O(gate445inter1));
  and2  gate1123(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate1124(.a(s_82), .O(gate445inter3));
  inv1  gate1125(.a(s_83), .O(gate445inter4));
  nand2 gate1126(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate1127(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate1128(.a(G14), .O(gate445inter7));
  inv1  gate1129(.a(G1171), .O(gate445inter8));
  nand2 gate1130(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate1131(.a(s_83), .b(gate445inter3), .O(gate445inter10));
  nor2  gate1132(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate1133(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate1134(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate1177(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate1178(.a(gate448inter0), .b(s_90), .O(gate448inter1));
  and2  gate1179(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate1180(.a(s_90), .O(gate448inter3));
  inv1  gate1181(.a(s_91), .O(gate448inter4));
  nand2 gate1182(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate1183(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate1184(.a(G1078), .O(gate448inter7));
  inv1  gate1185(.a(G1174), .O(gate448inter8));
  nand2 gate1186(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate1187(.a(s_91), .b(gate448inter3), .O(gate448inter10));
  nor2  gate1188(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate1189(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate1190(.a(gate448inter12), .b(gate448inter1), .O(G1257));
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );

  xor2  gate1373(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate1374(.a(gate452inter0), .b(s_118), .O(gate452inter1));
  and2  gate1375(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate1376(.a(s_118), .O(gate452inter3));
  inv1  gate1377(.a(s_119), .O(gate452inter4));
  nand2 gate1378(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate1379(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate1380(.a(G1084), .O(gate452inter7));
  inv1  gate1381(.a(G1180), .O(gate452inter8));
  nand2 gate1382(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate1383(.a(s_119), .b(gate452inter3), .O(gate452inter10));
  nor2  gate1384(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate1385(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate1386(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );

  xor2  gate1989(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate1990(.a(gate455inter0), .b(s_206), .O(gate455inter1));
  and2  gate1991(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate1992(.a(s_206), .O(gate455inter3));
  inv1  gate1993(.a(s_207), .O(gate455inter4));
  nand2 gate1994(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate1995(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate1996(.a(G19), .O(gate455inter7));
  inv1  gate1997(.a(G1186), .O(gate455inter8));
  nand2 gate1998(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate1999(.a(s_207), .b(gate455inter3), .O(gate455inter10));
  nor2  gate2000(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate2001(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate2002(.a(gate455inter12), .b(gate455inter1), .O(G1264));

  xor2  gate785(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate786(.a(gate456inter0), .b(s_34), .O(gate456inter1));
  and2  gate787(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate788(.a(s_34), .O(gate456inter3));
  inv1  gate789(.a(s_35), .O(gate456inter4));
  nand2 gate790(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate791(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate792(.a(G1090), .O(gate456inter7));
  inv1  gate793(.a(G1186), .O(gate456inter8));
  nand2 gate794(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate795(.a(s_35), .b(gate456inter3), .O(gate456inter10));
  nor2  gate796(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate797(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate798(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );

  xor2  gate2171(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate2172(.a(gate458inter0), .b(s_232), .O(gate458inter1));
  and2  gate2173(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate2174(.a(s_232), .O(gate458inter3));
  inv1  gate2175(.a(s_233), .O(gate458inter4));
  nand2 gate2176(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate2177(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate2178(.a(G1093), .O(gate458inter7));
  inv1  gate2179(.a(G1189), .O(gate458inter8));
  nand2 gate2180(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate2181(.a(s_233), .b(gate458inter3), .O(gate458inter10));
  nor2  gate2182(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate2183(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate2184(.a(gate458inter12), .b(gate458inter1), .O(G1267));
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate1653(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate1654(.a(gate463inter0), .b(s_158), .O(gate463inter1));
  and2  gate1655(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate1656(.a(s_158), .O(gate463inter3));
  inv1  gate1657(.a(s_159), .O(gate463inter4));
  nand2 gate1658(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate1659(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate1660(.a(G23), .O(gate463inter7));
  inv1  gate1661(.a(G1198), .O(gate463inter8));
  nand2 gate1662(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate1663(.a(s_159), .b(gate463inter3), .O(gate463inter10));
  nor2  gate1664(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate1665(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate1666(.a(gate463inter12), .b(gate463inter1), .O(G1272));

  xor2  gate981(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate982(.a(gate464inter0), .b(s_62), .O(gate464inter1));
  and2  gate983(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate984(.a(s_62), .O(gate464inter3));
  inv1  gate985(.a(s_63), .O(gate464inter4));
  nand2 gate986(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate987(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate988(.a(G1102), .O(gate464inter7));
  inv1  gate989(.a(G1198), .O(gate464inter8));
  nand2 gate990(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate991(.a(s_63), .b(gate464inter3), .O(gate464inter10));
  nor2  gate992(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate993(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate994(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate687(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate688(.a(gate466inter0), .b(s_20), .O(gate466inter1));
  and2  gate689(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate690(.a(s_20), .O(gate466inter3));
  inv1  gate691(.a(s_21), .O(gate466inter4));
  nand2 gate692(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate693(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate694(.a(G1105), .O(gate466inter7));
  inv1  gate695(.a(G1201), .O(gate466inter8));
  nand2 gate696(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate697(.a(s_21), .b(gate466inter3), .O(gate466inter10));
  nor2  gate698(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate699(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate700(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate1961(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate1962(.a(gate472inter0), .b(s_202), .O(gate472inter1));
  and2  gate1963(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate1964(.a(s_202), .O(gate472inter3));
  inv1  gate1965(.a(s_203), .O(gate472inter4));
  nand2 gate1966(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate1967(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate1968(.a(G1114), .O(gate472inter7));
  inv1  gate1969(.a(G1210), .O(gate472inter8));
  nand2 gate1970(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate1971(.a(s_203), .b(gate472inter3), .O(gate472inter10));
  nor2  gate1972(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate1973(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate1974(.a(gate472inter12), .b(gate472inter1), .O(G1281));

  xor2  gate813(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate814(.a(gate473inter0), .b(s_38), .O(gate473inter1));
  and2  gate815(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate816(.a(s_38), .O(gate473inter3));
  inv1  gate817(.a(s_39), .O(gate473inter4));
  nand2 gate818(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate819(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate820(.a(G28), .O(gate473inter7));
  inv1  gate821(.a(G1213), .O(gate473inter8));
  nand2 gate822(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate823(.a(s_39), .b(gate473inter3), .O(gate473inter10));
  nor2  gate824(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate825(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate826(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate1877(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate1878(.a(gate475inter0), .b(s_190), .O(gate475inter1));
  and2  gate1879(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate1880(.a(s_190), .O(gate475inter3));
  inv1  gate1881(.a(s_191), .O(gate475inter4));
  nand2 gate1882(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate1883(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate1884(.a(G29), .O(gate475inter7));
  inv1  gate1885(.a(G1216), .O(gate475inter8));
  nand2 gate1886(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate1887(.a(s_191), .b(gate475inter3), .O(gate475inter10));
  nor2  gate1888(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate1889(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate1890(.a(gate475inter12), .b(gate475inter1), .O(G1284));
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate1499(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate1500(.a(gate480inter0), .b(s_136), .O(gate480inter1));
  and2  gate1501(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate1502(.a(s_136), .O(gate480inter3));
  inv1  gate1503(.a(s_137), .O(gate480inter4));
  nand2 gate1504(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate1505(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate1506(.a(G1126), .O(gate480inter7));
  inv1  gate1507(.a(G1222), .O(gate480inter8));
  nand2 gate1508(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate1509(.a(s_137), .b(gate480inter3), .O(gate480inter10));
  nor2  gate1510(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate1511(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate1512(.a(gate480inter12), .b(gate480inter1), .O(G1289));

  xor2  gate2199(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate2200(.a(gate481inter0), .b(s_236), .O(gate481inter1));
  and2  gate2201(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate2202(.a(s_236), .O(gate481inter3));
  inv1  gate2203(.a(s_237), .O(gate481inter4));
  nand2 gate2204(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate2205(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate2206(.a(G32), .O(gate481inter7));
  inv1  gate2207(.a(G1225), .O(gate481inter8));
  nand2 gate2208(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate2209(.a(s_237), .b(gate481inter3), .O(gate481inter10));
  nor2  gate2210(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate2211(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate2212(.a(gate481inter12), .b(gate481inter1), .O(G1290));
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate1667(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate1668(.a(gate491inter0), .b(s_160), .O(gate491inter1));
  and2  gate1669(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate1670(.a(s_160), .O(gate491inter3));
  inv1  gate1671(.a(s_161), .O(gate491inter4));
  nand2 gate1672(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate1673(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate1674(.a(G1244), .O(gate491inter7));
  inv1  gate1675(.a(G1245), .O(gate491inter8));
  nand2 gate1676(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate1677(.a(s_161), .b(gate491inter3), .O(gate491inter10));
  nor2  gate1678(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate1679(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate1680(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate2213(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate2214(.a(gate493inter0), .b(s_238), .O(gate493inter1));
  and2  gate2215(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate2216(.a(s_238), .O(gate493inter3));
  inv1  gate2217(.a(s_239), .O(gate493inter4));
  nand2 gate2218(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate2219(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate2220(.a(G1248), .O(gate493inter7));
  inv1  gate2221(.a(G1249), .O(gate493inter8));
  nand2 gate2222(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate2223(.a(s_239), .b(gate493inter3), .O(gate493inter10));
  nor2  gate2224(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate2225(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate2226(.a(gate493inter12), .b(gate493inter1), .O(G1302));

  xor2  gate1891(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1892(.a(gate494inter0), .b(s_192), .O(gate494inter1));
  and2  gate1893(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1894(.a(s_192), .O(gate494inter3));
  inv1  gate1895(.a(s_193), .O(gate494inter4));
  nand2 gate1896(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1897(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1898(.a(G1250), .O(gate494inter7));
  inv1  gate1899(.a(G1251), .O(gate494inter8));
  nand2 gate1900(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1901(.a(s_193), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1902(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1903(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1904(.a(gate494inter12), .b(gate494inter1), .O(G1303));

  xor2  gate925(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate926(.a(gate495inter0), .b(s_54), .O(gate495inter1));
  and2  gate927(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate928(.a(s_54), .O(gate495inter3));
  inv1  gate929(.a(s_55), .O(gate495inter4));
  nand2 gate930(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate931(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate932(.a(G1252), .O(gate495inter7));
  inv1  gate933(.a(G1253), .O(gate495inter8));
  nand2 gate934(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate935(.a(s_55), .b(gate495inter3), .O(gate495inter10));
  nor2  gate936(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate937(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate938(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );

  xor2  gate1401(.a(G1257), .b(G1256), .O(gate497inter0));
  nand2 gate1402(.a(gate497inter0), .b(s_122), .O(gate497inter1));
  and2  gate1403(.a(G1257), .b(G1256), .O(gate497inter2));
  inv1  gate1404(.a(s_122), .O(gate497inter3));
  inv1  gate1405(.a(s_123), .O(gate497inter4));
  nand2 gate1406(.a(gate497inter4), .b(gate497inter3), .O(gate497inter5));
  nor2  gate1407(.a(gate497inter5), .b(gate497inter2), .O(gate497inter6));
  inv1  gate1408(.a(G1256), .O(gate497inter7));
  inv1  gate1409(.a(G1257), .O(gate497inter8));
  nand2 gate1410(.a(gate497inter8), .b(gate497inter7), .O(gate497inter9));
  nand2 gate1411(.a(s_123), .b(gate497inter3), .O(gate497inter10));
  nor2  gate1412(.a(gate497inter10), .b(gate497inter9), .O(gate497inter11));
  nor2  gate1413(.a(gate497inter11), .b(gate497inter6), .O(gate497inter12));
  nand2 gate1414(.a(gate497inter12), .b(gate497inter1), .O(G1306));
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate911(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate912(.a(gate500inter0), .b(s_52), .O(gate500inter1));
  and2  gate913(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate914(.a(s_52), .O(gate500inter3));
  inv1  gate915(.a(s_53), .O(gate500inter4));
  nand2 gate916(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate917(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate918(.a(G1262), .O(gate500inter7));
  inv1  gate919(.a(G1263), .O(gate500inter8));
  nand2 gate920(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate921(.a(s_53), .b(gate500inter3), .O(gate500inter10));
  nor2  gate922(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate923(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate924(.a(gate500inter12), .b(gate500inter1), .O(G1309));
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );

  xor2  gate1219(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate1220(.a(gate507inter0), .b(s_96), .O(gate507inter1));
  and2  gate1221(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate1222(.a(s_96), .O(gate507inter3));
  inv1  gate1223(.a(s_97), .O(gate507inter4));
  nand2 gate1224(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate1225(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate1226(.a(G1276), .O(gate507inter7));
  inv1  gate1227(.a(G1277), .O(gate507inter8));
  nand2 gate1228(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate1229(.a(s_97), .b(gate507inter3), .O(gate507inter10));
  nor2  gate1230(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate1231(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate1232(.a(gate507inter12), .b(gate507inter1), .O(G1316));
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule