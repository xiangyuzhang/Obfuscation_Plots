module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281, s_282, s_283, s_284, s_285, s_286, s_287, s_288, s_289, s_290, s_291, s_292, s_293, s_294, s_295, s_296, s_297, s_298, s_299, s_300, s_301, s_302, s_303, s_304, s_305, s_306, s_307, s_308, s_309, s_310, s_311, s_312, s_313, s_314, s_315, s_316, s_317, s_318, s_319, s_320, s_321, s_322, s_323, s_324, s_325, s_326, s_327, s_328, s_329, s_330, s_331, s_332, s_333, s_334, s_335, s_336, s_337, s_338, s_339, s_340, s_341, s_342, s_343, s_344, s_345, s_346, s_347, s_348, s_349, s_350, s_351;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate97inter0, gate97inter1, gate97inter2, gate97inter3, gate97inter4, gate97inter5, gate97inter6, gate97inter7, gate97inter8, gate97inter9, gate97inter10, gate97inter11, gate97inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate447inter0, gate447inter1, gate447inter2, gate447inter3, gate447inter4, gate447inter5, gate447inter6, gate447inter7, gate447inter8, gate447inter9, gate447inter10, gate447inter11, gate447inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate953(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate954(.a(gate17inter0), .b(s_58), .O(gate17inter1));
  and2  gate955(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate956(.a(s_58), .O(gate17inter3));
  inv1  gate957(.a(s_59), .O(gate17inter4));
  nand2 gate958(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate959(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate960(.a(G17), .O(gate17inter7));
  inv1  gate961(.a(G18), .O(gate17inter8));
  nand2 gate962(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate963(.a(s_59), .b(gate17inter3), .O(gate17inter10));
  nor2  gate964(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate965(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate966(.a(gate17inter12), .b(gate17inter1), .O(G290));

  xor2  gate967(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate968(.a(gate18inter0), .b(s_60), .O(gate18inter1));
  and2  gate969(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate970(.a(s_60), .O(gate18inter3));
  inv1  gate971(.a(s_61), .O(gate18inter4));
  nand2 gate972(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate973(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate974(.a(G19), .O(gate18inter7));
  inv1  gate975(.a(G20), .O(gate18inter8));
  nand2 gate976(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate977(.a(s_61), .b(gate18inter3), .O(gate18inter10));
  nor2  gate978(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate979(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate980(.a(gate18inter12), .b(gate18inter1), .O(G293));

  xor2  gate2437(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate2438(.a(gate19inter0), .b(s_270), .O(gate19inter1));
  and2  gate2439(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate2440(.a(s_270), .O(gate19inter3));
  inv1  gate2441(.a(s_271), .O(gate19inter4));
  nand2 gate2442(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate2443(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate2444(.a(G21), .O(gate19inter7));
  inv1  gate2445(.a(G22), .O(gate19inter8));
  nand2 gate2446(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate2447(.a(s_271), .b(gate19inter3), .O(gate19inter10));
  nor2  gate2448(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate2449(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate2450(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate939(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate940(.a(gate23inter0), .b(s_56), .O(gate23inter1));
  and2  gate941(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate942(.a(s_56), .O(gate23inter3));
  inv1  gate943(.a(s_57), .O(gate23inter4));
  nand2 gate944(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate945(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate946(.a(G29), .O(gate23inter7));
  inv1  gate947(.a(G30), .O(gate23inter8));
  nand2 gate948(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate949(.a(s_57), .b(gate23inter3), .O(gate23inter10));
  nor2  gate950(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate951(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate952(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate1205(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate1206(.a(gate25inter0), .b(s_94), .O(gate25inter1));
  and2  gate1207(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate1208(.a(s_94), .O(gate25inter3));
  inv1  gate1209(.a(s_95), .O(gate25inter4));
  nand2 gate1210(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate1211(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate1212(.a(G1), .O(gate25inter7));
  inv1  gate1213(.a(G5), .O(gate25inter8));
  nand2 gate1214(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate1215(.a(s_95), .b(gate25inter3), .O(gate25inter10));
  nor2  gate1216(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate1217(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate1218(.a(gate25inter12), .b(gate25inter1), .O(G314));

  xor2  gate2549(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate2550(.a(gate26inter0), .b(s_286), .O(gate26inter1));
  and2  gate2551(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate2552(.a(s_286), .O(gate26inter3));
  inv1  gate2553(.a(s_287), .O(gate26inter4));
  nand2 gate2554(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate2555(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate2556(.a(G9), .O(gate26inter7));
  inv1  gate2557(.a(G13), .O(gate26inter8));
  nand2 gate2558(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate2559(.a(s_287), .b(gate26inter3), .O(gate26inter10));
  nor2  gate2560(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate2561(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate2562(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate2199(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate2200(.a(gate28inter0), .b(s_236), .O(gate28inter1));
  and2  gate2201(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate2202(.a(s_236), .O(gate28inter3));
  inv1  gate2203(.a(s_237), .O(gate28inter4));
  nand2 gate2204(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate2205(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate2206(.a(G10), .O(gate28inter7));
  inv1  gate2207(.a(G14), .O(gate28inter8));
  nand2 gate2208(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate2209(.a(s_237), .b(gate28inter3), .O(gate28inter10));
  nor2  gate2210(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate2211(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate2212(.a(gate28inter12), .b(gate28inter1), .O(G323));
nand2 gate29( .a(G3), .b(G7), .O(G326) );

  xor2  gate715(.a(G15), .b(G11), .O(gate30inter0));
  nand2 gate716(.a(gate30inter0), .b(s_24), .O(gate30inter1));
  and2  gate717(.a(G15), .b(G11), .O(gate30inter2));
  inv1  gate718(.a(s_24), .O(gate30inter3));
  inv1  gate719(.a(s_25), .O(gate30inter4));
  nand2 gate720(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate721(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate722(.a(G11), .O(gate30inter7));
  inv1  gate723(.a(G15), .O(gate30inter8));
  nand2 gate724(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate725(.a(s_25), .b(gate30inter3), .O(gate30inter10));
  nor2  gate726(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate727(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate728(.a(gate30inter12), .b(gate30inter1), .O(G329));
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate2661(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate2662(.a(gate34inter0), .b(s_302), .O(gate34inter1));
  and2  gate2663(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate2664(.a(s_302), .O(gate34inter3));
  inv1  gate2665(.a(s_303), .O(gate34inter4));
  nand2 gate2666(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate2667(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate2668(.a(G25), .O(gate34inter7));
  inv1  gate2669(.a(G29), .O(gate34inter8));
  nand2 gate2670(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate2671(.a(s_303), .b(gate34inter3), .O(gate34inter10));
  nor2  gate2672(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate2673(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate2674(.a(gate34inter12), .b(gate34inter1), .O(G341));

  xor2  gate1121(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate1122(.a(gate35inter0), .b(s_82), .O(gate35inter1));
  and2  gate1123(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate1124(.a(s_82), .O(gate35inter3));
  inv1  gate1125(.a(s_83), .O(gate35inter4));
  nand2 gate1126(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate1127(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate1128(.a(G18), .O(gate35inter7));
  inv1  gate1129(.a(G22), .O(gate35inter8));
  nand2 gate1130(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate1131(.a(s_83), .b(gate35inter3), .O(gate35inter10));
  nor2  gate1132(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate1133(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate1134(.a(gate35inter12), .b(gate35inter1), .O(G344));
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate2325(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate2326(.a(gate39inter0), .b(s_254), .O(gate39inter1));
  and2  gate2327(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate2328(.a(s_254), .O(gate39inter3));
  inv1  gate2329(.a(s_255), .O(gate39inter4));
  nand2 gate2330(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate2331(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate2332(.a(G20), .O(gate39inter7));
  inv1  gate2333(.a(G24), .O(gate39inter8));
  nand2 gate2334(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate2335(.a(s_255), .b(gate39inter3), .O(gate39inter10));
  nor2  gate2336(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate2337(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate2338(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate561(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate562(.a(gate43inter0), .b(s_2), .O(gate43inter1));
  and2  gate563(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate564(.a(s_2), .O(gate43inter3));
  inv1  gate565(.a(s_3), .O(gate43inter4));
  nand2 gate566(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate567(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate568(.a(G3), .O(gate43inter7));
  inv1  gate569(.a(G269), .O(gate43inter8));
  nand2 gate570(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate571(.a(s_3), .b(gate43inter3), .O(gate43inter10));
  nor2  gate572(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate573(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate574(.a(gate43inter12), .b(gate43inter1), .O(G364));
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );

  xor2  gate1681(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate1682(.a(gate47inter0), .b(s_162), .O(gate47inter1));
  and2  gate1683(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate1684(.a(s_162), .O(gate47inter3));
  inv1  gate1685(.a(s_163), .O(gate47inter4));
  nand2 gate1686(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate1687(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate1688(.a(G7), .O(gate47inter7));
  inv1  gate1689(.a(G275), .O(gate47inter8));
  nand2 gate1690(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate1691(.a(s_163), .b(gate47inter3), .O(gate47inter10));
  nor2  gate1692(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate1693(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate1694(.a(gate47inter12), .b(gate47inter1), .O(G368));
nand2 gate48( .a(G8), .b(G275), .O(G369) );

  xor2  gate2423(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate2424(.a(gate49inter0), .b(s_268), .O(gate49inter1));
  and2  gate2425(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate2426(.a(s_268), .O(gate49inter3));
  inv1  gate2427(.a(s_269), .O(gate49inter4));
  nand2 gate2428(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate2429(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate2430(.a(G9), .O(gate49inter7));
  inv1  gate2431(.a(G278), .O(gate49inter8));
  nand2 gate2432(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate2433(.a(s_269), .b(gate49inter3), .O(gate49inter10));
  nor2  gate2434(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate2435(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate2436(.a(gate49inter12), .b(gate49inter1), .O(G370));

  xor2  gate2213(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate2214(.a(gate50inter0), .b(s_238), .O(gate50inter1));
  and2  gate2215(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate2216(.a(s_238), .O(gate50inter3));
  inv1  gate2217(.a(s_239), .O(gate50inter4));
  nand2 gate2218(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate2219(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate2220(.a(G10), .O(gate50inter7));
  inv1  gate2221(.a(G278), .O(gate50inter8));
  nand2 gate2222(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate2223(.a(s_239), .b(gate50inter3), .O(gate50inter10));
  nor2  gate2224(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate2225(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate2226(.a(gate50inter12), .b(gate50inter1), .O(G371));
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate2745(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate2746(.a(gate52inter0), .b(s_314), .O(gate52inter1));
  and2  gate2747(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate2748(.a(s_314), .O(gate52inter3));
  inv1  gate2749(.a(s_315), .O(gate52inter4));
  nand2 gate2750(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate2751(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate2752(.a(G12), .O(gate52inter7));
  inv1  gate2753(.a(G281), .O(gate52inter8));
  nand2 gate2754(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate2755(.a(s_315), .b(gate52inter3), .O(gate52inter10));
  nor2  gate2756(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate2757(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate2758(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );

  xor2  gate2493(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate2494(.a(gate56inter0), .b(s_278), .O(gate56inter1));
  and2  gate2495(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate2496(.a(s_278), .O(gate56inter3));
  inv1  gate2497(.a(s_279), .O(gate56inter4));
  nand2 gate2498(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate2499(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate2500(.a(G16), .O(gate56inter7));
  inv1  gate2501(.a(G287), .O(gate56inter8));
  nand2 gate2502(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate2503(.a(s_279), .b(gate56inter3), .O(gate56inter10));
  nor2  gate2504(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate2505(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate2506(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate785(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate786(.a(gate63inter0), .b(s_34), .O(gate63inter1));
  and2  gate787(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate788(.a(s_34), .O(gate63inter3));
  inv1  gate789(.a(s_35), .O(gate63inter4));
  nand2 gate790(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate791(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate792(.a(G23), .O(gate63inter7));
  inv1  gate793(.a(G299), .O(gate63inter8));
  nand2 gate794(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate795(.a(s_35), .b(gate63inter3), .O(gate63inter10));
  nor2  gate796(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate797(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate798(.a(gate63inter12), .b(gate63inter1), .O(G384));

  xor2  gate2843(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate2844(.a(gate64inter0), .b(s_328), .O(gate64inter1));
  and2  gate2845(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate2846(.a(s_328), .O(gate64inter3));
  inv1  gate2847(.a(s_329), .O(gate64inter4));
  nand2 gate2848(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate2849(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate2850(.a(G24), .O(gate64inter7));
  inv1  gate2851(.a(G299), .O(gate64inter8));
  nand2 gate2852(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate2853(.a(s_329), .b(gate64inter3), .O(gate64inter10));
  nor2  gate2854(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate2855(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate2856(.a(gate64inter12), .b(gate64inter1), .O(G385));
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate1149(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate1150(.a(gate69inter0), .b(s_86), .O(gate69inter1));
  and2  gate1151(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate1152(.a(s_86), .O(gate69inter3));
  inv1  gate1153(.a(s_87), .O(gate69inter4));
  nand2 gate1154(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate1155(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate1156(.a(G29), .O(gate69inter7));
  inv1  gate1157(.a(G308), .O(gate69inter8));
  nand2 gate1158(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate1159(.a(s_87), .b(gate69inter3), .O(gate69inter10));
  nor2  gate1160(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate1161(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate1162(.a(gate69inter12), .b(gate69inter1), .O(G390));

  xor2  gate1345(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate1346(.a(gate70inter0), .b(s_114), .O(gate70inter1));
  and2  gate1347(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate1348(.a(s_114), .O(gate70inter3));
  inv1  gate1349(.a(s_115), .O(gate70inter4));
  nand2 gate1350(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate1351(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate1352(.a(G30), .O(gate70inter7));
  inv1  gate1353(.a(G308), .O(gate70inter8));
  nand2 gate1354(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate1355(.a(s_115), .b(gate70inter3), .O(gate70inter10));
  nor2  gate1356(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate1357(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate1358(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );

  xor2  gate1653(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate1654(.a(gate73inter0), .b(s_158), .O(gate73inter1));
  and2  gate1655(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate1656(.a(s_158), .O(gate73inter3));
  inv1  gate1657(.a(s_159), .O(gate73inter4));
  nand2 gate1658(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate1659(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate1660(.a(G1), .O(gate73inter7));
  inv1  gate1661(.a(G314), .O(gate73inter8));
  nand2 gate1662(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate1663(.a(s_159), .b(gate73inter3), .O(gate73inter10));
  nor2  gate1664(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate1665(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate1666(.a(gate73inter12), .b(gate73inter1), .O(G394));
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );

  xor2  gate701(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate702(.a(gate76inter0), .b(s_22), .O(gate76inter1));
  and2  gate703(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate704(.a(s_22), .O(gate76inter3));
  inv1  gate705(.a(s_23), .O(gate76inter4));
  nand2 gate706(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate707(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate708(.a(G13), .O(gate76inter7));
  inv1  gate709(.a(G317), .O(gate76inter8));
  nand2 gate710(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate711(.a(s_23), .b(gate76inter3), .O(gate76inter10));
  nor2  gate712(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate713(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate714(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );

  xor2  gate841(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate842(.a(gate79inter0), .b(s_42), .O(gate79inter1));
  and2  gate843(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate844(.a(s_42), .O(gate79inter3));
  inv1  gate845(.a(s_43), .O(gate79inter4));
  nand2 gate846(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate847(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate848(.a(G10), .O(gate79inter7));
  inv1  gate849(.a(G323), .O(gate79inter8));
  nand2 gate850(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate851(.a(s_43), .b(gate79inter3), .O(gate79inter10));
  nor2  gate852(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate853(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate854(.a(gate79inter12), .b(gate79inter1), .O(G400));

  xor2  gate2073(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate2074(.a(gate80inter0), .b(s_218), .O(gate80inter1));
  and2  gate2075(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate2076(.a(s_218), .O(gate80inter3));
  inv1  gate2077(.a(s_219), .O(gate80inter4));
  nand2 gate2078(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate2079(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate2080(.a(G14), .O(gate80inter7));
  inv1  gate2081(.a(G323), .O(gate80inter8));
  nand2 gate2082(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate2083(.a(s_219), .b(gate80inter3), .O(gate80inter10));
  nor2  gate2084(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate2085(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate2086(.a(gate80inter12), .b(gate80inter1), .O(G401));

  xor2  gate2871(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate2872(.a(gate81inter0), .b(s_332), .O(gate81inter1));
  and2  gate2873(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate2874(.a(s_332), .O(gate81inter3));
  inv1  gate2875(.a(s_333), .O(gate81inter4));
  nand2 gate2876(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate2877(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate2878(.a(G3), .O(gate81inter7));
  inv1  gate2879(.a(G326), .O(gate81inter8));
  nand2 gate2880(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate2881(.a(s_333), .b(gate81inter3), .O(gate81inter10));
  nor2  gate2882(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate2883(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate2884(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );

  xor2  gate1555(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate1556(.a(gate84inter0), .b(s_144), .O(gate84inter1));
  and2  gate1557(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate1558(.a(s_144), .O(gate84inter3));
  inv1  gate1559(.a(s_145), .O(gate84inter4));
  nand2 gate1560(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate1561(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate1562(.a(G15), .O(gate84inter7));
  inv1  gate1563(.a(G329), .O(gate84inter8));
  nand2 gate1564(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate1565(.a(s_145), .b(gate84inter3), .O(gate84inter10));
  nor2  gate1566(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate1567(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate1568(.a(gate84inter12), .b(gate84inter1), .O(G405));

  xor2  gate1779(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate1780(.a(gate85inter0), .b(s_176), .O(gate85inter1));
  and2  gate1781(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate1782(.a(s_176), .O(gate85inter3));
  inv1  gate1783(.a(s_177), .O(gate85inter4));
  nand2 gate1784(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate1785(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate1786(.a(G4), .O(gate85inter7));
  inv1  gate1787(.a(G332), .O(gate85inter8));
  nand2 gate1788(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate1789(.a(s_177), .b(gate85inter3), .O(gate85inter10));
  nor2  gate1790(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate1791(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate1792(.a(gate85inter12), .b(gate85inter1), .O(G406));
nand2 gate86( .a(G8), .b(G332), .O(G407) );

  xor2  gate2031(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate2032(.a(gate87inter0), .b(s_212), .O(gate87inter1));
  and2  gate2033(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate2034(.a(s_212), .O(gate87inter3));
  inv1  gate2035(.a(s_213), .O(gate87inter4));
  nand2 gate2036(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate2037(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate2038(.a(G12), .O(gate87inter7));
  inv1  gate2039(.a(G335), .O(gate87inter8));
  nand2 gate2040(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate2041(.a(s_213), .b(gate87inter3), .O(gate87inter10));
  nor2  gate2042(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate2043(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate2044(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate2241(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate2242(.a(gate91inter0), .b(s_242), .O(gate91inter1));
  and2  gate2243(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate2244(.a(s_242), .O(gate91inter3));
  inv1  gate2245(.a(s_243), .O(gate91inter4));
  nand2 gate2246(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate2247(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate2248(.a(G25), .O(gate91inter7));
  inv1  gate2249(.a(G341), .O(gate91inter8));
  nand2 gate2250(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate2251(.a(s_243), .b(gate91inter3), .O(gate91inter10));
  nor2  gate2252(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate2253(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate2254(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );

  xor2  gate1135(.a(G350), .b(G19), .O(gate97inter0));
  nand2 gate1136(.a(gate97inter0), .b(s_84), .O(gate97inter1));
  and2  gate1137(.a(G350), .b(G19), .O(gate97inter2));
  inv1  gate1138(.a(s_84), .O(gate97inter3));
  inv1  gate1139(.a(s_85), .O(gate97inter4));
  nand2 gate1140(.a(gate97inter4), .b(gate97inter3), .O(gate97inter5));
  nor2  gate1141(.a(gate97inter5), .b(gate97inter2), .O(gate97inter6));
  inv1  gate1142(.a(G19), .O(gate97inter7));
  inv1  gate1143(.a(G350), .O(gate97inter8));
  nand2 gate1144(.a(gate97inter8), .b(gate97inter7), .O(gate97inter9));
  nand2 gate1145(.a(s_85), .b(gate97inter3), .O(gate97inter10));
  nor2  gate1146(.a(gate97inter10), .b(gate97inter9), .O(gate97inter11));
  nor2  gate1147(.a(gate97inter11), .b(gate97inter6), .O(gate97inter12));
  nand2 gate1148(.a(gate97inter12), .b(gate97inter1), .O(G418));

  xor2  gate757(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate758(.a(gate98inter0), .b(s_30), .O(gate98inter1));
  and2  gate759(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate760(.a(s_30), .O(gate98inter3));
  inv1  gate761(.a(s_31), .O(gate98inter4));
  nand2 gate762(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate763(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate764(.a(G23), .O(gate98inter7));
  inv1  gate765(.a(G350), .O(gate98inter8));
  nand2 gate766(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate767(.a(s_31), .b(gate98inter3), .O(gate98inter10));
  nor2  gate768(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate769(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate770(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate1415(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate1416(.a(gate100inter0), .b(s_124), .O(gate100inter1));
  and2  gate1417(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate1418(.a(s_124), .O(gate100inter3));
  inv1  gate1419(.a(s_125), .O(gate100inter4));
  nand2 gate1420(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate1421(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate1422(.a(G31), .O(gate100inter7));
  inv1  gate1423(.a(G353), .O(gate100inter8));
  nand2 gate1424(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate1425(.a(s_125), .b(gate100inter3), .O(gate100inter10));
  nor2  gate1426(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate1427(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate1428(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate1877(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate1878(.a(gate102inter0), .b(s_190), .O(gate102inter1));
  and2  gate1879(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate1880(.a(s_190), .O(gate102inter3));
  inv1  gate1881(.a(s_191), .O(gate102inter4));
  nand2 gate1882(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate1883(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate1884(.a(G24), .O(gate102inter7));
  inv1  gate1885(.a(G356), .O(gate102inter8));
  nand2 gate1886(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate1887(.a(s_191), .b(gate102inter3), .O(gate102inter10));
  nor2  gate1888(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate1889(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate1890(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate603(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate604(.a(gate104inter0), .b(s_8), .O(gate104inter1));
  and2  gate605(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate606(.a(s_8), .O(gate104inter3));
  inv1  gate607(.a(s_9), .O(gate104inter4));
  nand2 gate608(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate609(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate610(.a(G32), .O(gate104inter7));
  inv1  gate611(.a(G359), .O(gate104inter8));
  nand2 gate612(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate613(.a(s_9), .b(gate104inter3), .O(gate104inter10));
  nor2  gate614(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate615(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate616(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate2857(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate2858(.a(gate107inter0), .b(s_330), .O(gate107inter1));
  and2  gate2859(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate2860(.a(s_330), .O(gate107inter3));
  inv1  gate2861(.a(s_331), .O(gate107inter4));
  nand2 gate2862(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate2863(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate2864(.a(G366), .O(gate107inter7));
  inv1  gate2865(.a(G367), .O(gate107inter8));
  nand2 gate2866(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate2867(.a(s_331), .b(gate107inter3), .O(gate107inter10));
  nor2  gate2868(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate2869(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate2870(.a(gate107inter12), .b(gate107inter1), .O(G432));

  xor2  gate687(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate688(.a(gate108inter0), .b(s_20), .O(gate108inter1));
  and2  gate689(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate690(.a(s_20), .O(gate108inter3));
  inv1  gate691(.a(s_21), .O(gate108inter4));
  nand2 gate692(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate693(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate694(.a(G368), .O(gate108inter7));
  inv1  gate695(.a(G369), .O(gate108inter8));
  nand2 gate696(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate697(.a(s_21), .b(gate108inter3), .O(gate108inter10));
  nor2  gate698(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate699(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate700(.a(gate108inter12), .b(gate108inter1), .O(G435));
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );

  xor2  gate1093(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate1094(.a(gate111inter0), .b(s_78), .O(gate111inter1));
  and2  gate1095(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate1096(.a(s_78), .O(gate111inter3));
  inv1  gate1097(.a(s_79), .O(gate111inter4));
  nand2 gate1098(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate1099(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate1100(.a(G374), .O(gate111inter7));
  inv1  gate1101(.a(G375), .O(gate111inter8));
  nand2 gate1102(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate1103(.a(s_79), .b(gate111inter3), .O(gate111inter10));
  nor2  gate1104(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate1105(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate1106(.a(gate111inter12), .b(gate111inter1), .O(G444));

  xor2  gate2997(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate2998(.a(gate112inter0), .b(s_350), .O(gate112inter1));
  and2  gate2999(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate3000(.a(s_350), .O(gate112inter3));
  inv1  gate3001(.a(s_351), .O(gate112inter4));
  nand2 gate3002(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate3003(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate3004(.a(G376), .O(gate112inter7));
  inv1  gate3005(.a(G377), .O(gate112inter8));
  nand2 gate3006(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate3007(.a(s_351), .b(gate112inter3), .O(gate112inter10));
  nor2  gate3008(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate3009(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate3010(.a(gate112inter12), .b(gate112inter1), .O(G447));
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate2577(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate2578(.a(gate117inter0), .b(s_290), .O(gate117inter1));
  and2  gate2579(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate2580(.a(s_290), .O(gate117inter3));
  inv1  gate2581(.a(s_291), .O(gate117inter4));
  nand2 gate2582(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate2583(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate2584(.a(G386), .O(gate117inter7));
  inv1  gate2585(.a(G387), .O(gate117inter8));
  nand2 gate2586(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate2587(.a(s_291), .b(gate117inter3), .O(gate117inter10));
  nor2  gate2588(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate2589(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate2590(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate2507(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate2508(.a(gate125inter0), .b(s_280), .O(gate125inter1));
  and2  gate2509(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate2510(.a(s_280), .O(gate125inter3));
  inv1  gate2511(.a(s_281), .O(gate125inter4));
  nand2 gate2512(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate2513(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate2514(.a(G402), .O(gate125inter7));
  inv1  gate2515(.a(G403), .O(gate125inter8));
  nand2 gate2516(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate2517(.a(s_281), .b(gate125inter3), .O(gate125inter10));
  nor2  gate2518(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate2519(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate2520(.a(gate125inter12), .b(gate125inter1), .O(G486));

  xor2  gate2983(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate2984(.a(gate126inter0), .b(s_348), .O(gate126inter1));
  and2  gate2985(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate2986(.a(s_348), .O(gate126inter3));
  inv1  gate2987(.a(s_349), .O(gate126inter4));
  nand2 gate2988(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate2989(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate2990(.a(G404), .O(gate126inter7));
  inv1  gate2991(.a(G405), .O(gate126inter8));
  nand2 gate2992(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate2993(.a(s_349), .b(gate126inter3), .O(gate126inter10));
  nor2  gate2994(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate2995(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate2996(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );

  xor2  gate2759(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate2760(.a(gate129inter0), .b(s_316), .O(gate129inter1));
  and2  gate2761(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate2762(.a(s_316), .O(gate129inter3));
  inv1  gate2763(.a(s_317), .O(gate129inter4));
  nand2 gate2764(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate2765(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate2766(.a(G410), .O(gate129inter7));
  inv1  gate2767(.a(G411), .O(gate129inter8));
  nand2 gate2768(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate2769(.a(s_317), .b(gate129inter3), .O(gate129inter10));
  nor2  gate2770(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate2771(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate2772(.a(gate129inter12), .b(gate129inter1), .O(G498));
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate2045(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate2046(.a(gate131inter0), .b(s_214), .O(gate131inter1));
  and2  gate2047(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate2048(.a(s_214), .O(gate131inter3));
  inv1  gate2049(.a(s_215), .O(gate131inter4));
  nand2 gate2050(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate2051(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate2052(.a(G414), .O(gate131inter7));
  inv1  gate2053(.a(G415), .O(gate131inter8));
  nand2 gate2054(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate2055(.a(s_215), .b(gate131inter3), .O(gate131inter10));
  nor2  gate2056(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate2057(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate2058(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );

  xor2  gate547(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate548(.a(gate133inter0), .b(s_0), .O(gate133inter1));
  and2  gate549(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate550(.a(s_0), .O(gate133inter3));
  inv1  gate551(.a(s_1), .O(gate133inter4));
  nand2 gate552(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate553(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate554(.a(G418), .O(gate133inter7));
  inv1  gate555(.a(G419), .O(gate133inter8));
  nand2 gate556(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate557(.a(s_1), .b(gate133inter3), .O(gate133inter10));
  nor2  gate558(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate559(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate560(.a(gate133inter12), .b(gate133inter1), .O(G510));

  xor2  gate2479(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate2480(.a(gate134inter0), .b(s_276), .O(gate134inter1));
  and2  gate2481(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate2482(.a(s_276), .O(gate134inter3));
  inv1  gate2483(.a(s_277), .O(gate134inter4));
  nand2 gate2484(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate2485(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate2486(.a(G420), .O(gate134inter7));
  inv1  gate2487(.a(G421), .O(gate134inter8));
  nand2 gate2488(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate2489(.a(s_277), .b(gate134inter3), .O(gate134inter10));
  nor2  gate2490(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate2491(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate2492(.a(gate134inter12), .b(gate134inter1), .O(G513));

  xor2  gate1541(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate1542(.a(gate135inter0), .b(s_142), .O(gate135inter1));
  and2  gate1543(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate1544(.a(s_142), .O(gate135inter3));
  inv1  gate1545(.a(s_143), .O(gate135inter4));
  nand2 gate1546(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate1547(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate1548(.a(G422), .O(gate135inter7));
  inv1  gate1549(.a(G423), .O(gate135inter8));
  nand2 gate1550(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate1551(.a(s_143), .b(gate135inter3), .O(gate135inter10));
  nor2  gate1552(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate1553(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate1554(.a(gate135inter12), .b(gate135inter1), .O(G516));

  xor2  gate673(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate674(.a(gate136inter0), .b(s_18), .O(gate136inter1));
  and2  gate675(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate676(.a(s_18), .O(gate136inter3));
  inv1  gate677(.a(s_19), .O(gate136inter4));
  nand2 gate678(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate679(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate680(.a(G424), .O(gate136inter7));
  inv1  gate681(.a(G425), .O(gate136inter8));
  nand2 gate682(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate683(.a(s_19), .b(gate136inter3), .O(gate136inter10));
  nor2  gate684(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate685(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate686(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );

  xor2  gate1807(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate1808(.a(gate140inter0), .b(s_180), .O(gate140inter1));
  and2  gate1809(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate1810(.a(s_180), .O(gate140inter3));
  inv1  gate1811(.a(s_181), .O(gate140inter4));
  nand2 gate1812(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate1813(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate1814(.a(G444), .O(gate140inter7));
  inv1  gate1815(.a(G447), .O(gate140inter8));
  nand2 gate1816(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate1817(.a(s_181), .b(gate140inter3), .O(gate140inter10));
  nor2  gate1818(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate1819(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate1820(.a(gate140inter12), .b(gate140inter1), .O(G531));

  xor2  gate617(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate618(.a(gate141inter0), .b(s_10), .O(gate141inter1));
  and2  gate619(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate620(.a(s_10), .O(gate141inter3));
  inv1  gate621(.a(s_11), .O(gate141inter4));
  nand2 gate622(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate623(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate624(.a(G450), .O(gate141inter7));
  inv1  gate625(.a(G453), .O(gate141inter8));
  nand2 gate626(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate627(.a(s_11), .b(gate141inter3), .O(gate141inter10));
  nor2  gate628(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate629(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate630(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );

  xor2  gate1471(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate1472(.a(gate145inter0), .b(s_132), .O(gate145inter1));
  and2  gate1473(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate1474(.a(s_132), .O(gate145inter3));
  inv1  gate1475(.a(s_133), .O(gate145inter4));
  nand2 gate1476(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate1477(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate1478(.a(G474), .O(gate145inter7));
  inv1  gate1479(.a(G477), .O(gate145inter8));
  nand2 gate1480(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate1481(.a(s_133), .b(gate145inter3), .O(gate145inter10));
  nor2  gate1482(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate1483(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate1484(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate1765(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1766(.a(gate148inter0), .b(s_174), .O(gate148inter1));
  and2  gate1767(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1768(.a(s_174), .O(gate148inter3));
  inv1  gate1769(.a(s_175), .O(gate148inter4));
  nand2 gate1770(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1771(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1772(.a(G492), .O(gate148inter7));
  inv1  gate1773(.a(G495), .O(gate148inter8));
  nand2 gate1774(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1775(.a(s_175), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1776(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1777(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1778(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate1667(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate1668(.a(gate150inter0), .b(s_160), .O(gate150inter1));
  and2  gate1669(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate1670(.a(s_160), .O(gate150inter3));
  inv1  gate1671(.a(s_161), .O(gate150inter4));
  nand2 gate1672(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate1673(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate1674(.a(G504), .O(gate150inter7));
  inv1  gate1675(.a(G507), .O(gate150inter8));
  nand2 gate1676(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate1677(.a(s_161), .b(gate150inter3), .O(gate150inter10));
  nor2  gate1678(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate1679(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate1680(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate1289(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate1290(.a(gate153inter0), .b(s_106), .O(gate153inter1));
  and2  gate1291(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate1292(.a(s_106), .O(gate153inter3));
  inv1  gate1293(.a(s_107), .O(gate153inter4));
  nand2 gate1294(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate1295(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate1296(.a(G426), .O(gate153inter7));
  inv1  gate1297(.a(G522), .O(gate153inter8));
  nand2 gate1298(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate1299(.a(s_107), .b(gate153inter3), .O(gate153inter10));
  nor2  gate1300(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate1301(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate1302(.a(gate153inter12), .b(gate153inter1), .O(G570));

  xor2  gate2283(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate2284(.a(gate154inter0), .b(s_248), .O(gate154inter1));
  and2  gate2285(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate2286(.a(s_248), .O(gate154inter3));
  inv1  gate2287(.a(s_249), .O(gate154inter4));
  nand2 gate2288(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate2289(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate2290(.a(G429), .O(gate154inter7));
  inv1  gate2291(.a(G522), .O(gate154inter8));
  nand2 gate2292(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate2293(.a(s_249), .b(gate154inter3), .O(gate154inter10));
  nor2  gate2294(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate2295(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate2296(.a(gate154inter12), .b(gate154inter1), .O(G571));

  xor2  gate1723(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate1724(.a(gate155inter0), .b(s_168), .O(gate155inter1));
  and2  gate1725(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate1726(.a(s_168), .O(gate155inter3));
  inv1  gate1727(.a(s_169), .O(gate155inter4));
  nand2 gate1728(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1729(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1730(.a(G432), .O(gate155inter7));
  inv1  gate1731(.a(G525), .O(gate155inter8));
  nand2 gate1732(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1733(.a(s_169), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1734(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1735(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1736(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate813(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate814(.a(gate157inter0), .b(s_38), .O(gate157inter1));
  and2  gate815(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate816(.a(s_38), .O(gate157inter3));
  inv1  gate817(.a(s_39), .O(gate157inter4));
  nand2 gate818(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate819(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate820(.a(G438), .O(gate157inter7));
  inv1  gate821(.a(G528), .O(gate157inter8));
  nand2 gate822(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate823(.a(s_39), .b(gate157inter3), .O(gate157inter10));
  nor2  gate824(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate825(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate826(.a(gate157inter12), .b(gate157inter1), .O(G574));

  xor2  gate1387(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate1388(.a(gate158inter0), .b(s_120), .O(gate158inter1));
  and2  gate1389(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate1390(.a(s_120), .O(gate158inter3));
  inv1  gate1391(.a(s_121), .O(gate158inter4));
  nand2 gate1392(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate1393(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate1394(.a(G441), .O(gate158inter7));
  inv1  gate1395(.a(G528), .O(gate158inter8));
  nand2 gate1396(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate1397(.a(s_121), .b(gate158inter3), .O(gate158inter10));
  nor2  gate1398(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate1399(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate1400(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate2129(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate2130(.a(gate162inter0), .b(s_226), .O(gate162inter1));
  and2  gate2131(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate2132(.a(s_226), .O(gate162inter3));
  inv1  gate2133(.a(s_227), .O(gate162inter4));
  nand2 gate2134(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate2135(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate2136(.a(G453), .O(gate162inter7));
  inv1  gate2137(.a(G534), .O(gate162inter8));
  nand2 gate2138(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate2139(.a(s_227), .b(gate162inter3), .O(gate162inter10));
  nor2  gate2140(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate2141(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate2142(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate2829(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate2830(.a(gate164inter0), .b(s_326), .O(gate164inter1));
  and2  gate2831(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate2832(.a(s_326), .O(gate164inter3));
  inv1  gate2833(.a(s_327), .O(gate164inter4));
  nand2 gate2834(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate2835(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate2836(.a(G459), .O(gate164inter7));
  inv1  gate2837(.a(G537), .O(gate164inter8));
  nand2 gate2838(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate2839(.a(s_327), .b(gate164inter3), .O(gate164inter10));
  nor2  gate2840(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate2841(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate2842(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );

  xor2  gate1975(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate1976(.a(gate166inter0), .b(s_204), .O(gate166inter1));
  and2  gate1977(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate1978(.a(s_204), .O(gate166inter3));
  inv1  gate1979(.a(s_205), .O(gate166inter4));
  nand2 gate1980(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate1981(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate1982(.a(G465), .O(gate166inter7));
  inv1  gate1983(.a(G540), .O(gate166inter8));
  nand2 gate1984(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate1985(.a(s_205), .b(gate166inter3), .O(gate166inter10));
  nor2  gate1986(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate1987(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate1988(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );

  xor2  gate1051(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate1052(.a(gate168inter0), .b(s_72), .O(gate168inter1));
  and2  gate1053(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate1054(.a(s_72), .O(gate168inter3));
  inv1  gate1055(.a(s_73), .O(gate168inter4));
  nand2 gate1056(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate1057(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate1058(.a(G471), .O(gate168inter7));
  inv1  gate1059(.a(G543), .O(gate168inter8));
  nand2 gate1060(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate1061(.a(s_73), .b(gate168inter3), .O(gate168inter10));
  nor2  gate1062(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate1063(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate1064(.a(gate168inter12), .b(gate168inter1), .O(G585));
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate2297(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate2298(.a(gate173inter0), .b(s_250), .O(gate173inter1));
  and2  gate2299(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate2300(.a(s_250), .O(gate173inter3));
  inv1  gate2301(.a(s_251), .O(gate173inter4));
  nand2 gate2302(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate2303(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate2304(.a(G486), .O(gate173inter7));
  inv1  gate2305(.a(G552), .O(gate173inter8));
  nand2 gate2306(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate2307(.a(s_251), .b(gate173inter3), .O(gate173inter10));
  nor2  gate2308(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate2309(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate2310(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );

  xor2  gate1695(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate1696(.a(gate177inter0), .b(s_164), .O(gate177inter1));
  and2  gate1697(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate1698(.a(s_164), .O(gate177inter3));
  inv1  gate1699(.a(s_165), .O(gate177inter4));
  nand2 gate1700(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate1701(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate1702(.a(G498), .O(gate177inter7));
  inv1  gate1703(.a(G558), .O(gate177inter8));
  nand2 gate1704(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate1705(.a(s_165), .b(gate177inter3), .O(gate177inter10));
  nor2  gate1706(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate1707(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate1708(.a(gate177inter12), .b(gate177inter1), .O(G594));
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate1639(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate1640(.a(gate180inter0), .b(s_156), .O(gate180inter1));
  and2  gate1641(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate1642(.a(s_156), .O(gate180inter3));
  inv1  gate1643(.a(s_157), .O(gate180inter4));
  nand2 gate1644(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate1645(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate1646(.a(G507), .O(gate180inter7));
  inv1  gate1647(.a(G561), .O(gate180inter8));
  nand2 gate1648(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate1649(.a(s_157), .b(gate180inter3), .O(gate180inter10));
  nor2  gate1650(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate1651(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate1652(.a(gate180inter12), .b(gate180inter1), .O(G597));

  xor2  gate799(.a(G564), .b(G510), .O(gate181inter0));
  nand2 gate800(.a(gate181inter0), .b(s_36), .O(gate181inter1));
  and2  gate801(.a(G564), .b(G510), .O(gate181inter2));
  inv1  gate802(.a(s_36), .O(gate181inter3));
  inv1  gate803(.a(s_37), .O(gate181inter4));
  nand2 gate804(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate805(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate806(.a(G510), .O(gate181inter7));
  inv1  gate807(.a(G564), .O(gate181inter8));
  nand2 gate808(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate809(.a(s_37), .b(gate181inter3), .O(gate181inter10));
  nor2  gate810(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate811(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate812(.a(gate181inter12), .b(gate181inter1), .O(G598));

  xor2  gate2969(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate2970(.a(gate182inter0), .b(s_346), .O(gate182inter1));
  and2  gate2971(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate2972(.a(s_346), .O(gate182inter3));
  inv1  gate2973(.a(s_347), .O(gate182inter4));
  nand2 gate2974(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate2975(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate2976(.a(G513), .O(gate182inter7));
  inv1  gate2977(.a(G564), .O(gate182inter8));
  nand2 gate2978(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate2979(.a(s_347), .b(gate182inter3), .O(gate182inter10));
  nor2  gate2980(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate2981(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate2982(.a(gate182inter12), .b(gate182inter1), .O(G599));

  xor2  gate1107(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate1108(.a(gate183inter0), .b(s_80), .O(gate183inter1));
  and2  gate1109(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate1110(.a(s_80), .O(gate183inter3));
  inv1  gate1111(.a(s_81), .O(gate183inter4));
  nand2 gate1112(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate1113(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate1114(.a(G516), .O(gate183inter7));
  inv1  gate1115(.a(G567), .O(gate183inter8));
  nand2 gate1116(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate1117(.a(s_81), .b(gate183inter3), .O(gate183inter10));
  nor2  gate1118(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate1119(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate1120(.a(gate183inter12), .b(gate183inter1), .O(G600));

  xor2  gate2115(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate2116(.a(gate184inter0), .b(s_224), .O(gate184inter1));
  and2  gate2117(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate2118(.a(s_224), .O(gate184inter3));
  inv1  gate2119(.a(s_225), .O(gate184inter4));
  nand2 gate2120(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate2121(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate2122(.a(G519), .O(gate184inter7));
  inv1  gate2123(.a(G567), .O(gate184inter8));
  nand2 gate2124(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate2125(.a(s_225), .b(gate184inter3), .O(gate184inter10));
  nor2  gate2126(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate2127(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate2128(.a(gate184inter12), .b(gate184inter1), .O(G601));

  xor2  gate729(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate730(.a(gate185inter0), .b(s_26), .O(gate185inter1));
  and2  gate731(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate732(.a(s_26), .O(gate185inter3));
  inv1  gate733(.a(s_27), .O(gate185inter4));
  nand2 gate734(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate735(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate736(.a(G570), .O(gate185inter7));
  inv1  gate737(.a(G571), .O(gate185inter8));
  nand2 gate738(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate739(.a(s_27), .b(gate185inter3), .O(gate185inter10));
  nor2  gate740(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate741(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate742(.a(gate185inter12), .b(gate185inter1), .O(G602));
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate925(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate926(.a(gate187inter0), .b(s_54), .O(gate187inter1));
  and2  gate927(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate928(.a(s_54), .O(gate187inter3));
  inv1  gate929(.a(s_55), .O(gate187inter4));
  nand2 gate930(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate931(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate932(.a(G574), .O(gate187inter7));
  inv1  gate933(.a(G575), .O(gate187inter8));
  nand2 gate934(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate935(.a(s_55), .b(gate187inter3), .O(gate187inter10));
  nor2  gate936(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate937(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate938(.a(gate187inter12), .b(gate187inter1), .O(G612));

  xor2  gate2885(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate2886(.a(gate188inter0), .b(s_334), .O(gate188inter1));
  and2  gate2887(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate2888(.a(s_334), .O(gate188inter3));
  inv1  gate2889(.a(s_335), .O(gate188inter4));
  nand2 gate2890(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate2891(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate2892(.a(G576), .O(gate188inter7));
  inv1  gate2893(.a(G577), .O(gate188inter8));
  nand2 gate2894(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate2895(.a(s_335), .b(gate188inter3), .O(gate188inter10));
  nor2  gate2896(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate2897(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate2898(.a(gate188inter12), .b(gate188inter1), .O(G617));

  xor2  gate2633(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate2634(.a(gate189inter0), .b(s_298), .O(gate189inter1));
  and2  gate2635(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate2636(.a(s_298), .O(gate189inter3));
  inv1  gate2637(.a(s_299), .O(gate189inter4));
  nand2 gate2638(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate2639(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate2640(.a(G578), .O(gate189inter7));
  inv1  gate2641(.a(G579), .O(gate189inter8));
  nand2 gate2642(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate2643(.a(s_299), .b(gate189inter3), .O(gate189inter10));
  nor2  gate2644(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate2645(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate2646(.a(gate189inter12), .b(gate189inter1), .O(G622));
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate2731(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate2732(.a(gate191inter0), .b(s_312), .O(gate191inter1));
  and2  gate2733(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate2734(.a(s_312), .O(gate191inter3));
  inv1  gate2735(.a(s_313), .O(gate191inter4));
  nand2 gate2736(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate2737(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate2738(.a(G582), .O(gate191inter7));
  inv1  gate2739(.a(G583), .O(gate191inter8));
  nand2 gate2740(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate2741(.a(s_313), .b(gate191inter3), .O(gate191inter10));
  nor2  gate2742(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate2743(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate2744(.a(gate191inter12), .b(gate191inter1), .O(G632));

  xor2  gate1625(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate1626(.a(gate192inter0), .b(s_154), .O(gate192inter1));
  and2  gate1627(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate1628(.a(s_154), .O(gate192inter3));
  inv1  gate1629(.a(s_155), .O(gate192inter4));
  nand2 gate1630(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate1631(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate1632(.a(G584), .O(gate192inter7));
  inv1  gate1633(.a(G585), .O(gate192inter8));
  nand2 gate1634(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate1635(.a(s_155), .b(gate192inter3), .O(gate192inter10));
  nor2  gate1636(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate1637(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate1638(.a(gate192inter12), .b(gate192inter1), .O(G637));

  xor2  gate2395(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate2396(.a(gate193inter0), .b(s_264), .O(gate193inter1));
  and2  gate2397(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate2398(.a(s_264), .O(gate193inter3));
  inv1  gate2399(.a(s_265), .O(gate193inter4));
  nand2 gate2400(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate2401(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate2402(.a(G586), .O(gate193inter7));
  inv1  gate2403(.a(G587), .O(gate193inter8));
  nand2 gate2404(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate2405(.a(s_265), .b(gate193inter3), .O(gate193inter10));
  nor2  gate2406(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate2407(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate2408(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate2227(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate2228(.a(gate197inter0), .b(s_240), .O(gate197inter1));
  and2  gate2229(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate2230(.a(s_240), .O(gate197inter3));
  inv1  gate2231(.a(s_241), .O(gate197inter4));
  nand2 gate2232(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate2233(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate2234(.a(G594), .O(gate197inter7));
  inv1  gate2235(.a(G595), .O(gate197inter8));
  nand2 gate2236(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate2237(.a(s_241), .b(gate197inter3), .O(gate197inter10));
  nor2  gate2238(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate2239(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate2240(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate1933(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate1934(.a(gate200inter0), .b(s_198), .O(gate200inter1));
  and2  gate1935(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate1936(.a(s_198), .O(gate200inter3));
  inv1  gate1937(.a(s_199), .O(gate200inter4));
  nand2 gate1938(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate1939(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate1940(.a(G600), .O(gate200inter7));
  inv1  gate1941(.a(G601), .O(gate200inter8));
  nand2 gate1942(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate1943(.a(s_199), .b(gate200inter3), .O(gate200inter10));
  nor2  gate1944(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate1945(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate1946(.a(gate200inter12), .b(gate200inter1), .O(G663));

  xor2  gate1303(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate1304(.a(gate201inter0), .b(s_108), .O(gate201inter1));
  and2  gate1305(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate1306(.a(s_108), .O(gate201inter3));
  inv1  gate1307(.a(s_109), .O(gate201inter4));
  nand2 gate1308(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate1309(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate1310(.a(G602), .O(gate201inter7));
  inv1  gate1311(.a(G607), .O(gate201inter8));
  nand2 gate1312(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate1313(.a(s_109), .b(gate201inter3), .O(gate201inter10));
  nor2  gate1314(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate1315(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate1316(.a(gate201inter12), .b(gate201inter1), .O(G666));

  xor2  gate1275(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate1276(.a(gate202inter0), .b(s_104), .O(gate202inter1));
  and2  gate1277(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate1278(.a(s_104), .O(gate202inter3));
  inv1  gate1279(.a(s_105), .O(gate202inter4));
  nand2 gate1280(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate1281(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate1282(.a(G612), .O(gate202inter7));
  inv1  gate1283(.a(G617), .O(gate202inter8));
  nand2 gate1284(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate1285(.a(s_105), .b(gate202inter3), .O(gate202inter10));
  nor2  gate1286(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate1287(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate1288(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate2717(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate2718(.a(gate205inter0), .b(s_310), .O(gate205inter1));
  and2  gate2719(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate2720(.a(s_310), .O(gate205inter3));
  inv1  gate2721(.a(s_311), .O(gate205inter4));
  nand2 gate2722(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate2723(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate2724(.a(G622), .O(gate205inter7));
  inv1  gate2725(.a(G627), .O(gate205inter8));
  nand2 gate2726(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate2727(.a(s_311), .b(gate205inter3), .O(gate205inter10));
  nor2  gate2728(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate2729(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate2730(.a(gate205inter12), .b(gate205inter1), .O(G678));

  xor2  gate2773(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate2774(.a(gate206inter0), .b(s_318), .O(gate206inter1));
  and2  gate2775(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate2776(.a(s_318), .O(gate206inter3));
  inv1  gate2777(.a(s_319), .O(gate206inter4));
  nand2 gate2778(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate2779(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate2780(.a(G632), .O(gate206inter7));
  inv1  gate2781(.a(G637), .O(gate206inter8));
  nand2 gate2782(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate2783(.a(s_319), .b(gate206inter3), .O(gate206inter10));
  nor2  gate2784(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate2785(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate2786(.a(gate206inter12), .b(gate206inter1), .O(G681));

  xor2  gate1583(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate1584(.a(gate207inter0), .b(s_148), .O(gate207inter1));
  and2  gate1585(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate1586(.a(s_148), .O(gate207inter3));
  inv1  gate1587(.a(s_149), .O(gate207inter4));
  nand2 gate1588(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate1589(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate1590(.a(G622), .O(gate207inter7));
  inv1  gate1591(.a(G632), .O(gate207inter8));
  nand2 gate1592(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate1593(.a(s_149), .b(gate207inter3), .O(gate207inter10));
  nor2  gate1594(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate1595(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate1596(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate1233(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate1234(.a(gate211inter0), .b(s_98), .O(gate211inter1));
  and2  gate1235(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate1236(.a(s_98), .O(gate211inter3));
  inv1  gate1237(.a(s_99), .O(gate211inter4));
  nand2 gate1238(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate1239(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate1240(.a(G612), .O(gate211inter7));
  inv1  gate1241(.a(G669), .O(gate211inter8));
  nand2 gate1242(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate1243(.a(s_99), .b(gate211inter3), .O(gate211inter10));
  nor2  gate1244(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate1245(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate1246(.a(gate211inter12), .b(gate211inter1), .O(G692));
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate2815(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate2816(.a(gate214inter0), .b(s_324), .O(gate214inter1));
  and2  gate2817(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate2818(.a(s_324), .O(gate214inter3));
  inv1  gate2819(.a(s_325), .O(gate214inter4));
  nand2 gate2820(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate2821(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate2822(.a(G612), .O(gate214inter7));
  inv1  gate2823(.a(G672), .O(gate214inter8));
  nand2 gate2824(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate2825(.a(s_325), .b(gate214inter3), .O(gate214inter10));
  nor2  gate2826(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate2827(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate2828(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate911(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate912(.a(gate216inter0), .b(s_52), .O(gate216inter1));
  and2  gate913(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate914(.a(s_52), .O(gate216inter3));
  inv1  gate915(.a(s_53), .O(gate216inter4));
  nand2 gate916(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate917(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate918(.a(G617), .O(gate216inter7));
  inv1  gate919(.a(G675), .O(gate216inter8));
  nand2 gate920(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate921(.a(s_53), .b(gate216inter3), .O(gate216inter10));
  nor2  gate922(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate923(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate924(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate1261(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate1262(.a(gate218inter0), .b(s_102), .O(gate218inter1));
  and2  gate1263(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate1264(.a(s_102), .O(gate218inter3));
  inv1  gate1265(.a(s_103), .O(gate218inter4));
  nand2 gate1266(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate1267(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate1268(.a(G627), .O(gate218inter7));
  inv1  gate1269(.a(G678), .O(gate218inter8));
  nand2 gate1270(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate1271(.a(s_103), .b(gate218inter3), .O(gate218inter10));
  nor2  gate1272(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate1273(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate1274(.a(gate218inter12), .b(gate218inter1), .O(G699));
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate2689(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate2690(.a(gate220inter0), .b(s_306), .O(gate220inter1));
  and2  gate2691(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate2692(.a(s_306), .O(gate220inter3));
  inv1  gate2693(.a(s_307), .O(gate220inter4));
  nand2 gate2694(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate2695(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate2696(.a(G637), .O(gate220inter7));
  inv1  gate2697(.a(G681), .O(gate220inter8));
  nand2 gate2698(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate2699(.a(s_307), .b(gate220inter3), .O(gate220inter10));
  nor2  gate2700(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate2701(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate2702(.a(gate220inter12), .b(gate220inter1), .O(G701));
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate2955(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate2956(.a(gate223inter0), .b(s_344), .O(gate223inter1));
  and2  gate2957(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate2958(.a(s_344), .O(gate223inter3));
  inv1  gate2959(.a(s_345), .O(gate223inter4));
  nand2 gate2960(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate2961(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate2962(.a(G627), .O(gate223inter7));
  inv1  gate2963(.a(G687), .O(gate223inter8));
  nand2 gate2964(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate2965(.a(s_345), .b(gate223inter3), .O(gate223inter10));
  nor2  gate2966(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate2967(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate2968(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );

  xor2  gate2465(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate2466(.a(gate225inter0), .b(s_274), .O(gate225inter1));
  and2  gate2467(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate2468(.a(s_274), .O(gate225inter3));
  inv1  gate2469(.a(s_275), .O(gate225inter4));
  nand2 gate2470(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate2471(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate2472(.a(G690), .O(gate225inter7));
  inv1  gate2473(.a(G691), .O(gate225inter8));
  nand2 gate2474(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate2475(.a(s_275), .b(gate225inter3), .O(gate225inter10));
  nor2  gate2476(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate2477(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate2478(.a(gate225inter12), .b(gate225inter1), .O(G706));
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate981(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate982(.a(gate236inter0), .b(s_62), .O(gate236inter1));
  and2  gate983(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate984(.a(s_62), .O(gate236inter3));
  inv1  gate985(.a(s_63), .O(gate236inter4));
  nand2 gate986(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate987(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate988(.a(G251), .O(gate236inter7));
  inv1  gate989(.a(G727), .O(gate236inter8));
  nand2 gate990(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate991(.a(s_63), .b(gate236inter3), .O(gate236inter10));
  nor2  gate992(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate993(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate994(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate2157(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate2158(.a(gate241inter0), .b(s_230), .O(gate241inter1));
  and2  gate2159(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate2160(.a(s_230), .O(gate241inter3));
  inv1  gate2161(.a(s_231), .O(gate241inter4));
  nand2 gate2162(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate2163(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate2164(.a(G242), .O(gate241inter7));
  inv1  gate2165(.a(G730), .O(gate241inter8));
  nand2 gate2166(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate2167(.a(s_231), .b(gate241inter3), .O(gate241inter10));
  nor2  gate2168(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate2169(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate2170(.a(gate241inter12), .b(gate241inter1), .O(G754));

  xor2  gate2409(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate2410(.a(gate242inter0), .b(s_266), .O(gate242inter1));
  and2  gate2411(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate2412(.a(s_266), .O(gate242inter3));
  inv1  gate2413(.a(s_267), .O(gate242inter4));
  nand2 gate2414(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate2415(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate2416(.a(G718), .O(gate242inter7));
  inv1  gate2417(.a(G730), .O(gate242inter8));
  nand2 gate2418(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate2419(.a(s_267), .b(gate242inter3), .O(gate242inter10));
  nor2  gate2420(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate2421(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate2422(.a(gate242inter12), .b(gate242inter1), .O(G755));

  xor2  gate855(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate856(.a(gate243inter0), .b(s_44), .O(gate243inter1));
  and2  gate857(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate858(.a(s_44), .O(gate243inter3));
  inv1  gate859(.a(s_45), .O(gate243inter4));
  nand2 gate860(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate861(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate862(.a(G245), .O(gate243inter7));
  inv1  gate863(.a(G733), .O(gate243inter8));
  nand2 gate864(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate865(.a(s_45), .b(gate243inter3), .O(gate243inter10));
  nor2  gate866(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate867(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate868(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate1947(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate1948(.a(gate249inter0), .b(s_200), .O(gate249inter1));
  and2  gate1949(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate1950(.a(s_200), .O(gate249inter3));
  inv1  gate1951(.a(s_201), .O(gate249inter4));
  nand2 gate1952(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate1953(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate1954(.a(G254), .O(gate249inter7));
  inv1  gate1955(.a(G742), .O(gate249inter8));
  nand2 gate1956(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate1957(.a(s_201), .b(gate249inter3), .O(gate249inter10));
  nor2  gate1958(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate1959(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate1960(.a(gate249inter12), .b(gate249inter1), .O(G762));

  xor2  gate2941(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate2942(.a(gate250inter0), .b(s_342), .O(gate250inter1));
  and2  gate2943(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate2944(.a(s_342), .O(gate250inter3));
  inv1  gate2945(.a(s_343), .O(gate250inter4));
  nand2 gate2946(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate2947(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate2948(.a(G706), .O(gate250inter7));
  inv1  gate2949(.a(G742), .O(gate250inter8));
  nand2 gate2950(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate2951(.a(s_343), .b(gate250inter3), .O(gate250inter10));
  nor2  gate2952(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate2953(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate2954(.a(gate250inter12), .b(gate250inter1), .O(G763));

  xor2  gate1597(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate1598(.a(gate251inter0), .b(s_150), .O(gate251inter1));
  and2  gate1599(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate1600(.a(s_150), .O(gate251inter3));
  inv1  gate1601(.a(s_151), .O(gate251inter4));
  nand2 gate1602(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate1603(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate1604(.a(G257), .O(gate251inter7));
  inv1  gate1605(.a(G745), .O(gate251inter8));
  nand2 gate1606(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate1607(.a(s_151), .b(gate251inter3), .O(gate251inter10));
  nor2  gate1608(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate1609(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate1610(.a(gate251inter12), .b(gate251inter1), .O(G764));

  xor2  gate1177(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate1178(.a(gate252inter0), .b(s_90), .O(gate252inter1));
  and2  gate1179(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate1180(.a(s_90), .O(gate252inter3));
  inv1  gate1181(.a(s_91), .O(gate252inter4));
  nand2 gate1182(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate1183(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate1184(.a(G709), .O(gate252inter7));
  inv1  gate1185(.a(G745), .O(gate252inter8));
  nand2 gate1186(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate1187(.a(s_91), .b(gate252inter3), .O(gate252inter10));
  nor2  gate1188(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate1189(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate1190(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate1191(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate1192(.a(gate255inter0), .b(s_92), .O(gate255inter1));
  and2  gate1193(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate1194(.a(s_92), .O(gate255inter3));
  inv1  gate1195(.a(s_93), .O(gate255inter4));
  nand2 gate1196(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate1197(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate1198(.a(G263), .O(gate255inter7));
  inv1  gate1199(.a(G751), .O(gate255inter8));
  nand2 gate1200(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate1201(.a(s_93), .b(gate255inter3), .O(gate255inter10));
  nor2  gate1202(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate1203(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate1204(.a(gate255inter12), .b(gate255inter1), .O(G768));

  xor2  gate883(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate884(.a(gate256inter0), .b(s_48), .O(gate256inter1));
  and2  gate885(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate886(.a(s_48), .O(gate256inter3));
  inv1  gate887(.a(s_49), .O(gate256inter4));
  nand2 gate888(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate889(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate890(.a(G715), .O(gate256inter7));
  inv1  gate891(.a(G751), .O(gate256inter8));
  nand2 gate892(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate893(.a(s_49), .b(gate256inter3), .O(gate256inter10));
  nor2  gate894(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate895(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate896(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );

  xor2  gate771(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate772(.a(gate259inter0), .b(s_32), .O(gate259inter1));
  and2  gate773(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate774(.a(s_32), .O(gate259inter3));
  inv1  gate775(.a(s_33), .O(gate259inter4));
  nand2 gate776(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate777(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate778(.a(G758), .O(gate259inter7));
  inv1  gate779(.a(G759), .O(gate259inter8));
  nand2 gate780(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate781(.a(s_33), .b(gate259inter3), .O(gate259inter10));
  nor2  gate782(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate783(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate784(.a(gate259inter12), .b(gate259inter1), .O(G776));
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate827(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate828(.a(gate261inter0), .b(s_40), .O(gate261inter1));
  and2  gate829(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate830(.a(s_40), .O(gate261inter3));
  inv1  gate831(.a(s_41), .O(gate261inter4));
  nand2 gate832(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate833(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate834(.a(G762), .O(gate261inter7));
  inv1  gate835(.a(G763), .O(gate261inter8));
  nand2 gate836(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate837(.a(s_41), .b(gate261inter3), .O(gate261inter10));
  nor2  gate838(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate839(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate840(.a(gate261inter12), .b(gate261inter1), .O(G782));
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate2353(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate2354(.a(gate263inter0), .b(s_258), .O(gate263inter1));
  and2  gate2355(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate2356(.a(s_258), .O(gate263inter3));
  inv1  gate2357(.a(s_259), .O(gate263inter4));
  nand2 gate2358(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate2359(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate2360(.a(G766), .O(gate263inter7));
  inv1  gate2361(.a(G767), .O(gate263inter8));
  nand2 gate2362(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate2363(.a(s_259), .b(gate263inter3), .O(gate263inter10));
  nor2  gate2364(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate2365(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate2366(.a(gate263inter12), .b(gate263inter1), .O(G788));

  xor2  gate2563(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate2564(.a(gate264inter0), .b(s_288), .O(gate264inter1));
  and2  gate2565(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate2566(.a(s_288), .O(gate264inter3));
  inv1  gate2567(.a(s_289), .O(gate264inter4));
  nand2 gate2568(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate2569(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate2570(.a(G768), .O(gate264inter7));
  inv1  gate2571(.a(G769), .O(gate264inter8));
  nand2 gate2572(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate2573(.a(s_289), .b(gate264inter3), .O(gate264inter10));
  nor2  gate2574(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate2575(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate2576(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate2367(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate2368(.a(gate266inter0), .b(s_260), .O(gate266inter1));
  and2  gate2369(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate2370(.a(s_260), .O(gate266inter3));
  inv1  gate2371(.a(s_261), .O(gate266inter4));
  nand2 gate2372(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate2373(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate2374(.a(G645), .O(gate266inter7));
  inv1  gate2375(.a(G773), .O(gate266inter8));
  nand2 gate2376(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate2377(.a(s_261), .b(gate266inter3), .O(gate266inter10));
  nor2  gate2378(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate2379(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate2380(.a(gate266inter12), .b(gate266inter1), .O(G797));

  xor2  gate2311(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate2312(.a(gate267inter0), .b(s_252), .O(gate267inter1));
  and2  gate2313(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate2314(.a(s_252), .O(gate267inter3));
  inv1  gate2315(.a(s_253), .O(gate267inter4));
  nand2 gate2316(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate2317(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate2318(.a(G648), .O(gate267inter7));
  inv1  gate2319(.a(G776), .O(gate267inter8));
  nand2 gate2320(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate2321(.a(s_253), .b(gate267inter3), .O(gate267inter10));
  nor2  gate2322(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate2323(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate2324(.a(gate267inter12), .b(gate267inter1), .O(G800));

  xor2  gate2675(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate2676(.a(gate268inter0), .b(s_304), .O(gate268inter1));
  and2  gate2677(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate2678(.a(s_304), .O(gate268inter3));
  inv1  gate2679(.a(s_305), .O(gate268inter4));
  nand2 gate2680(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate2681(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate2682(.a(G651), .O(gate268inter7));
  inv1  gate2683(.a(G779), .O(gate268inter8));
  nand2 gate2684(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate2685(.a(s_305), .b(gate268inter3), .O(gate268inter10));
  nor2  gate2686(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate2687(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate2688(.a(gate268inter12), .b(gate268inter1), .O(G803));

  xor2  gate1905(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate1906(.a(gate269inter0), .b(s_194), .O(gate269inter1));
  and2  gate1907(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate1908(.a(s_194), .O(gate269inter3));
  inv1  gate1909(.a(s_195), .O(gate269inter4));
  nand2 gate1910(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate1911(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate1912(.a(G654), .O(gate269inter7));
  inv1  gate1913(.a(G782), .O(gate269inter8));
  nand2 gate1914(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate1915(.a(s_195), .b(gate269inter3), .O(gate269inter10));
  nor2  gate1916(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate1917(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate1918(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate2255(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate2256(.a(gate274inter0), .b(s_244), .O(gate274inter1));
  and2  gate2257(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate2258(.a(s_244), .O(gate274inter3));
  inv1  gate2259(.a(s_245), .O(gate274inter4));
  nand2 gate2260(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate2261(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate2262(.a(G770), .O(gate274inter7));
  inv1  gate2263(.a(G794), .O(gate274inter8));
  nand2 gate2264(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate2265(.a(s_245), .b(gate274inter3), .O(gate274inter10));
  nor2  gate2266(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate2267(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate2268(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate2339(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate2340(.a(gate278inter0), .b(s_256), .O(gate278inter1));
  and2  gate2341(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate2342(.a(s_256), .O(gate278inter3));
  inv1  gate2343(.a(s_257), .O(gate278inter4));
  nand2 gate2344(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate2345(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate2346(.a(G776), .O(gate278inter7));
  inv1  gate2347(.a(G800), .O(gate278inter8));
  nand2 gate2348(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate2349(.a(s_257), .b(gate278inter3), .O(gate278inter10));
  nor2  gate2350(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate2351(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate2352(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate1989(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate1990(.a(gate282inter0), .b(s_206), .O(gate282inter1));
  and2  gate1991(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate1992(.a(s_206), .O(gate282inter3));
  inv1  gate1993(.a(s_207), .O(gate282inter4));
  nand2 gate1994(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate1995(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate1996(.a(G782), .O(gate282inter7));
  inv1  gate1997(.a(G806), .O(gate282inter8));
  nand2 gate1998(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate1999(.a(s_207), .b(gate282inter3), .O(gate282inter10));
  nor2  gate2000(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate2001(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate2002(.a(gate282inter12), .b(gate282inter1), .O(G827));

  xor2  gate1485(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate1486(.a(gate283inter0), .b(s_134), .O(gate283inter1));
  and2  gate1487(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate1488(.a(s_134), .O(gate283inter3));
  inv1  gate1489(.a(s_135), .O(gate283inter4));
  nand2 gate1490(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate1491(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate1492(.a(G657), .O(gate283inter7));
  inv1  gate1493(.a(G809), .O(gate283inter8));
  nand2 gate1494(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate1495(.a(s_135), .b(gate283inter3), .O(gate283inter10));
  nor2  gate1496(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate1497(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate1498(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate1737(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate1738(.a(gate285inter0), .b(s_170), .O(gate285inter1));
  and2  gate1739(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate1740(.a(s_170), .O(gate285inter3));
  inv1  gate1741(.a(s_171), .O(gate285inter4));
  nand2 gate1742(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate1743(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate1744(.a(G660), .O(gate285inter7));
  inv1  gate1745(.a(G812), .O(gate285inter8));
  nand2 gate1746(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate1747(.a(s_171), .b(gate285inter3), .O(gate285inter10));
  nor2  gate1748(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate1749(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate1750(.a(gate285inter12), .b(gate285inter1), .O(G830));

  xor2  gate1331(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate1332(.a(gate286inter0), .b(s_112), .O(gate286inter1));
  and2  gate1333(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate1334(.a(s_112), .O(gate286inter3));
  inv1  gate1335(.a(s_113), .O(gate286inter4));
  nand2 gate1336(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate1337(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate1338(.a(G788), .O(gate286inter7));
  inv1  gate1339(.a(G812), .O(gate286inter8));
  nand2 gate1340(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate1341(.a(s_113), .b(gate286inter3), .O(gate286inter10));
  nor2  gate1342(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate1343(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate1344(.a(gate286inter12), .b(gate286inter1), .O(G831));

  xor2  gate645(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate646(.a(gate287inter0), .b(s_14), .O(gate287inter1));
  and2  gate647(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate648(.a(s_14), .O(gate287inter3));
  inv1  gate649(.a(s_15), .O(gate287inter4));
  nand2 gate650(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate651(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate652(.a(G663), .O(gate287inter7));
  inv1  gate653(.a(G815), .O(gate287inter8));
  nand2 gate654(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate655(.a(s_15), .b(gate287inter3), .O(gate287inter10));
  nor2  gate656(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate657(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate658(.a(gate287inter12), .b(gate287inter1), .O(G832));

  xor2  gate659(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate660(.a(gate288inter0), .b(s_16), .O(gate288inter1));
  and2  gate661(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate662(.a(s_16), .O(gate288inter3));
  inv1  gate663(.a(s_17), .O(gate288inter4));
  nand2 gate664(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate665(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate666(.a(G791), .O(gate288inter7));
  inv1  gate667(.a(G815), .O(gate288inter8));
  nand2 gate668(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate669(.a(s_17), .b(gate288inter3), .O(gate288inter10));
  nor2  gate670(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate671(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate672(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate1373(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate1374(.a(gate291inter0), .b(s_118), .O(gate291inter1));
  and2  gate1375(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate1376(.a(s_118), .O(gate291inter3));
  inv1  gate1377(.a(s_119), .O(gate291inter4));
  nand2 gate1378(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate1379(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate1380(.a(G822), .O(gate291inter7));
  inv1  gate1381(.a(G823), .O(gate291inter8));
  nand2 gate1382(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate1383(.a(s_119), .b(gate291inter3), .O(gate291inter10));
  nor2  gate1384(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate1385(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate1386(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate1961(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate1962(.a(gate295inter0), .b(s_202), .O(gate295inter1));
  and2  gate1963(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate1964(.a(s_202), .O(gate295inter3));
  inv1  gate1965(.a(s_203), .O(gate295inter4));
  nand2 gate1966(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate1967(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate1968(.a(G830), .O(gate295inter7));
  inv1  gate1969(.a(G831), .O(gate295inter8));
  nand2 gate1970(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate1971(.a(s_203), .b(gate295inter3), .O(gate295inter10));
  nor2  gate1972(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate1973(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate1974(.a(gate295inter12), .b(gate295inter1), .O(G912));

  xor2  gate1835(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate1836(.a(gate296inter0), .b(s_184), .O(gate296inter1));
  and2  gate1837(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate1838(.a(s_184), .O(gate296inter3));
  inv1  gate1839(.a(s_185), .O(gate296inter4));
  nand2 gate1840(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate1841(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate1842(.a(G826), .O(gate296inter7));
  inv1  gate1843(.a(G827), .O(gate296inter8));
  nand2 gate1844(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate1845(.a(s_185), .b(gate296inter3), .O(gate296inter10));
  nor2  gate1846(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate1847(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate1848(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate2017(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate2018(.a(gate389inter0), .b(s_210), .O(gate389inter1));
  and2  gate2019(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate2020(.a(s_210), .O(gate389inter3));
  inv1  gate2021(.a(s_211), .O(gate389inter4));
  nand2 gate2022(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate2023(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate2024(.a(G3), .O(gate389inter7));
  inv1  gate2025(.a(G1042), .O(gate389inter8));
  nand2 gate2026(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate2027(.a(s_211), .b(gate389inter3), .O(gate389inter10));
  nor2  gate2028(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate2029(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate2030(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate2269(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate2270(.a(gate391inter0), .b(s_246), .O(gate391inter1));
  and2  gate2271(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate2272(.a(s_246), .O(gate391inter3));
  inv1  gate2273(.a(s_247), .O(gate391inter4));
  nand2 gate2274(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate2275(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate2276(.a(G5), .O(gate391inter7));
  inv1  gate2277(.a(G1048), .O(gate391inter8));
  nand2 gate2278(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate2279(.a(s_247), .b(gate391inter3), .O(gate391inter10));
  nor2  gate2280(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate2281(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate2282(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate1611(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate1612(.a(gate394inter0), .b(s_152), .O(gate394inter1));
  and2  gate1613(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate1614(.a(s_152), .O(gate394inter3));
  inv1  gate1615(.a(s_153), .O(gate394inter4));
  nand2 gate1616(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate1617(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate1618(.a(G8), .O(gate394inter7));
  inv1  gate1619(.a(G1057), .O(gate394inter8));
  nand2 gate1620(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate1621(.a(s_153), .b(gate394inter3), .O(gate394inter10));
  nor2  gate1622(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate1623(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate1624(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );

  xor2  gate1443(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate1444(.a(gate396inter0), .b(s_128), .O(gate396inter1));
  and2  gate1445(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate1446(.a(s_128), .O(gate396inter3));
  inv1  gate1447(.a(s_129), .O(gate396inter4));
  nand2 gate1448(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate1449(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate1450(.a(G10), .O(gate396inter7));
  inv1  gate1451(.a(G1063), .O(gate396inter8));
  nand2 gate1452(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate1453(.a(s_129), .b(gate396inter3), .O(gate396inter10));
  nor2  gate1454(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate1455(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate1456(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate1359(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate1360(.a(gate398inter0), .b(s_116), .O(gate398inter1));
  and2  gate1361(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate1362(.a(s_116), .O(gate398inter3));
  inv1  gate1363(.a(s_117), .O(gate398inter4));
  nand2 gate1364(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate1365(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate1366(.a(G12), .O(gate398inter7));
  inv1  gate1367(.a(G1069), .O(gate398inter8));
  nand2 gate1368(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate1369(.a(s_117), .b(gate398inter3), .O(gate398inter10));
  nor2  gate1370(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate1371(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate1372(.a(gate398inter12), .b(gate398inter1), .O(G1165));

  xor2  gate1023(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate1024(.a(gate399inter0), .b(s_68), .O(gate399inter1));
  and2  gate1025(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate1026(.a(s_68), .O(gate399inter3));
  inv1  gate1027(.a(s_69), .O(gate399inter4));
  nand2 gate1028(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate1029(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate1030(.a(G13), .O(gate399inter7));
  inv1  gate1031(.a(G1072), .O(gate399inter8));
  nand2 gate1032(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate1033(.a(s_69), .b(gate399inter3), .O(gate399inter10));
  nor2  gate1034(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate1035(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate1036(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate1079(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate1080(.a(gate403inter0), .b(s_76), .O(gate403inter1));
  and2  gate1081(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate1082(.a(s_76), .O(gate403inter3));
  inv1  gate1083(.a(s_77), .O(gate403inter4));
  nand2 gate1084(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate1085(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate1086(.a(G17), .O(gate403inter7));
  inv1  gate1087(.a(G1084), .O(gate403inter8));
  nand2 gate1088(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate1089(.a(s_77), .b(gate403inter3), .O(gate403inter10));
  nor2  gate1090(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate1091(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate1092(.a(gate403inter12), .b(gate403inter1), .O(G1180));
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate2899(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate2900(.a(gate407inter0), .b(s_336), .O(gate407inter1));
  and2  gate2901(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate2902(.a(s_336), .O(gate407inter3));
  inv1  gate2903(.a(s_337), .O(gate407inter4));
  nand2 gate2904(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate2905(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate2906(.a(G21), .O(gate407inter7));
  inv1  gate2907(.a(G1096), .O(gate407inter8));
  nand2 gate2908(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate2909(.a(s_337), .b(gate407inter3), .O(gate407inter10));
  nor2  gate2910(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate2911(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate2912(.a(gate407inter12), .b(gate407inter1), .O(G1192));

  xor2  gate2087(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate2088(.a(gate408inter0), .b(s_220), .O(gate408inter1));
  and2  gate2089(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate2090(.a(s_220), .O(gate408inter3));
  inv1  gate2091(.a(s_221), .O(gate408inter4));
  nand2 gate2092(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate2093(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate2094(.a(G22), .O(gate408inter7));
  inv1  gate2095(.a(G1099), .O(gate408inter8));
  nand2 gate2096(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate2097(.a(s_221), .b(gate408inter3), .O(gate408inter10));
  nor2  gate2098(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate2099(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate2100(.a(gate408inter12), .b(gate408inter1), .O(G1195));

  xor2  gate1317(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate1318(.a(gate409inter0), .b(s_110), .O(gate409inter1));
  and2  gate1319(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate1320(.a(s_110), .O(gate409inter3));
  inv1  gate1321(.a(s_111), .O(gate409inter4));
  nand2 gate1322(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate1323(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate1324(.a(G23), .O(gate409inter7));
  inv1  gate1325(.a(G1102), .O(gate409inter8));
  nand2 gate1326(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate1327(.a(s_111), .b(gate409inter3), .O(gate409inter10));
  nor2  gate1328(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate1329(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate1330(.a(gate409inter12), .b(gate409inter1), .O(G1198));

  xor2  gate1919(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate1920(.a(gate410inter0), .b(s_196), .O(gate410inter1));
  and2  gate1921(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate1922(.a(s_196), .O(gate410inter3));
  inv1  gate1923(.a(s_197), .O(gate410inter4));
  nand2 gate1924(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate1925(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate1926(.a(G24), .O(gate410inter7));
  inv1  gate1927(.a(G1105), .O(gate410inter8));
  nand2 gate1928(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate1929(.a(s_197), .b(gate410inter3), .O(gate410inter10));
  nor2  gate1930(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate1931(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate1932(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );

  xor2  gate2913(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate2914(.a(gate412inter0), .b(s_338), .O(gate412inter1));
  and2  gate2915(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate2916(.a(s_338), .O(gate412inter3));
  inv1  gate2917(.a(s_339), .O(gate412inter4));
  nand2 gate2918(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate2919(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate2920(.a(G26), .O(gate412inter7));
  inv1  gate2921(.a(G1111), .O(gate412inter8));
  nand2 gate2922(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate2923(.a(s_339), .b(gate412inter3), .O(gate412inter10));
  nor2  gate2924(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate2925(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate2926(.a(gate412inter12), .b(gate412inter1), .O(G1207));

  xor2  gate2927(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate2928(.a(gate413inter0), .b(s_340), .O(gate413inter1));
  and2  gate2929(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate2930(.a(s_340), .O(gate413inter3));
  inv1  gate2931(.a(s_341), .O(gate413inter4));
  nand2 gate2932(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate2933(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate2934(.a(G27), .O(gate413inter7));
  inv1  gate2935(.a(G1114), .O(gate413inter8));
  nand2 gate2936(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate2937(.a(s_341), .b(gate413inter3), .O(gate413inter10));
  nor2  gate2938(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate2939(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate2940(.a(gate413inter12), .b(gate413inter1), .O(G1210));

  xor2  gate2451(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate2452(.a(gate414inter0), .b(s_272), .O(gate414inter1));
  and2  gate2453(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate2454(.a(s_272), .O(gate414inter3));
  inv1  gate2455(.a(s_273), .O(gate414inter4));
  nand2 gate2456(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate2457(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate2458(.a(G28), .O(gate414inter7));
  inv1  gate2459(.a(G1117), .O(gate414inter8));
  nand2 gate2460(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate2461(.a(s_273), .b(gate414inter3), .O(gate414inter10));
  nor2  gate2462(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate2463(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate2464(.a(gate414inter12), .b(gate414inter1), .O(G1213));

  xor2  gate897(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate898(.a(gate415inter0), .b(s_50), .O(gate415inter1));
  and2  gate899(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate900(.a(s_50), .O(gate415inter3));
  inv1  gate901(.a(s_51), .O(gate415inter4));
  nand2 gate902(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate903(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate904(.a(G29), .O(gate415inter7));
  inv1  gate905(.a(G1120), .O(gate415inter8));
  nand2 gate906(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate907(.a(s_51), .b(gate415inter3), .O(gate415inter10));
  nor2  gate908(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate909(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate910(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate2003(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate2004(.a(gate421inter0), .b(s_208), .O(gate421inter1));
  and2  gate2005(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate2006(.a(s_208), .O(gate421inter3));
  inv1  gate2007(.a(s_209), .O(gate421inter4));
  nand2 gate2008(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate2009(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate2010(.a(G2), .O(gate421inter7));
  inv1  gate2011(.a(G1135), .O(gate421inter8));
  nand2 gate2012(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate2013(.a(s_209), .b(gate421inter3), .O(gate421inter10));
  nor2  gate2014(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate2015(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate2016(.a(gate421inter12), .b(gate421inter1), .O(G1230));

  xor2  gate575(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate576(.a(gate422inter0), .b(s_4), .O(gate422inter1));
  and2  gate577(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate578(.a(s_4), .O(gate422inter3));
  inv1  gate579(.a(s_5), .O(gate422inter4));
  nand2 gate580(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate581(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate582(.a(G1039), .O(gate422inter7));
  inv1  gate583(.a(G1135), .O(gate422inter8));
  nand2 gate584(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate585(.a(s_5), .b(gate422inter3), .O(gate422inter10));
  nor2  gate586(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate587(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate588(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );

  xor2  gate1569(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate1570(.a(gate424inter0), .b(s_146), .O(gate424inter1));
  and2  gate1571(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate1572(.a(s_146), .O(gate424inter3));
  inv1  gate1573(.a(s_147), .O(gate424inter4));
  nand2 gate1574(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate1575(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate1576(.a(G1042), .O(gate424inter7));
  inv1  gate1577(.a(G1138), .O(gate424inter8));
  nand2 gate1578(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate1579(.a(s_147), .b(gate424inter3), .O(gate424inter10));
  nor2  gate1580(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate1581(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate1582(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate2703(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate2704(.a(gate430inter0), .b(s_308), .O(gate430inter1));
  and2  gate2705(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate2706(.a(s_308), .O(gate430inter3));
  inv1  gate2707(.a(s_309), .O(gate430inter4));
  nand2 gate2708(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate2709(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate2710(.a(G1051), .O(gate430inter7));
  inv1  gate2711(.a(G1147), .O(gate430inter8));
  nand2 gate2712(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate2713(.a(s_309), .b(gate430inter3), .O(gate430inter10));
  nor2  gate2714(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate2715(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate2716(.a(gate430inter12), .b(gate430inter1), .O(G1239));
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );

  xor2  gate1247(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate1248(.a(gate432inter0), .b(s_100), .O(gate432inter1));
  and2  gate1249(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate1250(.a(s_100), .O(gate432inter3));
  inv1  gate1251(.a(s_101), .O(gate432inter4));
  nand2 gate1252(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate1253(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate1254(.a(G1054), .O(gate432inter7));
  inv1  gate1255(.a(G1150), .O(gate432inter8));
  nand2 gate1256(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate1257(.a(s_101), .b(gate432inter3), .O(gate432inter10));
  nor2  gate1258(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate1259(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate1260(.a(gate432inter12), .b(gate432inter1), .O(G1241));
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate995(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate996(.a(gate434inter0), .b(s_64), .O(gate434inter1));
  and2  gate997(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate998(.a(s_64), .O(gate434inter3));
  inv1  gate999(.a(s_65), .O(gate434inter4));
  nand2 gate1000(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate1001(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate1002(.a(G1057), .O(gate434inter7));
  inv1  gate1003(.a(G1153), .O(gate434inter8));
  nand2 gate1004(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate1005(.a(s_65), .b(gate434inter3), .O(gate434inter10));
  nor2  gate1006(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate1007(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate1008(.a(gate434inter12), .b(gate434inter1), .O(G1243));
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate1457(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate1458(.a(gate437inter0), .b(s_130), .O(gate437inter1));
  and2  gate1459(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate1460(.a(s_130), .O(gate437inter3));
  inv1  gate1461(.a(s_131), .O(gate437inter4));
  nand2 gate1462(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate1463(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate1464(.a(G10), .O(gate437inter7));
  inv1  gate1465(.a(G1159), .O(gate437inter8));
  nand2 gate1466(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate1467(.a(s_131), .b(gate437inter3), .O(gate437inter10));
  nor2  gate1468(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate1469(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate1470(.a(gate437inter12), .b(gate437inter1), .O(G1246));

  xor2  gate631(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate632(.a(gate438inter0), .b(s_12), .O(gate438inter1));
  and2  gate633(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate634(.a(s_12), .O(gate438inter3));
  inv1  gate635(.a(s_13), .O(gate438inter4));
  nand2 gate636(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate637(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate638(.a(G1063), .O(gate438inter7));
  inv1  gate639(.a(G1159), .O(gate438inter8));
  nand2 gate640(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate641(.a(s_13), .b(gate438inter3), .O(gate438inter10));
  nor2  gate642(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate643(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate644(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );

  xor2  gate1709(.a(G1174), .b(G15), .O(gate447inter0));
  nand2 gate1710(.a(gate447inter0), .b(s_166), .O(gate447inter1));
  and2  gate1711(.a(G1174), .b(G15), .O(gate447inter2));
  inv1  gate1712(.a(s_166), .O(gate447inter3));
  inv1  gate1713(.a(s_167), .O(gate447inter4));
  nand2 gate1714(.a(gate447inter4), .b(gate447inter3), .O(gate447inter5));
  nor2  gate1715(.a(gate447inter5), .b(gate447inter2), .O(gate447inter6));
  inv1  gate1716(.a(G15), .O(gate447inter7));
  inv1  gate1717(.a(G1174), .O(gate447inter8));
  nand2 gate1718(.a(gate447inter8), .b(gate447inter7), .O(gate447inter9));
  nand2 gate1719(.a(s_167), .b(gate447inter3), .O(gate447inter10));
  nor2  gate1720(.a(gate447inter10), .b(gate447inter9), .O(gate447inter11));
  nor2  gate1721(.a(gate447inter11), .b(gate447inter6), .O(gate447inter12));
  nand2 gate1722(.a(gate447inter12), .b(gate447inter1), .O(G1256));
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );

  xor2  gate1401(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate1402(.a(gate449inter0), .b(s_122), .O(gate449inter1));
  and2  gate1403(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate1404(.a(s_122), .O(gate449inter3));
  inv1  gate1405(.a(s_123), .O(gate449inter4));
  nand2 gate1406(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate1407(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate1408(.a(G16), .O(gate449inter7));
  inv1  gate1409(.a(G1177), .O(gate449inter8));
  nand2 gate1410(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate1411(.a(s_123), .b(gate449inter3), .O(gate449inter10));
  nor2  gate1412(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate1413(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate1414(.a(gate449inter12), .b(gate449inter1), .O(G1258));

  xor2  gate2171(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate2172(.a(gate450inter0), .b(s_232), .O(gate450inter1));
  and2  gate2173(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate2174(.a(s_232), .O(gate450inter3));
  inv1  gate2175(.a(s_233), .O(gate450inter4));
  nand2 gate2176(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate2177(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate2178(.a(G1081), .O(gate450inter7));
  inv1  gate2179(.a(G1177), .O(gate450inter8));
  nand2 gate2180(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate2181(.a(s_233), .b(gate450inter3), .O(gate450inter10));
  nor2  gate2182(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate2183(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate2184(.a(gate450inter12), .b(gate450inter1), .O(G1259));
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );

  xor2  gate1751(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate1752(.a(gate455inter0), .b(s_172), .O(gate455inter1));
  and2  gate1753(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate1754(.a(s_172), .O(gate455inter3));
  inv1  gate1755(.a(s_173), .O(gate455inter4));
  nand2 gate1756(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate1757(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate1758(.a(G19), .O(gate455inter7));
  inv1  gate1759(.a(G1186), .O(gate455inter8));
  nand2 gate1760(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate1761(.a(s_173), .b(gate455inter3), .O(gate455inter10));
  nor2  gate1762(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate1763(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate1764(.a(gate455inter12), .b(gate455inter1), .O(G1264));

  xor2  gate2185(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate2186(.a(gate456inter0), .b(s_234), .O(gate456inter1));
  and2  gate2187(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate2188(.a(s_234), .O(gate456inter3));
  inv1  gate2189(.a(s_235), .O(gate456inter4));
  nand2 gate2190(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate2191(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate2192(.a(G1090), .O(gate456inter7));
  inv1  gate2193(.a(G1186), .O(gate456inter8));
  nand2 gate2194(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate2195(.a(s_235), .b(gate456inter3), .O(gate456inter10));
  nor2  gate2196(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate2197(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate2198(.a(gate456inter12), .b(gate456inter1), .O(G1265));
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );

  xor2  gate2591(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate2592(.a(gate458inter0), .b(s_292), .O(gate458inter1));
  and2  gate2593(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate2594(.a(s_292), .O(gate458inter3));
  inv1  gate2595(.a(s_293), .O(gate458inter4));
  nand2 gate2596(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate2597(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate2598(.a(G1093), .O(gate458inter7));
  inv1  gate2599(.a(G1189), .O(gate458inter8));
  nand2 gate2600(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate2601(.a(s_293), .b(gate458inter3), .O(gate458inter10));
  nor2  gate2602(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate2603(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate2604(.a(gate458inter12), .b(gate458inter1), .O(G1267));

  xor2  gate1499(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate1500(.a(gate459inter0), .b(s_136), .O(gate459inter1));
  and2  gate1501(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate1502(.a(s_136), .O(gate459inter3));
  inv1  gate1503(.a(s_137), .O(gate459inter4));
  nand2 gate1504(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate1505(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate1506(.a(G21), .O(gate459inter7));
  inv1  gate1507(.a(G1192), .O(gate459inter8));
  nand2 gate1508(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate1509(.a(s_137), .b(gate459inter3), .O(gate459inter10));
  nor2  gate1510(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate1511(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate1512(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate2647(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate2648(.a(gate461inter0), .b(s_300), .O(gate461inter1));
  and2  gate2649(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate2650(.a(s_300), .O(gate461inter3));
  inv1  gate2651(.a(s_301), .O(gate461inter4));
  nand2 gate2652(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate2653(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate2654(.a(G22), .O(gate461inter7));
  inv1  gate2655(.a(G1195), .O(gate461inter8));
  nand2 gate2656(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate2657(.a(s_301), .b(gate461inter3), .O(gate461inter10));
  nor2  gate2658(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate2659(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate2660(.a(gate461inter12), .b(gate461inter1), .O(G1270));
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );

  xor2  gate1037(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate1038(.a(gate469inter0), .b(s_70), .O(gate469inter1));
  and2  gate1039(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate1040(.a(s_70), .O(gate469inter3));
  inv1  gate1041(.a(s_71), .O(gate469inter4));
  nand2 gate1042(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate1043(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate1044(.a(G26), .O(gate469inter7));
  inv1  gate1045(.a(G1207), .O(gate469inter8));
  nand2 gate1046(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate1047(.a(s_71), .b(gate469inter3), .O(gate469inter10));
  nor2  gate1048(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate1049(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate1050(.a(gate469inter12), .b(gate469inter1), .O(G1278));
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate589(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate590(.a(gate471inter0), .b(s_6), .O(gate471inter1));
  and2  gate591(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate592(.a(s_6), .O(gate471inter3));
  inv1  gate593(.a(s_7), .O(gate471inter4));
  nand2 gate594(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate595(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate596(.a(G27), .O(gate471inter7));
  inv1  gate597(.a(G1210), .O(gate471inter8));
  nand2 gate598(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate599(.a(s_7), .b(gate471inter3), .O(gate471inter10));
  nor2  gate600(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate601(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate602(.a(gate471inter12), .b(gate471inter1), .O(G1280));

  xor2  gate2535(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate2536(.a(gate472inter0), .b(s_284), .O(gate472inter1));
  and2  gate2537(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate2538(.a(s_284), .O(gate472inter3));
  inv1  gate2539(.a(s_285), .O(gate472inter4));
  nand2 gate2540(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate2541(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate2542(.a(G1114), .O(gate472inter7));
  inv1  gate2543(.a(G1210), .O(gate472inter8));
  nand2 gate2544(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate2545(.a(s_285), .b(gate472inter3), .O(gate472inter10));
  nor2  gate2546(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate2547(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate2548(.a(gate472inter12), .b(gate472inter1), .O(G1281));

  xor2  gate1219(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate1220(.a(gate473inter0), .b(s_96), .O(gate473inter1));
  and2  gate1221(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate1222(.a(s_96), .O(gate473inter3));
  inv1  gate1223(.a(s_97), .O(gate473inter4));
  nand2 gate1224(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate1225(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate1226(.a(G28), .O(gate473inter7));
  inv1  gate1227(.a(G1213), .O(gate473inter8));
  nand2 gate1228(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate1229(.a(s_97), .b(gate473inter3), .O(gate473inter10));
  nor2  gate1230(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate1231(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate1232(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate2787(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate2788(.a(gate475inter0), .b(s_320), .O(gate475inter1));
  and2  gate2789(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate2790(.a(s_320), .O(gate475inter3));
  inv1  gate2791(.a(s_321), .O(gate475inter4));
  nand2 gate2792(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate2793(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate2794(.a(G29), .O(gate475inter7));
  inv1  gate2795(.a(G1216), .O(gate475inter8));
  nand2 gate2796(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate2797(.a(s_321), .b(gate475inter3), .O(gate475inter10));
  nor2  gate2798(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate2799(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate2800(.a(gate475inter12), .b(gate475inter1), .O(G1284));
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );

  xor2  gate2605(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate2606(.a(gate483inter0), .b(s_294), .O(gate483inter1));
  and2  gate2607(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate2608(.a(s_294), .O(gate483inter3));
  inv1  gate2609(.a(s_295), .O(gate483inter4));
  nand2 gate2610(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate2611(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate2612(.a(G1228), .O(gate483inter7));
  inv1  gate2613(.a(G1229), .O(gate483inter8));
  nand2 gate2614(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate2615(.a(s_295), .b(gate483inter3), .O(gate483inter10));
  nor2  gate2616(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate2617(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate2618(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate743(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate744(.a(gate485inter0), .b(s_28), .O(gate485inter1));
  and2  gate745(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate746(.a(s_28), .O(gate485inter3));
  inv1  gate747(.a(s_29), .O(gate485inter4));
  nand2 gate748(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate749(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate750(.a(G1232), .O(gate485inter7));
  inv1  gate751(.a(G1233), .O(gate485inter8));
  nand2 gate752(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate753(.a(s_29), .b(gate485inter3), .O(gate485inter10));
  nor2  gate754(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate755(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate756(.a(gate485inter12), .b(gate485inter1), .O(G1294));

  xor2  gate1163(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate1164(.a(gate486inter0), .b(s_88), .O(gate486inter1));
  and2  gate1165(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate1166(.a(s_88), .O(gate486inter3));
  inv1  gate1167(.a(s_89), .O(gate486inter4));
  nand2 gate1168(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate1169(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate1170(.a(G1234), .O(gate486inter7));
  inv1  gate1171(.a(G1235), .O(gate486inter8));
  nand2 gate1172(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate1173(.a(s_89), .b(gate486inter3), .O(gate486inter10));
  nor2  gate1174(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate1175(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate1176(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate1527(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate1528(.a(gate488inter0), .b(s_140), .O(gate488inter1));
  and2  gate1529(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate1530(.a(s_140), .O(gate488inter3));
  inv1  gate1531(.a(s_141), .O(gate488inter4));
  nand2 gate1532(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate1533(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate1534(.a(G1238), .O(gate488inter7));
  inv1  gate1535(.a(G1239), .O(gate488inter8));
  nand2 gate1536(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate1537(.a(s_141), .b(gate488inter3), .O(gate488inter10));
  nor2  gate1538(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate1539(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate1540(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate2059(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate2060(.a(gate490inter0), .b(s_216), .O(gate490inter1));
  and2  gate2061(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate2062(.a(s_216), .O(gate490inter3));
  inv1  gate2063(.a(s_217), .O(gate490inter4));
  nand2 gate2064(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate2065(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate2066(.a(G1242), .O(gate490inter7));
  inv1  gate2067(.a(G1243), .O(gate490inter8));
  nand2 gate2068(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate2069(.a(s_217), .b(gate490inter3), .O(gate490inter10));
  nor2  gate2070(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate2071(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate2072(.a(gate490inter12), .b(gate490inter1), .O(G1299));

  xor2  gate1513(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate1514(.a(gate491inter0), .b(s_138), .O(gate491inter1));
  and2  gate1515(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate1516(.a(s_138), .O(gate491inter3));
  inv1  gate1517(.a(s_139), .O(gate491inter4));
  nand2 gate1518(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate1519(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate1520(.a(G1244), .O(gate491inter7));
  inv1  gate1521(.a(G1245), .O(gate491inter8));
  nand2 gate1522(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate1523(.a(s_139), .b(gate491inter3), .O(gate491inter10));
  nor2  gate1524(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate1525(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate1526(.a(gate491inter12), .b(gate491inter1), .O(G1300));

  xor2  gate1429(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate1430(.a(gate492inter0), .b(s_126), .O(gate492inter1));
  and2  gate1431(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate1432(.a(s_126), .O(gate492inter3));
  inv1  gate1433(.a(s_127), .O(gate492inter4));
  nand2 gate1434(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate1435(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate1436(.a(G1246), .O(gate492inter7));
  inv1  gate1437(.a(G1247), .O(gate492inter8));
  nand2 gate1438(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate1439(.a(s_127), .b(gate492inter3), .O(gate492inter10));
  nor2  gate1440(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate1441(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate1442(.a(gate492inter12), .b(gate492inter1), .O(G1301));

  xor2  gate2619(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate2620(.a(gate493inter0), .b(s_296), .O(gate493inter1));
  and2  gate2621(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate2622(.a(s_296), .O(gate493inter3));
  inv1  gate2623(.a(s_297), .O(gate493inter4));
  nand2 gate2624(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate2625(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate2626(.a(G1248), .O(gate493inter7));
  inv1  gate2627(.a(G1249), .O(gate493inter8));
  nand2 gate2628(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate2629(.a(s_297), .b(gate493inter3), .O(gate493inter10));
  nor2  gate2630(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate2631(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate2632(.a(gate493inter12), .b(gate493inter1), .O(G1302));
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );

  xor2  gate2143(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate2144(.a(gate498inter0), .b(s_228), .O(gate498inter1));
  and2  gate2145(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate2146(.a(s_228), .O(gate498inter3));
  inv1  gate2147(.a(s_229), .O(gate498inter4));
  nand2 gate2148(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate2149(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate2150(.a(G1258), .O(gate498inter7));
  inv1  gate2151(.a(G1259), .O(gate498inter8));
  nand2 gate2152(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate2153(.a(s_229), .b(gate498inter3), .O(gate498inter10));
  nor2  gate2154(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate2155(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate2156(.a(gate498inter12), .b(gate498inter1), .O(G1307));

  xor2  gate1009(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate1010(.a(gate499inter0), .b(s_66), .O(gate499inter1));
  and2  gate1011(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate1012(.a(s_66), .O(gate499inter3));
  inv1  gate1013(.a(s_67), .O(gate499inter4));
  nand2 gate1014(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate1015(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate1016(.a(G1260), .O(gate499inter7));
  inv1  gate1017(.a(G1261), .O(gate499inter8));
  nand2 gate1018(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate1019(.a(s_67), .b(gate499inter3), .O(gate499inter10));
  nor2  gate1020(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate1021(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate1022(.a(gate499inter12), .b(gate499inter1), .O(G1308));
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate1849(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate1850(.a(gate503inter0), .b(s_186), .O(gate503inter1));
  and2  gate1851(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate1852(.a(s_186), .O(gate503inter3));
  inv1  gate1853(.a(s_187), .O(gate503inter4));
  nand2 gate1854(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate1855(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate1856(.a(G1268), .O(gate503inter7));
  inv1  gate1857(.a(G1269), .O(gate503inter8));
  nand2 gate1858(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate1859(.a(s_187), .b(gate503inter3), .O(gate503inter10));
  nor2  gate1860(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate1861(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate1862(.a(gate503inter12), .b(gate503inter1), .O(G1312));

  xor2  gate2521(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate2522(.a(gate504inter0), .b(s_282), .O(gate504inter1));
  and2  gate2523(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate2524(.a(s_282), .O(gate504inter3));
  inv1  gate2525(.a(s_283), .O(gate504inter4));
  nand2 gate2526(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate2527(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate2528(.a(G1270), .O(gate504inter7));
  inv1  gate2529(.a(G1271), .O(gate504inter8));
  nand2 gate2530(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate2531(.a(s_283), .b(gate504inter3), .O(gate504inter10));
  nor2  gate2532(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate2533(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate2534(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate1793(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate1794(.a(gate506inter0), .b(s_178), .O(gate506inter1));
  and2  gate1795(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate1796(.a(s_178), .O(gate506inter3));
  inv1  gate1797(.a(s_179), .O(gate506inter4));
  nand2 gate1798(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate1799(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate1800(.a(G1274), .O(gate506inter7));
  inv1  gate1801(.a(G1275), .O(gate506inter8));
  nand2 gate1802(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate1803(.a(s_179), .b(gate506inter3), .O(gate506inter10));
  nor2  gate1804(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate1805(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate1806(.a(gate506inter12), .b(gate506inter1), .O(G1315));

  xor2  gate1065(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate1066(.a(gate507inter0), .b(s_74), .O(gate507inter1));
  and2  gate1067(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate1068(.a(s_74), .O(gate507inter3));
  inv1  gate1069(.a(s_75), .O(gate507inter4));
  nand2 gate1070(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate1071(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate1072(.a(G1276), .O(gate507inter7));
  inv1  gate1073(.a(G1277), .O(gate507inter8));
  nand2 gate1074(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate1075(.a(s_75), .b(gate507inter3), .O(gate507inter10));
  nor2  gate1076(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate1077(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate1078(.a(gate507inter12), .b(gate507inter1), .O(G1316));

  xor2  gate2381(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate2382(.a(gate508inter0), .b(s_262), .O(gate508inter1));
  and2  gate2383(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate2384(.a(s_262), .O(gate508inter3));
  inv1  gate2385(.a(s_263), .O(gate508inter4));
  nand2 gate2386(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate2387(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate2388(.a(G1278), .O(gate508inter7));
  inv1  gate2389(.a(G1279), .O(gate508inter8));
  nand2 gate2390(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate2391(.a(s_263), .b(gate508inter3), .O(gate508inter10));
  nor2  gate2392(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate2393(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate2394(.a(gate508inter12), .b(gate508inter1), .O(G1317));

  xor2  gate2801(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate2802(.a(gate509inter0), .b(s_322), .O(gate509inter1));
  and2  gate2803(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate2804(.a(s_322), .O(gate509inter3));
  inv1  gate2805(.a(s_323), .O(gate509inter4));
  nand2 gate2806(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate2807(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate2808(.a(G1280), .O(gate509inter7));
  inv1  gate2809(.a(G1281), .O(gate509inter8));
  nand2 gate2810(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate2811(.a(s_323), .b(gate509inter3), .O(gate509inter10));
  nor2  gate2812(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate2813(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate2814(.a(gate509inter12), .b(gate509inter1), .O(G1318));

  xor2  gate1863(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate1864(.a(gate510inter0), .b(s_188), .O(gate510inter1));
  and2  gate1865(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate1866(.a(s_188), .O(gate510inter3));
  inv1  gate1867(.a(s_189), .O(gate510inter4));
  nand2 gate1868(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate1869(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate1870(.a(G1282), .O(gate510inter7));
  inv1  gate1871(.a(G1283), .O(gate510inter8));
  nand2 gate1872(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate1873(.a(s_189), .b(gate510inter3), .O(gate510inter10));
  nor2  gate1874(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate1875(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate1876(.a(gate510inter12), .b(gate510inter1), .O(G1319));

  xor2  gate1891(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate1892(.a(gate511inter0), .b(s_192), .O(gate511inter1));
  and2  gate1893(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate1894(.a(s_192), .O(gate511inter3));
  inv1  gate1895(.a(s_193), .O(gate511inter4));
  nand2 gate1896(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate1897(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate1898(.a(G1284), .O(gate511inter7));
  inv1  gate1899(.a(G1285), .O(gate511inter8));
  nand2 gate1900(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate1901(.a(s_193), .b(gate511inter3), .O(gate511inter10));
  nor2  gate1902(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate1903(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate1904(.a(gate511inter12), .b(gate511inter1), .O(G1320));

  xor2  gate869(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate870(.a(gate512inter0), .b(s_46), .O(gate512inter1));
  and2  gate871(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate872(.a(s_46), .O(gate512inter3));
  inv1  gate873(.a(s_47), .O(gate512inter4));
  nand2 gate874(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate875(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate876(.a(G1286), .O(gate512inter7));
  inv1  gate877(.a(G1287), .O(gate512inter8));
  nand2 gate878(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate879(.a(s_47), .b(gate512inter3), .O(gate512inter10));
  nor2  gate880(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate881(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate882(.a(gate512inter12), .b(gate512inter1), .O(G1321));

  xor2  gate2101(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate2102(.a(gate513inter0), .b(s_222), .O(gate513inter1));
  and2  gate2103(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate2104(.a(s_222), .O(gate513inter3));
  inv1  gate2105(.a(s_223), .O(gate513inter4));
  nand2 gate2106(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate2107(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate2108(.a(G1288), .O(gate513inter7));
  inv1  gate2109(.a(G1289), .O(gate513inter8));
  nand2 gate2110(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate2111(.a(s_223), .b(gate513inter3), .O(gate513inter10));
  nor2  gate2112(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate2113(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate2114(.a(gate513inter12), .b(gate513inter1), .O(G1322));

  xor2  gate1821(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate1822(.a(gate514inter0), .b(s_182), .O(gate514inter1));
  and2  gate1823(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate1824(.a(s_182), .O(gate514inter3));
  inv1  gate1825(.a(s_183), .O(gate514inter4));
  nand2 gate1826(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate1827(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate1828(.a(G1290), .O(gate514inter7));
  inv1  gate1829(.a(G1291), .O(gate514inter8));
  nand2 gate1830(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate1831(.a(s_183), .b(gate514inter3), .O(gate514inter10));
  nor2  gate1832(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate1833(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate1834(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule