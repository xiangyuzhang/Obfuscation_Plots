module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate121inter0, gate121inter1, gate121inter2, gate121inter3, gate121inter4, gate121inter5, gate121inter6, gate121inter7, gate121inter8, gate121inter9, gate121inter10, gate121inter11, gate121inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate269inter0, gate269inter1, gate269inter2, gate269inter3, gate269inter4, gate269inter5, gate269inter6, gate269inter7, gate269inter8, gate269inter9, gate269inter10, gate269inter11, gate269inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate855(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate856(.a(gate12inter0), .b(s_44), .O(gate12inter1));
  and2  gate857(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate858(.a(s_44), .O(gate12inter3));
  inv1  gate859(.a(s_45), .O(gate12inter4));
  nand2 gate860(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate861(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate862(.a(G7), .O(gate12inter7));
  inv1  gate863(.a(G8), .O(gate12inter8));
  nand2 gate864(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate865(.a(s_45), .b(gate12inter3), .O(gate12inter10));
  nor2  gate866(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate867(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate868(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate1387(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate1388(.a(gate23inter0), .b(s_120), .O(gate23inter1));
  and2  gate1389(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate1390(.a(s_120), .O(gate23inter3));
  inv1  gate1391(.a(s_121), .O(gate23inter4));
  nand2 gate1392(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate1393(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate1394(.a(G29), .O(gate23inter7));
  inv1  gate1395(.a(G30), .O(gate23inter8));
  nand2 gate1396(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate1397(.a(s_121), .b(gate23inter3), .O(gate23inter10));
  nor2  gate1398(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate1399(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate1400(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate1261(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate1262(.a(gate31inter0), .b(s_102), .O(gate31inter1));
  and2  gate1263(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate1264(.a(s_102), .O(gate31inter3));
  inv1  gate1265(.a(s_103), .O(gate31inter4));
  nand2 gate1266(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate1267(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate1268(.a(G4), .O(gate31inter7));
  inv1  gate1269(.a(G8), .O(gate31inter8));
  nand2 gate1270(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate1271(.a(s_103), .b(gate31inter3), .O(gate31inter10));
  nor2  gate1272(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate1273(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate1274(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate617(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate618(.a(gate65inter0), .b(s_10), .O(gate65inter1));
  and2  gate619(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate620(.a(s_10), .O(gate65inter3));
  inv1  gate621(.a(s_11), .O(gate65inter4));
  nand2 gate622(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate623(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate624(.a(G25), .O(gate65inter7));
  inv1  gate625(.a(G302), .O(gate65inter8));
  nand2 gate626(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate627(.a(s_11), .b(gate65inter3), .O(gate65inter10));
  nor2  gate628(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate629(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate630(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate1275(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate1276(.a(gate69inter0), .b(s_104), .O(gate69inter1));
  and2  gate1277(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate1278(.a(s_104), .O(gate69inter3));
  inv1  gate1279(.a(s_105), .O(gate69inter4));
  nand2 gate1280(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate1281(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate1282(.a(G29), .O(gate69inter7));
  inv1  gate1283(.a(G308), .O(gate69inter8));
  nand2 gate1284(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate1285(.a(s_105), .b(gate69inter3), .O(gate69inter10));
  nor2  gate1286(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate1287(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate1288(.a(gate69inter12), .b(gate69inter1), .O(G390));
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate1191(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate1192(.a(gate80inter0), .b(s_92), .O(gate80inter1));
  and2  gate1193(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate1194(.a(s_92), .O(gate80inter3));
  inv1  gate1195(.a(s_93), .O(gate80inter4));
  nand2 gate1196(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate1197(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate1198(.a(G14), .O(gate80inter7));
  inv1  gate1199(.a(G323), .O(gate80inter8));
  nand2 gate1200(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate1201(.a(s_93), .b(gate80inter3), .O(gate80inter10));
  nor2  gate1202(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate1203(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate1204(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );

  xor2  gate757(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate758(.a(gate87inter0), .b(s_30), .O(gate87inter1));
  and2  gate759(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate760(.a(s_30), .O(gate87inter3));
  inv1  gate761(.a(s_31), .O(gate87inter4));
  nand2 gate762(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate763(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate764(.a(G12), .O(gate87inter7));
  inv1  gate765(.a(G335), .O(gate87inter8));
  nand2 gate766(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate767(.a(s_31), .b(gate87inter3), .O(gate87inter10));
  nor2  gate768(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate769(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate770(.a(gate87inter12), .b(gate87inter1), .O(G408));

  xor2  gate1331(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate1332(.a(gate88inter0), .b(s_112), .O(gate88inter1));
  and2  gate1333(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate1334(.a(s_112), .O(gate88inter3));
  inv1  gate1335(.a(s_113), .O(gate88inter4));
  nand2 gate1336(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate1337(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate1338(.a(G16), .O(gate88inter7));
  inv1  gate1339(.a(G335), .O(gate88inter8));
  nand2 gate1340(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate1341(.a(s_113), .b(gate88inter3), .O(gate88inter10));
  nor2  gate1342(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate1343(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate1344(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate701(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate702(.a(gate91inter0), .b(s_22), .O(gate91inter1));
  and2  gate703(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate704(.a(s_22), .O(gate91inter3));
  inv1  gate705(.a(s_23), .O(gate91inter4));
  nand2 gate706(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate707(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate708(.a(G25), .O(gate91inter7));
  inv1  gate709(.a(G341), .O(gate91inter8));
  nand2 gate710(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate711(.a(s_23), .b(gate91inter3), .O(gate91inter10));
  nor2  gate712(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate713(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate714(.a(gate91inter12), .b(gate91inter1), .O(G412));
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate1037(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate1038(.a(gate98inter0), .b(s_70), .O(gate98inter1));
  and2  gate1039(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate1040(.a(s_70), .O(gate98inter3));
  inv1  gate1041(.a(s_71), .O(gate98inter4));
  nand2 gate1042(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1043(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1044(.a(G23), .O(gate98inter7));
  inv1  gate1045(.a(G350), .O(gate98inter8));
  nand2 gate1046(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1047(.a(s_71), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1048(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1049(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1050(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );

  xor2  gate981(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate982(.a(gate103inter0), .b(s_62), .O(gate103inter1));
  and2  gate983(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate984(.a(s_62), .O(gate103inter3));
  inv1  gate985(.a(s_63), .O(gate103inter4));
  nand2 gate986(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate987(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate988(.a(G28), .O(gate103inter7));
  inv1  gate989(.a(G359), .O(gate103inter8));
  nand2 gate990(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate991(.a(s_63), .b(gate103inter3), .O(gate103inter10));
  nor2  gate992(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate993(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate994(.a(gate103inter12), .b(gate103inter1), .O(G424));
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate1317(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate1318(.a(gate106inter0), .b(s_110), .O(gate106inter1));
  and2  gate1319(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate1320(.a(s_110), .O(gate106inter3));
  inv1  gate1321(.a(s_111), .O(gate106inter4));
  nand2 gate1322(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate1323(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate1324(.a(G364), .O(gate106inter7));
  inv1  gate1325(.a(G365), .O(gate106inter8));
  nand2 gate1326(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate1327(.a(s_111), .b(gate106inter3), .O(gate106inter10));
  nor2  gate1328(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate1329(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate1330(.a(gate106inter12), .b(gate106inter1), .O(G429));

  xor2  gate1079(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate1080(.a(gate107inter0), .b(s_76), .O(gate107inter1));
  and2  gate1081(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate1082(.a(s_76), .O(gate107inter3));
  inv1  gate1083(.a(s_77), .O(gate107inter4));
  nand2 gate1084(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate1085(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate1086(.a(G366), .O(gate107inter7));
  inv1  gate1087(.a(G367), .O(gate107inter8));
  nand2 gate1088(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate1089(.a(s_77), .b(gate107inter3), .O(gate107inter10));
  nor2  gate1090(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate1091(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate1092(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate1107(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate1108(.a(gate110inter0), .b(s_80), .O(gate110inter1));
  and2  gate1109(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate1110(.a(s_80), .O(gate110inter3));
  inv1  gate1111(.a(s_81), .O(gate110inter4));
  nand2 gate1112(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1113(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1114(.a(G372), .O(gate110inter7));
  inv1  gate1115(.a(G373), .O(gate110inter8));
  nand2 gate1116(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1117(.a(s_81), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1118(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1119(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1120(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate715(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate716(.a(gate115inter0), .b(s_24), .O(gate115inter1));
  and2  gate717(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate718(.a(s_24), .O(gate115inter3));
  inv1  gate719(.a(s_25), .O(gate115inter4));
  nand2 gate720(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate721(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate722(.a(G382), .O(gate115inter7));
  inv1  gate723(.a(G383), .O(gate115inter8));
  nand2 gate724(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate725(.a(s_25), .b(gate115inter3), .O(gate115inter10));
  nor2  gate726(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate727(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate728(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );

  xor2  gate561(.a(G395), .b(G394), .O(gate121inter0));
  nand2 gate562(.a(gate121inter0), .b(s_2), .O(gate121inter1));
  and2  gate563(.a(G395), .b(G394), .O(gate121inter2));
  inv1  gate564(.a(s_2), .O(gate121inter3));
  inv1  gate565(.a(s_3), .O(gate121inter4));
  nand2 gate566(.a(gate121inter4), .b(gate121inter3), .O(gate121inter5));
  nor2  gate567(.a(gate121inter5), .b(gate121inter2), .O(gate121inter6));
  inv1  gate568(.a(G394), .O(gate121inter7));
  inv1  gate569(.a(G395), .O(gate121inter8));
  nand2 gate570(.a(gate121inter8), .b(gate121inter7), .O(gate121inter9));
  nand2 gate571(.a(s_3), .b(gate121inter3), .O(gate121inter10));
  nor2  gate572(.a(gate121inter10), .b(gate121inter9), .O(gate121inter11));
  nor2  gate573(.a(gate121inter11), .b(gate121inter6), .O(gate121inter12));
  nand2 gate574(.a(gate121inter12), .b(gate121inter1), .O(G474));
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate1233(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate1234(.a(gate124inter0), .b(s_98), .O(gate124inter1));
  and2  gate1235(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate1236(.a(s_98), .O(gate124inter3));
  inv1  gate1237(.a(s_99), .O(gate124inter4));
  nand2 gate1238(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate1239(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate1240(.a(G400), .O(gate124inter7));
  inv1  gate1241(.a(G401), .O(gate124inter8));
  nand2 gate1242(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate1243(.a(s_99), .b(gate124inter3), .O(gate124inter10));
  nor2  gate1244(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate1245(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate1246(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate827(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate828(.a(gate128inter0), .b(s_40), .O(gate128inter1));
  and2  gate829(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate830(.a(s_40), .O(gate128inter3));
  inv1  gate831(.a(s_41), .O(gate128inter4));
  nand2 gate832(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate833(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate834(.a(G408), .O(gate128inter7));
  inv1  gate835(.a(G409), .O(gate128inter8));
  nand2 gate836(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate837(.a(s_41), .b(gate128inter3), .O(gate128inter10));
  nor2  gate838(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate839(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate840(.a(gate128inter12), .b(gate128inter1), .O(G495));
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );

  xor2  gate1149(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate1150(.a(gate133inter0), .b(s_86), .O(gate133inter1));
  and2  gate1151(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate1152(.a(s_86), .O(gate133inter3));
  inv1  gate1153(.a(s_87), .O(gate133inter4));
  nand2 gate1154(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate1155(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate1156(.a(G418), .O(gate133inter7));
  inv1  gate1157(.a(G419), .O(gate133inter8));
  nand2 gate1158(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate1159(.a(s_87), .b(gate133inter3), .O(gate133inter10));
  nor2  gate1160(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate1161(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate1162(.a(gate133inter12), .b(gate133inter1), .O(G510));
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate1205(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate1206(.a(gate144inter0), .b(s_94), .O(gate144inter1));
  and2  gate1207(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate1208(.a(s_94), .O(gate144inter3));
  inv1  gate1209(.a(s_95), .O(gate144inter4));
  nand2 gate1210(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate1211(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate1212(.a(G468), .O(gate144inter7));
  inv1  gate1213(.a(G471), .O(gate144inter8));
  nand2 gate1214(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate1215(.a(s_95), .b(gate144inter3), .O(gate144inter10));
  nor2  gate1216(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate1217(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate1218(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );

  xor2  gate687(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate688(.a(gate146inter0), .b(s_20), .O(gate146inter1));
  and2  gate689(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate690(.a(s_20), .O(gate146inter3));
  inv1  gate691(.a(s_21), .O(gate146inter4));
  nand2 gate692(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate693(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate694(.a(G480), .O(gate146inter7));
  inv1  gate695(.a(G483), .O(gate146inter8));
  nand2 gate696(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate697(.a(s_21), .b(gate146inter3), .O(gate146inter10));
  nor2  gate698(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate699(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate700(.a(gate146inter12), .b(gate146inter1), .O(G549));
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate673(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate674(.a(gate153inter0), .b(s_18), .O(gate153inter1));
  and2  gate675(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate676(.a(s_18), .O(gate153inter3));
  inv1  gate677(.a(s_19), .O(gate153inter4));
  nand2 gate678(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate679(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate680(.a(G426), .O(gate153inter7));
  inv1  gate681(.a(G522), .O(gate153inter8));
  nand2 gate682(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate683(.a(s_19), .b(gate153inter3), .O(gate153inter10));
  nor2  gate684(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate685(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate686(.a(gate153inter12), .b(gate153inter1), .O(G570));
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate995(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate996(.a(gate159inter0), .b(s_64), .O(gate159inter1));
  and2  gate997(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate998(.a(s_64), .O(gate159inter3));
  inv1  gate999(.a(s_65), .O(gate159inter4));
  nand2 gate1000(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate1001(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate1002(.a(G444), .O(gate159inter7));
  inv1  gate1003(.a(G531), .O(gate159inter8));
  nand2 gate1004(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate1005(.a(s_65), .b(gate159inter3), .O(gate159inter10));
  nor2  gate1006(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate1007(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate1008(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );

  xor2  gate1163(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate1164(.a(gate163inter0), .b(s_88), .O(gate163inter1));
  and2  gate1165(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate1166(.a(s_88), .O(gate163inter3));
  inv1  gate1167(.a(s_89), .O(gate163inter4));
  nand2 gate1168(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate1169(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate1170(.a(G456), .O(gate163inter7));
  inv1  gate1171(.a(G537), .O(gate163inter8));
  nand2 gate1172(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate1173(.a(s_89), .b(gate163inter3), .O(gate163inter10));
  nor2  gate1174(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate1175(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate1176(.a(gate163inter12), .b(gate163inter1), .O(G580));
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );

  xor2  gate645(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate646(.a(gate166inter0), .b(s_14), .O(gate166inter1));
  and2  gate647(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate648(.a(s_14), .O(gate166inter3));
  inv1  gate649(.a(s_15), .O(gate166inter4));
  nand2 gate650(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate651(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate652(.a(G465), .O(gate166inter7));
  inv1  gate653(.a(G540), .O(gate166inter8));
  nand2 gate654(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate655(.a(s_15), .b(gate166inter3), .O(gate166inter10));
  nor2  gate656(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate657(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate658(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate785(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate786(.a(gate173inter0), .b(s_34), .O(gate173inter1));
  and2  gate787(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate788(.a(s_34), .O(gate173inter3));
  inv1  gate789(.a(s_35), .O(gate173inter4));
  nand2 gate790(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate791(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate792(.a(G486), .O(gate173inter7));
  inv1  gate793(.a(G552), .O(gate173inter8));
  nand2 gate794(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate795(.a(s_35), .b(gate173inter3), .O(gate173inter10));
  nor2  gate796(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate797(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate798(.a(gate173inter12), .b(gate173inter1), .O(G590));

  xor2  gate925(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate926(.a(gate174inter0), .b(s_54), .O(gate174inter1));
  and2  gate927(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate928(.a(s_54), .O(gate174inter3));
  inv1  gate929(.a(s_55), .O(gate174inter4));
  nand2 gate930(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate931(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate932(.a(G489), .O(gate174inter7));
  inv1  gate933(.a(G552), .O(gate174inter8));
  nand2 gate934(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate935(.a(s_55), .b(gate174inter3), .O(gate174inter10));
  nor2  gate936(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate937(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate938(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate813(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate814(.a(gate180inter0), .b(s_38), .O(gate180inter1));
  and2  gate815(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate816(.a(s_38), .O(gate180inter3));
  inv1  gate817(.a(s_39), .O(gate180inter4));
  nand2 gate818(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate819(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate820(.a(G507), .O(gate180inter7));
  inv1  gate821(.a(G561), .O(gate180inter8));
  nand2 gate822(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate823(.a(s_39), .b(gate180inter3), .O(gate180inter10));
  nor2  gate824(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate825(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate826(.a(gate180inter12), .b(gate180inter1), .O(G597));
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate799(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate800(.a(gate187inter0), .b(s_36), .O(gate187inter1));
  and2  gate801(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate802(.a(s_36), .O(gate187inter3));
  inv1  gate803(.a(s_37), .O(gate187inter4));
  nand2 gate804(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate805(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate806(.a(G574), .O(gate187inter7));
  inv1  gate807(.a(G575), .O(gate187inter8));
  nand2 gate808(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate809(.a(s_37), .b(gate187inter3), .O(gate187inter10));
  nor2  gate810(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate811(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate812(.a(gate187inter12), .b(gate187inter1), .O(G612));
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate547(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate548(.a(gate193inter0), .b(s_0), .O(gate193inter1));
  and2  gate549(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate550(.a(s_0), .O(gate193inter3));
  inv1  gate551(.a(s_1), .O(gate193inter4));
  nand2 gate552(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate553(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate554(.a(G586), .O(gate193inter7));
  inv1  gate555(.a(G587), .O(gate193inter8));
  nand2 gate556(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate557(.a(s_1), .b(gate193inter3), .O(gate193inter10));
  nor2  gate558(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate559(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate560(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate841(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate842(.a(gate213inter0), .b(s_42), .O(gate213inter1));
  and2  gate843(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate844(.a(s_42), .O(gate213inter3));
  inv1  gate845(.a(s_43), .O(gate213inter4));
  nand2 gate846(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate847(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate848(.a(G602), .O(gate213inter7));
  inv1  gate849(.a(G672), .O(gate213inter8));
  nand2 gate850(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate851(.a(s_43), .b(gate213inter3), .O(gate213inter10));
  nor2  gate852(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate853(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate854(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate953(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate954(.a(gate219inter0), .b(s_58), .O(gate219inter1));
  and2  gate955(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate956(.a(s_58), .O(gate219inter3));
  inv1  gate957(.a(s_59), .O(gate219inter4));
  nand2 gate958(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate959(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate960(.a(G632), .O(gate219inter7));
  inv1  gate961(.a(G681), .O(gate219inter8));
  nand2 gate962(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate963(.a(s_59), .b(gate219inter3), .O(gate219inter10));
  nor2  gate964(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate965(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate966(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate1065(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate1066(.a(gate237inter0), .b(s_74), .O(gate237inter1));
  and2  gate1067(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate1068(.a(s_74), .O(gate237inter3));
  inv1  gate1069(.a(s_75), .O(gate237inter4));
  nand2 gate1070(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1071(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1072(.a(G254), .O(gate237inter7));
  inv1  gate1073(.a(G706), .O(gate237inter8));
  nand2 gate1074(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1075(.a(s_75), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1076(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1077(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1078(.a(gate237inter12), .b(gate237inter1), .O(G742));

  xor2  gate1051(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate1052(.a(gate238inter0), .b(s_72), .O(gate238inter1));
  and2  gate1053(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate1054(.a(s_72), .O(gate238inter3));
  inv1  gate1055(.a(s_73), .O(gate238inter4));
  nand2 gate1056(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate1057(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate1058(.a(G257), .O(gate238inter7));
  inv1  gate1059(.a(G709), .O(gate238inter8));
  nand2 gate1060(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate1061(.a(s_73), .b(gate238inter3), .O(gate238inter10));
  nor2  gate1062(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate1063(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate1064(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate1135(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate1136(.a(gate241inter0), .b(s_84), .O(gate241inter1));
  and2  gate1137(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate1138(.a(s_84), .O(gate241inter3));
  inv1  gate1139(.a(s_85), .O(gate241inter4));
  nand2 gate1140(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate1141(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate1142(.a(G242), .O(gate241inter7));
  inv1  gate1143(.a(G730), .O(gate241inter8));
  nand2 gate1144(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate1145(.a(s_85), .b(gate241inter3), .O(gate241inter10));
  nor2  gate1146(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate1147(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate1148(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate883(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate884(.a(gate243inter0), .b(s_48), .O(gate243inter1));
  and2  gate885(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate886(.a(s_48), .O(gate243inter3));
  inv1  gate887(.a(s_49), .O(gate243inter4));
  nand2 gate888(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate889(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate890(.a(G245), .O(gate243inter7));
  inv1  gate891(.a(G733), .O(gate243inter8));
  nand2 gate892(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate893(.a(s_49), .b(gate243inter3), .O(gate243inter10));
  nor2  gate894(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate895(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate896(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );

  xor2  gate897(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate898(.a(gate254inter0), .b(s_50), .O(gate254inter1));
  and2  gate899(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate900(.a(s_50), .O(gate254inter3));
  inv1  gate901(.a(s_51), .O(gate254inter4));
  nand2 gate902(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate903(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate904(.a(G712), .O(gate254inter7));
  inv1  gate905(.a(G748), .O(gate254inter8));
  nand2 gate906(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate907(.a(s_51), .b(gate254inter3), .O(gate254inter10));
  nor2  gate908(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate909(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate910(.a(gate254inter12), .b(gate254inter1), .O(G767));
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate1177(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate1178(.a(gate257inter0), .b(s_90), .O(gate257inter1));
  and2  gate1179(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate1180(.a(s_90), .O(gate257inter3));
  inv1  gate1181(.a(s_91), .O(gate257inter4));
  nand2 gate1182(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate1183(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate1184(.a(G754), .O(gate257inter7));
  inv1  gate1185(.a(G755), .O(gate257inter8));
  nand2 gate1186(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate1187(.a(s_91), .b(gate257inter3), .O(gate257inter10));
  nor2  gate1188(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate1189(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate1190(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );

  xor2  gate743(.a(G782), .b(G654), .O(gate269inter0));
  nand2 gate744(.a(gate269inter0), .b(s_28), .O(gate269inter1));
  and2  gate745(.a(G782), .b(G654), .O(gate269inter2));
  inv1  gate746(.a(s_28), .O(gate269inter3));
  inv1  gate747(.a(s_29), .O(gate269inter4));
  nand2 gate748(.a(gate269inter4), .b(gate269inter3), .O(gate269inter5));
  nor2  gate749(.a(gate269inter5), .b(gate269inter2), .O(gate269inter6));
  inv1  gate750(.a(G654), .O(gate269inter7));
  inv1  gate751(.a(G782), .O(gate269inter8));
  nand2 gate752(.a(gate269inter8), .b(gate269inter7), .O(gate269inter9));
  nand2 gate753(.a(s_29), .b(gate269inter3), .O(gate269inter10));
  nor2  gate754(.a(gate269inter10), .b(gate269inter9), .O(gate269inter11));
  nor2  gate755(.a(gate269inter11), .b(gate269inter6), .O(gate269inter12));
  nand2 gate756(.a(gate269inter12), .b(gate269inter1), .O(G806));
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate575(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate576(.a(gate280inter0), .b(s_4), .O(gate280inter1));
  and2  gate577(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate578(.a(s_4), .O(gate280inter3));
  inv1  gate579(.a(s_5), .O(gate280inter4));
  nand2 gate580(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate581(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate582(.a(G779), .O(gate280inter7));
  inv1  gate583(.a(G803), .O(gate280inter8));
  nand2 gate584(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate585(.a(s_5), .b(gate280inter3), .O(gate280inter10));
  nor2  gate586(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate587(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate588(.a(gate280inter12), .b(gate280inter1), .O(G825));

  xor2  gate1023(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate1024(.a(gate281inter0), .b(s_68), .O(gate281inter1));
  and2  gate1025(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate1026(.a(s_68), .O(gate281inter3));
  inv1  gate1027(.a(s_69), .O(gate281inter4));
  nand2 gate1028(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate1029(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate1030(.a(G654), .O(gate281inter7));
  inv1  gate1031(.a(G806), .O(gate281inter8));
  nand2 gate1032(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate1033(.a(s_69), .b(gate281inter3), .O(gate281inter10));
  nor2  gate1034(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate1035(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate1036(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate729(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate730(.a(gate296inter0), .b(s_26), .O(gate296inter1));
  and2  gate731(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate732(.a(s_26), .O(gate296inter3));
  inv1  gate733(.a(s_27), .O(gate296inter4));
  nand2 gate734(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate735(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate736(.a(G826), .O(gate296inter7));
  inv1  gate737(.a(G827), .O(gate296inter8));
  nand2 gate738(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate739(.a(s_27), .b(gate296inter3), .O(gate296inter10));
  nor2  gate740(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate741(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate742(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate1289(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate1290(.a(gate387inter0), .b(s_106), .O(gate387inter1));
  and2  gate1291(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate1292(.a(s_106), .O(gate387inter3));
  inv1  gate1293(.a(s_107), .O(gate387inter4));
  nand2 gate1294(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1295(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1296(.a(G1), .O(gate387inter7));
  inv1  gate1297(.a(G1036), .O(gate387inter8));
  nand2 gate1298(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1299(.a(s_107), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1300(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1301(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate1302(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );

  xor2  gate939(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate940(.a(gate408inter0), .b(s_56), .O(gate408inter1));
  and2  gate941(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate942(.a(s_56), .O(gate408inter3));
  inv1  gate943(.a(s_57), .O(gate408inter4));
  nand2 gate944(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate945(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate946(.a(G22), .O(gate408inter7));
  inv1  gate947(.a(G1099), .O(gate408inter8));
  nand2 gate948(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate949(.a(s_57), .b(gate408inter3), .O(gate408inter10));
  nor2  gate950(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate951(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate952(.a(gate408inter12), .b(gate408inter1), .O(G1195));

  xor2  gate1093(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate1094(.a(gate409inter0), .b(s_78), .O(gate409inter1));
  and2  gate1095(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate1096(.a(s_78), .O(gate409inter3));
  inv1  gate1097(.a(s_79), .O(gate409inter4));
  nand2 gate1098(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate1099(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate1100(.a(G23), .O(gate409inter7));
  inv1  gate1101(.a(G1102), .O(gate409inter8));
  nand2 gate1102(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate1103(.a(s_79), .b(gate409inter3), .O(gate409inter10));
  nor2  gate1104(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate1105(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate1106(.a(gate409inter12), .b(gate409inter1), .O(G1198));
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate1219(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate1220(.a(gate411inter0), .b(s_96), .O(gate411inter1));
  and2  gate1221(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate1222(.a(s_96), .O(gate411inter3));
  inv1  gate1223(.a(s_97), .O(gate411inter4));
  nand2 gate1224(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate1225(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate1226(.a(G25), .O(gate411inter7));
  inv1  gate1227(.a(G1108), .O(gate411inter8));
  nand2 gate1228(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate1229(.a(s_97), .b(gate411inter3), .O(gate411inter10));
  nor2  gate1230(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate1231(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate1232(.a(gate411inter12), .b(gate411inter1), .O(G1204));

  xor2  gate631(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate632(.a(gate412inter0), .b(s_12), .O(gate412inter1));
  and2  gate633(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate634(.a(s_12), .O(gate412inter3));
  inv1  gate635(.a(s_13), .O(gate412inter4));
  nand2 gate636(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate637(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate638(.a(G26), .O(gate412inter7));
  inv1  gate639(.a(G1111), .O(gate412inter8));
  nand2 gate640(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate641(.a(s_13), .b(gate412inter3), .O(gate412inter10));
  nor2  gate642(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate643(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate644(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate1121(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate1122(.a(gate419inter0), .b(s_82), .O(gate419inter1));
  and2  gate1123(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate1124(.a(s_82), .O(gate419inter3));
  inv1  gate1125(.a(s_83), .O(gate419inter4));
  nand2 gate1126(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate1127(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate1128(.a(G1), .O(gate419inter7));
  inv1  gate1129(.a(G1132), .O(gate419inter8));
  nand2 gate1130(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate1131(.a(s_83), .b(gate419inter3), .O(gate419inter10));
  nor2  gate1132(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate1133(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate1134(.a(gate419inter12), .b(gate419inter1), .O(G1228));
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate771(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate772(.a(gate428inter0), .b(s_32), .O(gate428inter1));
  and2  gate773(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate774(.a(s_32), .O(gate428inter3));
  inv1  gate775(.a(s_33), .O(gate428inter4));
  nand2 gate776(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate777(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate778(.a(G1048), .O(gate428inter7));
  inv1  gate779(.a(G1144), .O(gate428inter8));
  nand2 gate780(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate781(.a(s_33), .b(gate428inter3), .O(gate428inter10));
  nor2  gate782(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate783(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate784(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate659(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate660(.a(gate443inter0), .b(s_16), .O(gate443inter1));
  and2  gate661(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate662(.a(s_16), .O(gate443inter3));
  inv1  gate663(.a(s_17), .O(gate443inter4));
  nand2 gate664(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate665(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate666(.a(G13), .O(gate443inter7));
  inv1  gate667(.a(G1168), .O(gate443inter8));
  nand2 gate668(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate669(.a(s_17), .b(gate443inter3), .O(gate443inter10));
  nor2  gate670(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate671(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate672(.a(gate443inter12), .b(gate443inter1), .O(G1252));

  xor2  gate1247(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate1248(.a(gate444inter0), .b(s_100), .O(gate444inter1));
  and2  gate1249(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate1250(.a(s_100), .O(gate444inter3));
  inv1  gate1251(.a(s_101), .O(gate444inter4));
  nand2 gate1252(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate1253(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate1254(.a(G1072), .O(gate444inter7));
  inv1  gate1255(.a(G1168), .O(gate444inter8));
  nand2 gate1256(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate1257(.a(s_101), .b(gate444inter3), .O(gate444inter10));
  nor2  gate1258(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate1259(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate1260(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate1303(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate1304(.a(gate464inter0), .b(s_108), .O(gate464inter1));
  and2  gate1305(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate1306(.a(s_108), .O(gate464inter3));
  inv1  gate1307(.a(s_109), .O(gate464inter4));
  nand2 gate1308(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate1309(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate1310(.a(G1102), .O(gate464inter7));
  inv1  gate1311(.a(G1198), .O(gate464inter8));
  nand2 gate1312(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate1313(.a(s_109), .b(gate464inter3), .O(gate464inter10));
  nor2  gate1314(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate1315(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate1316(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );

  xor2  gate967(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate968(.a(gate468inter0), .b(s_60), .O(gate468inter1));
  and2  gate969(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate970(.a(s_60), .O(gate468inter3));
  inv1  gate971(.a(s_61), .O(gate468inter4));
  nand2 gate972(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate973(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate974(.a(G1108), .O(gate468inter7));
  inv1  gate975(.a(G1204), .O(gate468inter8));
  nand2 gate976(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate977(.a(s_61), .b(gate468inter3), .O(gate468inter10));
  nor2  gate978(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate979(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate980(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate1345(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate1346(.a(gate474inter0), .b(s_114), .O(gate474inter1));
  and2  gate1347(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate1348(.a(s_114), .O(gate474inter3));
  inv1  gate1349(.a(s_115), .O(gate474inter4));
  nand2 gate1350(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate1351(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate1352(.a(G1117), .O(gate474inter7));
  inv1  gate1353(.a(G1213), .O(gate474inter8));
  nand2 gate1354(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate1355(.a(s_115), .b(gate474inter3), .O(gate474inter10));
  nor2  gate1356(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate1357(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate1358(.a(gate474inter12), .b(gate474inter1), .O(G1283));
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate869(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate870(.a(gate476inter0), .b(s_46), .O(gate476inter1));
  and2  gate871(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate872(.a(s_46), .O(gate476inter3));
  inv1  gate873(.a(s_47), .O(gate476inter4));
  nand2 gate874(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate875(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate876(.a(G1120), .O(gate476inter7));
  inv1  gate877(.a(G1216), .O(gate476inter8));
  nand2 gate878(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate879(.a(s_47), .b(gate476inter3), .O(gate476inter10));
  nor2  gate880(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate881(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate882(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate1359(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate1360(.a(gate485inter0), .b(s_116), .O(gate485inter1));
  and2  gate1361(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate1362(.a(s_116), .O(gate485inter3));
  inv1  gate1363(.a(s_117), .O(gate485inter4));
  nand2 gate1364(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate1365(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate1366(.a(G1232), .O(gate485inter7));
  inv1  gate1367(.a(G1233), .O(gate485inter8));
  nand2 gate1368(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate1369(.a(s_117), .b(gate485inter3), .O(gate485inter10));
  nor2  gate1370(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate1371(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate1372(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate911(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate912(.a(gate493inter0), .b(s_52), .O(gate493inter1));
  and2  gate913(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate914(.a(s_52), .O(gate493inter3));
  inv1  gate915(.a(s_53), .O(gate493inter4));
  nand2 gate916(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate917(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate918(.a(G1248), .O(gate493inter7));
  inv1  gate919(.a(G1249), .O(gate493inter8));
  nand2 gate920(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate921(.a(s_53), .b(gate493inter3), .O(gate493inter10));
  nor2  gate922(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate923(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate924(.a(gate493inter12), .b(gate493inter1), .O(G1302));
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate603(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate604(.a(gate503inter0), .b(s_8), .O(gate503inter1));
  and2  gate605(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate606(.a(s_8), .O(gate503inter3));
  inv1  gate607(.a(s_9), .O(gate503inter4));
  nand2 gate608(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate609(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate610(.a(G1268), .O(gate503inter7));
  inv1  gate611(.a(G1269), .O(gate503inter8));
  nand2 gate612(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate613(.a(s_9), .b(gate503inter3), .O(gate503inter10));
  nor2  gate614(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate615(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate616(.a(gate503inter12), .b(gate503inter1), .O(G1312));
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );

  xor2  gate1009(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate1010(.a(gate505inter0), .b(s_66), .O(gate505inter1));
  and2  gate1011(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate1012(.a(s_66), .O(gate505inter3));
  inv1  gate1013(.a(s_67), .O(gate505inter4));
  nand2 gate1014(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate1015(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate1016(.a(G1272), .O(gate505inter7));
  inv1  gate1017(.a(G1273), .O(gate505inter8));
  nand2 gate1018(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate1019(.a(s_67), .b(gate505inter3), .O(gate505inter10));
  nor2  gate1020(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate1021(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate1022(.a(gate505inter12), .b(gate505inter1), .O(G1314));

  xor2  gate1373(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate1374(.a(gate506inter0), .b(s_118), .O(gate506inter1));
  and2  gate1375(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate1376(.a(s_118), .O(gate506inter3));
  inv1  gate1377(.a(s_119), .O(gate506inter4));
  nand2 gate1378(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate1379(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate1380(.a(G1274), .O(gate506inter7));
  inv1  gate1381(.a(G1275), .O(gate506inter8));
  nand2 gate1382(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate1383(.a(s_119), .b(gate506inter3), .O(gate506inter10));
  nor2  gate1384(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate1385(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate1386(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate589(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate590(.a(gate514inter0), .b(s_6), .O(gate514inter1));
  and2  gate591(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate592(.a(s_6), .O(gate514inter3));
  inv1  gate593(.a(s_7), .O(gate514inter4));
  nand2 gate594(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate595(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate596(.a(G1290), .O(gate514inter7));
  inv1  gate597(.a(G1291), .O(gate514inter8));
  nand2 gate598(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate599(.a(s_7), .b(gate514inter3), .O(gate514inter10));
  nor2  gate600(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate601(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate602(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule