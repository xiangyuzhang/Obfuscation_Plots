module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281, s_282, s_283, s_284, s_285, s_286, s_287, s_288, s_289, s_290, s_291, s_292, s_293, s_294, s_295, s_296, s_297, s_298, s_299, s_300, s_301;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate18inter0, gate18inter1, gate18inter2, gate18inter3, gate18inter4, gate18inter5, gate18inter6, gate18inter7, gate18inter8, gate18inter9, gate18inter10, gate18inter11, gate18inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate499inter0, gate499inter1, gate499inter2, gate499inter3, gate499inter4, gate499inter5, gate499inter6, gate499inter7, gate499inter8, gate499inter9, gate499inter10, gate499inter11, gate499inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate101inter0, gate101inter1, gate101inter2, gate101inter3, gate101inter4, gate101inter5, gate101inter6, gate101inter7, gate101inter8, gate101inter9, gate101inter10, gate101inter11, gate101inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate266inter0, gate266inter1, gate266inter2, gate266inter3, gate266inter4, gate266inter5, gate266inter6, gate266inter7, gate266inter8, gate266inter9, gate266inter10, gate266inter11, gate266inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate513inter0, gate513inter1, gate513inter2, gate513inter3, gate513inter4, gate513inter5, gate513inter6, gate513inter7, gate513inter8, gate513inter9, gate513inter10, gate513inter11, gate513inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate2157(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate2158(.a(gate12inter0), .b(s_230), .O(gate12inter1));
  and2  gate2159(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate2160(.a(s_230), .O(gate12inter3));
  inv1  gate2161(.a(s_231), .O(gate12inter4));
  nand2 gate2162(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate2163(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate2164(.a(G7), .O(gate12inter7));
  inv1  gate2165(.a(G8), .O(gate12inter8));
  nand2 gate2166(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate2167(.a(s_231), .b(gate12inter3), .O(gate12inter10));
  nor2  gate2168(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate2169(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate2170(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );

  xor2  gate1079(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate1080(.a(gate14inter0), .b(s_76), .O(gate14inter1));
  and2  gate1081(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate1082(.a(s_76), .O(gate14inter3));
  inv1  gate1083(.a(s_77), .O(gate14inter4));
  nand2 gate1084(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate1085(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate1086(.a(G11), .O(gate14inter7));
  inv1  gate1087(.a(G12), .O(gate14inter8));
  nand2 gate1088(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate1089(.a(s_77), .b(gate14inter3), .O(gate14inter10));
  nor2  gate1090(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate1091(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate1092(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate1765(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate1766(.a(gate16inter0), .b(s_174), .O(gate16inter1));
  and2  gate1767(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate1768(.a(s_174), .O(gate16inter3));
  inv1  gate1769(.a(s_175), .O(gate16inter4));
  nand2 gate1770(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate1771(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate1772(.a(G15), .O(gate16inter7));
  inv1  gate1773(.a(G16), .O(gate16inter8));
  nand2 gate1774(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate1775(.a(s_175), .b(gate16inter3), .O(gate16inter10));
  nor2  gate1776(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate1777(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate1778(.a(gate16inter12), .b(gate16inter1), .O(G287));

  xor2  gate2297(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate2298(.a(gate17inter0), .b(s_250), .O(gate17inter1));
  and2  gate2299(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate2300(.a(s_250), .O(gate17inter3));
  inv1  gate2301(.a(s_251), .O(gate17inter4));
  nand2 gate2302(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate2303(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate2304(.a(G17), .O(gate17inter7));
  inv1  gate2305(.a(G18), .O(gate17inter8));
  nand2 gate2306(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate2307(.a(s_251), .b(gate17inter3), .O(gate17inter10));
  nor2  gate2308(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate2309(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate2310(.a(gate17inter12), .b(gate17inter1), .O(G290));

  xor2  gate645(.a(G20), .b(G19), .O(gate18inter0));
  nand2 gate646(.a(gate18inter0), .b(s_14), .O(gate18inter1));
  and2  gate647(.a(G20), .b(G19), .O(gate18inter2));
  inv1  gate648(.a(s_14), .O(gate18inter3));
  inv1  gate649(.a(s_15), .O(gate18inter4));
  nand2 gate650(.a(gate18inter4), .b(gate18inter3), .O(gate18inter5));
  nor2  gate651(.a(gate18inter5), .b(gate18inter2), .O(gate18inter6));
  inv1  gate652(.a(G19), .O(gate18inter7));
  inv1  gate653(.a(G20), .O(gate18inter8));
  nand2 gate654(.a(gate18inter8), .b(gate18inter7), .O(gate18inter9));
  nand2 gate655(.a(s_15), .b(gate18inter3), .O(gate18inter10));
  nor2  gate656(.a(gate18inter10), .b(gate18inter9), .O(gate18inter11));
  nor2  gate657(.a(gate18inter11), .b(gate18inter6), .O(gate18inter12));
  nand2 gate658(.a(gate18inter12), .b(gate18inter1), .O(G293));
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate1219(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate1220(.a(gate20inter0), .b(s_96), .O(gate20inter1));
  and2  gate1221(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate1222(.a(s_96), .O(gate20inter3));
  inv1  gate1223(.a(s_97), .O(gate20inter4));
  nand2 gate1224(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate1225(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate1226(.a(G23), .O(gate20inter7));
  inv1  gate1227(.a(G24), .O(gate20inter8));
  nand2 gate1228(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate1229(.a(s_97), .b(gate20inter3), .O(gate20inter10));
  nor2  gate1230(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate1231(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate1232(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate2283(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate2284(.a(gate25inter0), .b(s_248), .O(gate25inter1));
  and2  gate2285(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate2286(.a(s_248), .O(gate25inter3));
  inv1  gate2287(.a(s_249), .O(gate25inter4));
  nand2 gate2288(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate2289(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate2290(.a(G1), .O(gate25inter7));
  inv1  gate2291(.a(G5), .O(gate25inter8));
  nand2 gate2292(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate2293(.a(s_249), .b(gate25inter3), .O(gate25inter10));
  nor2  gate2294(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate2295(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate2296(.a(gate25inter12), .b(gate25inter1), .O(G314));

  xor2  gate1807(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate1808(.a(gate26inter0), .b(s_180), .O(gate26inter1));
  and2  gate1809(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate1810(.a(s_180), .O(gate26inter3));
  inv1  gate1811(.a(s_181), .O(gate26inter4));
  nand2 gate1812(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate1813(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate1814(.a(G9), .O(gate26inter7));
  inv1  gate1815(.a(G13), .O(gate26inter8));
  nand2 gate1816(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate1817(.a(s_181), .b(gate26inter3), .O(gate26inter10));
  nor2  gate1818(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate1819(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate1820(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );

  xor2  gate869(.a(G14), .b(G10), .O(gate28inter0));
  nand2 gate870(.a(gate28inter0), .b(s_46), .O(gate28inter1));
  and2  gate871(.a(G14), .b(G10), .O(gate28inter2));
  inv1  gate872(.a(s_46), .O(gate28inter3));
  inv1  gate873(.a(s_47), .O(gate28inter4));
  nand2 gate874(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate875(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate876(.a(G10), .O(gate28inter7));
  inv1  gate877(.a(G14), .O(gate28inter8));
  nand2 gate878(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate879(.a(s_47), .b(gate28inter3), .O(gate28inter10));
  nor2  gate880(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate881(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate882(.a(gate28inter12), .b(gate28inter1), .O(G323));

  xor2  gate2619(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate2620(.a(gate29inter0), .b(s_296), .O(gate29inter1));
  and2  gate2621(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate2622(.a(s_296), .O(gate29inter3));
  inv1  gate2623(.a(s_297), .O(gate29inter4));
  nand2 gate2624(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate2625(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate2626(.a(G3), .O(gate29inter7));
  inv1  gate2627(.a(G7), .O(gate29inter8));
  nand2 gate2628(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate2629(.a(s_297), .b(gate29inter3), .O(gate29inter10));
  nor2  gate2630(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate2631(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate2632(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );

  xor2  gate1737(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate1738(.a(gate32inter0), .b(s_170), .O(gate32inter1));
  and2  gate1739(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate1740(.a(s_170), .O(gate32inter3));
  inv1  gate1741(.a(s_171), .O(gate32inter4));
  nand2 gate1742(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate1743(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate1744(.a(G12), .O(gate32inter7));
  inv1  gate1745(.a(G16), .O(gate32inter8));
  nand2 gate1746(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate1747(.a(s_171), .b(gate32inter3), .O(gate32inter10));
  nor2  gate1748(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate1749(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate1750(.a(gate32inter12), .b(gate32inter1), .O(G335));
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate911(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate912(.a(gate34inter0), .b(s_52), .O(gate34inter1));
  and2  gate913(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate914(.a(s_52), .O(gate34inter3));
  inv1  gate915(.a(s_53), .O(gate34inter4));
  nand2 gate916(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate917(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate918(.a(G25), .O(gate34inter7));
  inv1  gate919(.a(G29), .O(gate34inter8));
  nand2 gate920(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate921(.a(s_53), .b(gate34inter3), .O(gate34inter10));
  nor2  gate922(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate923(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate924(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate1779(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate1780(.a(gate37inter0), .b(s_176), .O(gate37inter1));
  and2  gate1781(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate1782(.a(s_176), .O(gate37inter3));
  inv1  gate1783(.a(s_177), .O(gate37inter4));
  nand2 gate1784(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate1785(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate1786(.a(G19), .O(gate37inter7));
  inv1  gate1787(.a(G23), .O(gate37inter8));
  nand2 gate1788(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate1789(.a(s_177), .b(gate37inter3), .O(gate37inter10));
  nor2  gate1790(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate1791(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate1792(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );

  xor2  gate2563(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate2564(.a(gate42inter0), .b(s_288), .O(gate42inter1));
  and2  gate2565(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate2566(.a(s_288), .O(gate42inter3));
  inv1  gate2567(.a(s_289), .O(gate42inter4));
  nand2 gate2568(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate2569(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate2570(.a(G2), .O(gate42inter7));
  inv1  gate2571(.a(G266), .O(gate42inter8));
  nand2 gate2572(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate2573(.a(s_289), .b(gate42inter3), .O(gate42inter10));
  nor2  gate2574(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate2575(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate2576(.a(gate42inter12), .b(gate42inter1), .O(G363));
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );

  xor2  gate1625(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate1626(.a(gate45inter0), .b(s_154), .O(gate45inter1));
  and2  gate1627(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate1628(.a(s_154), .O(gate45inter3));
  inv1  gate1629(.a(s_155), .O(gate45inter4));
  nand2 gate1630(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate1631(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate1632(.a(G5), .O(gate45inter7));
  inv1  gate1633(.a(G272), .O(gate45inter8));
  nand2 gate1634(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate1635(.a(s_155), .b(gate45inter3), .O(gate45inter10));
  nor2  gate1636(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate1637(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate1638(.a(gate45inter12), .b(gate45inter1), .O(G366));

  xor2  gate1317(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate1318(.a(gate46inter0), .b(s_110), .O(gate46inter1));
  and2  gate1319(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate1320(.a(s_110), .O(gate46inter3));
  inv1  gate1321(.a(s_111), .O(gate46inter4));
  nand2 gate1322(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate1323(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate1324(.a(G6), .O(gate46inter7));
  inv1  gate1325(.a(G272), .O(gate46inter8));
  nand2 gate1326(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate1327(.a(s_111), .b(gate46inter3), .O(gate46inter10));
  nor2  gate1328(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate1329(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate1330(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );

  xor2  gate967(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate968(.a(gate50inter0), .b(s_60), .O(gate50inter1));
  and2  gate969(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate970(.a(s_60), .O(gate50inter3));
  inv1  gate971(.a(s_61), .O(gate50inter4));
  nand2 gate972(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate973(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate974(.a(G10), .O(gate50inter7));
  inv1  gate975(.a(G278), .O(gate50inter8));
  nand2 gate976(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate977(.a(s_61), .b(gate50inter3), .O(gate50inter10));
  nor2  gate978(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate979(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate980(.a(gate50inter12), .b(gate50inter1), .O(G371));
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate1695(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate1696(.a(gate52inter0), .b(s_164), .O(gate52inter1));
  and2  gate1697(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate1698(.a(s_164), .O(gate52inter3));
  inv1  gate1699(.a(s_165), .O(gate52inter4));
  nand2 gate1700(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate1701(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate1702(.a(G12), .O(gate52inter7));
  inv1  gate1703(.a(G281), .O(gate52inter8));
  nand2 gate1704(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate1705(.a(s_165), .b(gate52inter3), .O(gate52inter10));
  nor2  gate1706(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate1707(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate1708(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate1877(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate1878(.a(gate54inter0), .b(s_190), .O(gate54inter1));
  and2  gate1879(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate1880(.a(s_190), .O(gate54inter3));
  inv1  gate1881(.a(s_191), .O(gate54inter4));
  nand2 gate1882(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate1883(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate1884(.a(G14), .O(gate54inter7));
  inv1  gate1885(.a(G284), .O(gate54inter8));
  nand2 gate1886(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate1887(.a(s_191), .b(gate54inter3), .O(gate54inter10));
  nor2  gate1888(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate1889(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate1890(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate2115(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate2116(.a(gate58inter0), .b(s_224), .O(gate58inter1));
  and2  gate2117(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate2118(.a(s_224), .O(gate58inter3));
  inv1  gate2119(.a(s_225), .O(gate58inter4));
  nand2 gate2120(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate2121(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate2122(.a(G18), .O(gate58inter7));
  inv1  gate2123(.a(G290), .O(gate58inter8));
  nand2 gate2124(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate2125(.a(s_225), .b(gate58inter3), .O(gate58inter10));
  nor2  gate2126(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate2127(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate2128(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate589(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate590(.a(gate60inter0), .b(s_6), .O(gate60inter1));
  and2  gate591(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate592(.a(s_6), .O(gate60inter3));
  inv1  gate593(.a(s_7), .O(gate60inter4));
  nand2 gate594(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate595(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate596(.a(G20), .O(gate60inter7));
  inv1  gate597(.a(G293), .O(gate60inter8));
  nand2 gate598(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate599(.a(s_7), .b(gate60inter3), .O(gate60inter10));
  nor2  gate600(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate601(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate602(.a(gate60inter12), .b(gate60inter1), .O(G381));
nand2 gate61( .a(G21), .b(G296), .O(G382) );

  xor2  gate2395(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate2396(.a(gate62inter0), .b(s_264), .O(gate62inter1));
  and2  gate2397(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate2398(.a(s_264), .O(gate62inter3));
  inv1  gate2399(.a(s_265), .O(gate62inter4));
  nand2 gate2400(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate2401(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate2402(.a(G22), .O(gate62inter7));
  inv1  gate2403(.a(G296), .O(gate62inter8));
  nand2 gate2404(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate2405(.a(s_265), .b(gate62inter3), .O(gate62inter10));
  nor2  gate2406(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate2407(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate2408(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );

  xor2  gate2605(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate2606(.a(gate66inter0), .b(s_294), .O(gate66inter1));
  and2  gate2607(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate2608(.a(s_294), .O(gate66inter3));
  inv1  gate2609(.a(s_295), .O(gate66inter4));
  nand2 gate2610(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate2611(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate2612(.a(G26), .O(gate66inter7));
  inv1  gate2613(.a(G302), .O(gate66inter8));
  nand2 gate2614(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate2615(.a(s_295), .b(gate66inter3), .O(gate66inter10));
  nor2  gate2616(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate2617(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate2618(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate1331(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate1332(.a(gate70inter0), .b(s_112), .O(gate70inter1));
  and2  gate1333(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate1334(.a(s_112), .O(gate70inter3));
  inv1  gate1335(.a(s_113), .O(gate70inter4));
  nand2 gate1336(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate1337(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate1338(.a(G30), .O(gate70inter7));
  inv1  gate1339(.a(G308), .O(gate70inter8));
  nand2 gate1340(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate1341(.a(s_113), .b(gate70inter3), .O(gate70inter10));
  nor2  gate1342(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate1343(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate1344(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate1821(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate1822(.a(gate74inter0), .b(s_182), .O(gate74inter1));
  and2  gate1823(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate1824(.a(s_182), .O(gate74inter3));
  inv1  gate1825(.a(s_183), .O(gate74inter4));
  nand2 gate1826(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate1827(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate1828(.a(G5), .O(gate74inter7));
  inv1  gate1829(.a(G314), .O(gate74inter8));
  nand2 gate1830(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate1831(.a(s_183), .b(gate74inter3), .O(gate74inter10));
  nor2  gate1832(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate1833(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate1834(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );

  xor2  gate2227(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate2228(.a(gate76inter0), .b(s_240), .O(gate76inter1));
  and2  gate2229(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate2230(.a(s_240), .O(gate76inter3));
  inv1  gate2231(.a(s_241), .O(gate76inter4));
  nand2 gate2232(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate2233(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate2234(.a(G13), .O(gate76inter7));
  inv1  gate2235(.a(G317), .O(gate76inter8));
  nand2 gate2236(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate2237(.a(s_241), .b(gate76inter3), .O(gate76inter10));
  nor2  gate2238(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate2239(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate2240(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate1275(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate1276(.a(gate82inter0), .b(s_104), .O(gate82inter1));
  and2  gate1277(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate1278(.a(s_104), .O(gate82inter3));
  inv1  gate1279(.a(s_105), .O(gate82inter4));
  nand2 gate1280(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate1281(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate1282(.a(G7), .O(gate82inter7));
  inv1  gate1283(.a(G326), .O(gate82inter8));
  nand2 gate1284(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate1285(.a(s_105), .b(gate82inter3), .O(gate82inter10));
  nor2  gate1286(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate1287(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate1288(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );

  xor2  gate1541(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate1542(.a(gate84inter0), .b(s_142), .O(gate84inter1));
  and2  gate1543(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate1544(.a(s_142), .O(gate84inter3));
  inv1  gate1545(.a(s_143), .O(gate84inter4));
  nand2 gate1546(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate1547(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate1548(.a(G15), .O(gate84inter7));
  inv1  gate1549(.a(G329), .O(gate84inter8));
  nand2 gate1550(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate1551(.a(s_143), .b(gate84inter3), .O(gate84inter10));
  nor2  gate1552(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate1553(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate1554(.a(gate84inter12), .b(gate84inter1), .O(G405));

  xor2  gate1653(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate1654(.a(gate85inter0), .b(s_158), .O(gate85inter1));
  and2  gate1655(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate1656(.a(s_158), .O(gate85inter3));
  inv1  gate1657(.a(s_159), .O(gate85inter4));
  nand2 gate1658(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate1659(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate1660(.a(G4), .O(gate85inter7));
  inv1  gate1661(.a(G332), .O(gate85inter8));
  nand2 gate1662(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate1663(.a(s_159), .b(gate85inter3), .O(gate85inter10));
  nor2  gate1664(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate1665(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate1666(.a(gate85inter12), .b(gate85inter1), .O(G406));

  xor2  gate1709(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate1710(.a(gate86inter0), .b(s_166), .O(gate86inter1));
  and2  gate1711(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate1712(.a(s_166), .O(gate86inter3));
  inv1  gate1713(.a(s_167), .O(gate86inter4));
  nand2 gate1714(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate1715(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate1716(.a(G8), .O(gate86inter7));
  inv1  gate1717(.a(G332), .O(gate86inter8));
  nand2 gate1718(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate1719(.a(s_167), .b(gate86inter3), .O(gate86inter10));
  nor2  gate1720(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate1721(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate1722(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );

  xor2  gate673(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate674(.a(gate89inter0), .b(s_18), .O(gate89inter1));
  and2  gate675(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate676(.a(s_18), .O(gate89inter3));
  inv1  gate677(.a(s_19), .O(gate89inter4));
  nand2 gate678(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate679(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate680(.a(G17), .O(gate89inter7));
  inv1  gate681(.a(G338), .O(gate89inter8));
  nand2 gate682(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate683(.a(s_19), .b(gate89inter3), .O(gate89inter10));
  nor2  gate684(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate685(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate686(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );

  xor2  gate2633(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate2634(.a(gate93inter0), .b(s_298), .O(gate93inter1));
  and2  gate2635(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate2636(.a(s_298), .O(gate93inter3));
  inv1  gate2637(.a(s_299), .O(gate93inter4));
  nand2 gate2638(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate2639(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate2640(.a(G18), .O(gate93inter7));
  inv1  gate2641(.a(G344), .O(gate93inter8));
  nand2 gate2642(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate2643(.a(s_299), .b(gate93inter3), .O(gate93inter10));
  nor2  gate2644(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate2645(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate2646(.a(gate93inter12), .b(gate93inter1), .O(G414));
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate785(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate786(.a(gate95inter0), .b(s_34), .O(gate95inter1));
  and2  gate787(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate788(.a(s_34), .O(gate95inter3));
  inv1  gate789(.a(s_35), .O(gate95inter4));
  nand2 gate790(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate791(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate792(.a(G26), .O(gate95inter7));
  inv1  gate793(.a(G347), .O(gate95inter8));
  nand2 gate794(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate795(.a(s_35), .b(gate95inter3), .O(gate95inter10));
  nor2  gate796(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate797(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate798(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate1373(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate1374(.a(gate98inter0), .b(s_118), .O(gate98inter1));
  and2  gate1375(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate1376(.a(s_118), .O(gate98inter3));
  inv1  gate1377(.a(s_119), .O(gate98inter4));
  nand2 gate1378(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate1379(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate1380(.a(G23), .O(gate98inter7));
  inv1  gate1381(.a(G350), .O(gate98inter8));
  nand2 gate1382(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate1383(.a(s_119), .b(gate98inter3), .O(gate98inter10));
  nor2  gate1384(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate1385(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate1386(.a(gate98inter12), .b(gate98inter1), .O(G419));

  xor2  gate1555(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate1556(.a(gate99inter0), .b(s_144), .O(gate99inter1));
  and2  gate1557(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate1558(.a(s_144), .O(gate99inter3));
  inv1  gate1559(.a(s_145), .O(gate99inter4));
  nand2 gate1560(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate1561(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate1562(.a(G27), .O(gate99inter7));
  inv1  gate1563(.a(G353), .O(gate99inter8));
  nand2 gate1564(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate1565(.a(s_145), .b(gate99inter3), .O(gate99inter10));
  nor2  gate1566(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate1567(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate1568(.a(gate99inter12), .b(gate99inter1), .O(G420));

  xor2  gate1961(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate1962(.a(gate100inter0), .b(s_202), .O(gate100inter1));
  and2  gate1963(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate1964(.a(s_202), .O(gate100inter3));
  inv1  gate1965(.a(s_203), .O(gate100inter4));
  nand2 gate1966(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate1967(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate1968(.a(G31), .O(gate100inter7));
  inv1  gate1969(.a(G353), .O(gate100inter8));
  nand2 gate1970(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate1971(.a(s_203), .b(gate100inter3), .O(gate100inter10));
  nor2  gate1972(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate1973(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate1974(.a(gate100inter12), .b(gate100inter1), .O(G421));

  xor2  gate1345(.a(G356), .b(G20), .O(gate101inter0));
  nand2 gate1346(.a(gate101inter0), .b(s_114), .O(gate101inter1));
  and2  gate1347(.a(G356), .b(G20), .O(gate101inter2));
  inv1  gate1348(.a(s_114), .O(gate101inter3));
  inv1  gate1349(.a(s_115), .O(gate101inter4));
  nand2 gate1350(.a(gate101inter4), .b(gate101inter3), .O(gate101inter5));
  nor2  gate1351(.a(gate101inter5), .b(gate101inter2), .O(gate101inter6));
  inv1  gate1352(.a(G20), .O(gate101inter7));
  inv1  gate1353(.a(G356), .O(gate101inter8));
  nand2 gate1354(.a(gate101inter8), .b(gate101inter7), .O(gate101inter9));
  nand2 gate1355(.a(s_115), .b(gate101inter3), .O(gate101inter10));
  nor2  gate1356(.a(gate101inter10), .b(gate101inter9), .O(gate101inter11));
  nor2  gate1357(.a(gate101inter11), .b(gate101inter6), .O(gate101inter12));
  nand2 gate1358(.a(gate101inter12), .b(gate101inter1), .O(G422));
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );

  xor2  gate2591(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate2592(.a(gate105inter0), .b(s_292), .O(gate105inter1));
  and2  gate2593(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate2594(.a(s_292), .O(gate105inter3));
  inv1  gate2595(.a(s_293), .O(gate105inter4));
  nand2 gate2596(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate2597(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate2598(.a(G362), .O(gate105inter7));
  inv1  gate2599(.a(G363), .O(gate105inter8));
  nand2 gate2600(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate2601(.a(s_293), .b(gate105inter3), .O(gate105inter10));
  nor2  gate2602(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate2603(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate2604(.a(gate105inter12), .b(gate105inter1), .O(G426));

  xor2  gate883(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate884(.a(gate106inter0), .b(s_48), .O(gate106inter1));
  and2  gate885(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate886(.a(s_48), .O(gate106inter3));
  inv1  gate887(.a(s_49), .O(gate106inter4));
  nand2 gate888(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate889(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate890(.a(G364), .O(gate106inter7));
  inv1  gate891(.a(G365), .O(gate106inter8));
  nand2 gate892(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate893(.a(s_49), .b(gate106inter3), .O(gate106inter10));
  nor2  gate894(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate895(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate896(.a(gate106inter12), .b(gate106inter1), .O(G429));

  xor2  gate757(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate758(.a(gate107inter0), .b(s_30), .O(gate107inter1));
  and2  gate759(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate760(.a(s_30), .O(gate107inter3));
  inv1  gate761(.a(s_31), .O(gate107inter4));
  nand2 gate762(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate763(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate764(.a(G366), .O(gate107inter7));
  inv1  gate765(.a(G367), .O(gate107inter8));
  nand2 gate766(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate767(.a(s_31), .b(gate107inter3), .O(gate107inter10));
  nor2  gate768(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate769(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate770(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate1177(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate1178(.a(gate110inter0), .b(s_90), .O(gate110inter1));
  and2  gate1179(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate1180(.a(s_90), .O(gate110inter3));
  inv1  gate1181(.a(s_91), .O(gate110inter4));
  nand2 gate1182(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1183(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1184(.a(G372), .O(gate110inter7));
  inv1  gate1185(.a(G373), .O(gate110inter8));
  nand2 gate1186(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1187(.a(s_91), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1188(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1189(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1190(.a(gate110inter12), .b(gate110inter1), .O(G441));

  xor2  gate2171(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate2172(.a(gate111inter0), .b(s_232), .O(gate111inter1));
  and2  gate2173(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate2174(.a(s_232), .O(gate111inter3));
  inv1  gate2175(.a(s_233), .O(gate111inter4));
  nand2 gate2176(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate2177(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate2178(.a(G374), .O(gate111inter7));
  inv1  gate2179(.a(G375), .O(gate111inter8));
  nand2 gate2180(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate2181(.a(s_233), .b(gate111inter3), .O(gate111inter10));
  nor2  gate2182(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate2183(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate2184(.a(gate111inter12), .b(gate111inter1), .O(G444));
nand2 gate112( .a(G376), .b(G377), .O(G447) );

  xor2  gate743(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate744(.a(gate113inter0), .b(s_28), .O(gate113inter1));
  and2  gate745(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate746(.a(s_28), .O(gate113inter3));
  inv1  gate747(.a(s_29), .O(gate113inter4));
  nand2 gate748(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate749(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate750(.a(G378), .O(gate113inter7));
  inv1  gate751(.a(G379), .O(gate113inter8));
  nand2 gate752(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate753(.a(s_29), .b(gate113inter3), .O(gate113inter10));
  nor2  gate754(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate755(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate756(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate2269(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate2270(.a(gate117inter0), .b(s_246), .O(gate117inter1));
  and2  gate2271(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate2272(.a(s_246), .O(gate117inter3));
  inv1  gate2273(.a(s_247), .O(gate117inter4));
  nand2 gate2274(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate2275(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate2276(.a(G386), .O(gate117inter7));
  inv1  gate2277(.a(G387), .O(gate117inter8));
  nand2 gate2278(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate2279(.a(s_247), .b(gate117inter3), .O(gate117inter10));
  nor2  gate2280(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate2281(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate2282(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );

  xor2  gate1247(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate1248(.a(gate120inter0), .b(s_100), .O(gate120inter1));
  and2  gate1249(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate1250(.a(s_100), .O(gate120inter3));
  inv1  gate1251(.a(s_101), .O(gate120inter4));
  nand2 gate1252(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate1253(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate1254(.a(G392), .O(gate120inter7));
  inv1  gate1255(.a(G393), .O(gate120inter8));
  nand2 gate1256(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate1257(.a(s_101), .b(gate120inter3), .O(gate120inter10));
  nor2  gate1258(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate1259(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate1260(.a(gate120inter12), .b(gate120inter1), .O(G471));
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate2549(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate2550(.a(gate124inter0), .b(s_286), .O(gate124inter1));
  and2  gate2551(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate2552(.a(s_286), .O(gate124inter3));
  inv1  gate2553(.a(s_287), .O(gate124inter4));
  nand2 gate2554(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate2555(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate2556(.a(G400), .O(gate124inter7));
  inv1  gate2557(.a(G401), .O(gate124inter8));
  nand2 gate2558(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate2559(.a(s_287), .b(gate124inter3), .O(gate124inter10));
  nor2  gate2560(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate2561(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate2562(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate2577(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate2578(.a(gate126inter0), .b(s_290), .O(gate126inter1));
  and2  gate2579(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate2580(.a(s_290), .O(gate126inter3));
  inv1  gate2581(.a(s_291), .O(gate126inter4));
  nand2 gate2582(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate2583(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate2584(.a(G404), .O(gate126inter7));
  inv1  gate2585(.a(G405), .O(gate126inter8));
  nand2 gate2586(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate2587(.a(s_291), .b(gate126inter3), .O(gate126inter10));
  nor2  gate2588(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate2589(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate2590(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );

  xor2  gate701(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate702(.a(gate129inter0), .b(s_22), .O(gate129inter1));
  and2  gate703(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate704(.a(s_22), .O(gate129inter3));
  inv1  gate705(.a(s_23), .O(gate129inter4));
  nand2 gate706(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate707(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate708(.a(G410), .O(gate129inter7));
  inv1  gate709(.a(G411), .O(gate129inter8));
  nand2 gate710(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate711(.a(s_23), .b(gate129inter3), .O(gate129inter10));
  nor2  gate712(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate713(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate714(.a(gate129inter12), .b(gate129inter1), .O(G498));
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate1975(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate1976(.a(gate132inter0), .b(s_204), .O(gate132inter1));
  and2  gate1977(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate1978(.a(s_204), .O(gate132inter3));
  inv1  gate1979(.a(s_205), .O(gate132inter4));
  nand2 gate1980(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate1981(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate1982(.a(G416), .O(gate132inter7));
  inv1  gate1983(.a(G417), .O(gate132inter8));
  nand2 gate1984(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate1985(.a(s_205), .b(gate132inter3), .O(gate132inter10));
  nor2  gate1986(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate1987(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate1988(.a(gate132inter12), .b(gate132inter1), .O(G507));

  xor2  gate631(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate632(.a(gate133inter0), .b(s_12), .O(gate133inter1));
  and2  gate633(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate634(.a(s_12), .O(gate133inter3));
  inv1  gate635(.a(s_13), .O(gate133inter4));
  nand2 gate636(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate637(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate638(.a(G418), .O(gate133inter7));
  inv1  gate639(.a(G419), .O(gate133inter8));
  nand2 gate640(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate641(.a(s_13), .b(gate133inter3), .O(gate133inter10));
  nor2  gate642(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate643(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate644(.a(gate133inter12), .b(gate133inter1), .O(G510));
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate2423(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate2424(.a(gate135inter0), .b(s_268), .O(gate135inter1));
  and2  gate2425(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate2426(.a(s_268), .O(gate135inter3));
  inv1  gate2427(.a(s_269), .O(gate135inter4));
  nand2 gate2428(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate2429(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate2430(.a(G422), .O(gate135inter7));
  inv1  gate2431(.a(G423), .O(gate135inter8));
  nand2 gate2432(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate2433(.a(s_269), .b(gate135inter3), .O(gate135inter10));
  nor2  gate2434(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate2435(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate2436(.a(gate135inter12), .b(gate135inter1), .O(G516));
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate1527(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate1528(.a(gate144inter0), .b(s_140), .O(gate144inter1));
  and2  gate1529(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate1530(.a(s_140), .O(gate144inter3));
  inv1  gate1531(.a(s_141), .O(gate144inter4));
  nand2 gate1532(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate1533(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate1534(.a(G468), .O(gate144inter7));
  inv1  gate1535(.a(G471), .O(gate144inter8));
  nand2 gate1536(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate1537(.a(s_141), .b(gate144inter3), .O(gate144inter10));
  nor2  gate1538(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate1539(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate1540(.a(gate144inter12), .b(gate144inter1), .O(G543));

  xor2  gate1583(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate1584(.a(gate145inter0), .b(s_148), .O(gate145inter1));
  and2  gate1585(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate1586(.a(s_148), .O(gate145inter3));
  inv1  gate1587(.a(s_149), .O(gate145inter4));
  nand2 gate1588(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate1589(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate1590(.a(G474), .O(gate145inter7));
  inv1  gate1591(.a(G477), .O(gate145inter8));
  nand2 gate1592(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate1593(.a(s_149), .b(gate145inter3), .O(gate145inter10));
  nor2  gate1594(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate1595(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate1596(.a(gate145inter12), .b(gate145inter1), .O(G546));

  xor2  gate2143(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate2144(.a(gate146inter0), .b(s_228), .O(gate146inter1));
  and2  gate2145(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate2146(.a(s_228), .O(gate146inter3));
  inv1  gate2147(.a(s_229), .O(gate146inter4));
  nand2 gate2148(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate2149(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate2150(.a(G480), .O(gate146inter7));
  inv1  gate2151(.a(G483), .O(gate146inter8));
  nand2 gate2152(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate2153(.a(s_229), .b(gate146inter3), .O(gate146inter10));
  nor2  gate2154(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate2155(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate2156(.a(gate146inter12), .b(gate146inter1), .O(G549));

  xor2  gate2073(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate2074(.a(gate147inter0), .b(s_218), .O(gate147inter1));
  and2  gate2075(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate2076(.a(s_218), .O(gate147inter3));
  inv1  gate2077(.a(s_219), .O(gate147inter4));
  nand2 gate2078(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate2079(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate2080(.a(G486), .O(gate147inter7));
  inv1  gate2081(.a(G489), .O(gate147inter8));
  nand2 gate2082(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate2083(.a(s_219), .b(gate147inter3), .O(gate147inter10));
  nor2  gate2084(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate2085(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate2086(.a(gate147inter12), .b(gate147inter1), .O(G552));

  xor2  gate1387(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1388(.a(gate148inter0), .b(s_120), .O(gate148inter1));
  and2  gate1389(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1390(.a(s_120), .O(gate148inter3));
  inv1  gate1391(.a(s_121), .O(gate148inter4));
  nand2 gate1392(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1393(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1394(.a(G492), .O(gate148inter7));
  inv1  gate1395(.a(G495), .O(gate148inter8));
  nand2 gate1396(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1397(.a(s_121), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1398(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1399(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1400(.a(gate148inter12), .b(gate148inter1), .O(G555));

  xor2  gate995(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate996(.a(gate149inter0), .b(s_64), .O(gate149inter1));
  and2  gate997(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate998(.a(s_64), .O(gate149inter3));
  inv1  gate999(.a(s_65), .O(gate149inter4));
  nand2 gate1000(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate1001(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate1002(.a(G498), .O(gate149inter7));
  inv1  gate1003(.a(G501), .O(gate149inter8));
  nand2 gate1004(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate1005(.a(s_65), .b(gate149inter3), .O(gate149inter10));
  nor2  gate1006(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate1007(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate1008(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate1303(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate1304(.a(gate156inter0), .b(s_108), .O(gate156inter1));
  and2  gate1305(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate1306(.a(s_108), .O(gate156inter3));
  inv1  gate1307(.a(s_109), .O(gate156inter4));
  nand2 gate1308(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate1309(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate1310(.a(G435), .O(gate156inter7));
  inv1  gate1311(.a(G525), .O(gate156inter8));
  nand2 gate1312(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate1313(.a(s_109), .b(gate156inter3), .O(gate156inter10));
  nor2  gate1314(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate1315(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate1316(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate1457(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate1458(.a(gate160inter0), .b(s_130), .O(gate160inter1));
  and2  gate1459(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate1460(.a(s_130), .O(gate160inter3));
  inv1  gate1461(.a(s_131), .O(gate160inter4));
  nand2 gate1462(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate1463(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate1464(.a(G447), .O(gate160inter7));
  inv1  gate1465(.a(G531), .O(gate160inter8));
  nand2 gate1466(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate1467(.a(s_131), .b(gate160inter3), .O(gate160inter10));
  nor2  gate1468(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate1469(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate1470(.a(gate160inter12), .b(gate160inter1), .O(G577));

  xor2  gate2087(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate2088(.a(gate161inter0), .b(s_220), .O(gate161inter1));
  and2  gate2089(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate2090(.a(s_220), .O(gate161inter3));
  inv1  gate2091(.a(s_221), .O(gate161inter4));
  nand2 gate2092(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate2093(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate2094(.a(G450), .O(gate161inter7));
  inv1  gate2095(.a(G534), .O(gate161inter8));
  nand2 gate2096(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate2097(.a(s_221), .b(gate161inter3), .O(gate161inter10));
  nor2  gate2098(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate2099(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate2100(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate617(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate618(.a(gate164inter0), .b(s_10), .O(gate164inter1));
  and2  gate619(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate620(.a(s_10), .O(gate164inter3));
  inv1  gate621(.a(s_11), .O(gate164inter4));
  nand2 gate622(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate623(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate624(.a(G459), .O(gate164inter7));
  inv1  gate625(.a(G537), .O(gate164inter8));
  nand2 gate626(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate627(.a(s_11), .b(gate164inter3), .O(gate164inter10));
  nor2  gate628(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate629(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate630(.a(gate164inter12), .b(gate164inter1), .O(G581));

  xor2  gate603(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate604(.a(gate165inter0), .b(s_8), .O(gate165inter1));
  and2  gate605(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate606(.a(s_8), .O(gate165inter3));
  inv1  gate607(.a(s_9), .O(gate165inter4));
  nand2 gate608(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate609(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate610(.a(G462), .O(gate165inter7));
  inv1  gate611(.a(G540), .O(gate165inter8));
  nand2 gate612(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate613(.a(s_9), .b(gate165inter3), .O(gate165inter10));
  nor2  gate614(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate615(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate616(.a(gate165inter12), .b(gate165inter1), .O(G582));

  xor2  gate2059(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate2060(.a(gate166inter0), .b(s_216), .O(gate166inter1));
  and2  gate2061(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate2062(.a(s_216), .O(gate166inter3));
  inv1  gate2063(.a(s_217), .O(gate166inter4));
  nand2 gate2064(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate2065(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate2066(.a(G465), .O(gate166inter7));
  inv1  gate2067(.a(G540), .O(gate166inter8));
  nand2 gate2068(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate2069(.a(s_217), .b(gate166inter3), .O(gate166inter10));
  nor2  gate2070(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate2071(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate2072(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate2199(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate2200(.a(gate173inter0), .b(s_236), .O(gate173inter1));
  and2  gate2201(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate2202(.a(s_236), .O(gate173inter3));
  inv1  gate2203(.a(s_237), .O(gate173inter4));
  nand2 gate2204(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate2205(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate2206(.a(G486), .O(gate173inter7));
  inv1  gate2207(.a(G552), .O(gate173inter8));
  nand2 gate2208(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate2209(.a(s_237), .b(gate173inter3), .O(gate173inter10));
  nor2  gate2210(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate2211(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate2212(.a(gate173inter12), .b(gate173inter1), .O(G590));

  xor2  gate1849(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate1850(.a(gate174inter0), .b(s_186), .O(gate174inter1));
  and2  gate1851(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate1852(.a(s_186), .O(gate174inter3));
  inv1  gate1853(.a(s_187), .O(gate174inter4));
  nand2 gate1854(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate1855(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate1856(.a(G489), .O(gate174inter7));
  inv1  gate1857(.a(G552), .O(gate174inter8));
  nand2 gate1858(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate1859(.a(s_187), .b(gate174inter3), .O(gate174inter10));
  nor2  gate1860(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate1861(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate1862(.a(gate174inter12), .b(gate174inter1), .O(G591));

  xor2  gate1681(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate1682(.a(gate175inter0), .b(s_162), .O(gate175inter1));
  and2  gate1683(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate1684(.a(s_162), .O(gate175inter3));
  inv1  gate1685(.a(s_163), .O(gate175inter4));
  nand2 gate1686(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1687(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1688(.a(G492), .O(gate175inter7));
  inv1  gate1689(.a(G555), .O(gate175inter8));
  nand2 gate1690(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1691(.a(s_163), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1692(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1693(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1694(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate1933(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1934(.a(gate186inter0), .b(s_198), .O(gate186inter1));
  and2  gate1935(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1936(.a(s_198), .O(gate186inter3));
  inv1  gate1937(.a(s_199), .O(gate186inter4));
  nand2 gate1938(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1939(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1940(.a(G572), .O(gate186inter7));
  inv1  gate1941(.a(G573), .O(gate186inter8));
  nand2 gate1942(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1943(.a(s_199), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1944(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1945(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1946(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );

  xor2  gate2241(.a(G579), .b(G578), .O(gate189inter0));
  nand2 gate2242(.a(gate189inter0), .b(s_242), .O(gate189inter1));
  and2  gate2243(.a(G579), .b(G578), .O(gate189inter2));
  inv1  gate2244(.a(s_242), .O(gate189inter3));
  inv1  gate2245(.a(s_243), .O(gate189inter4));
  nand2 gate2246(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate2247(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate2248(.a(G578), .O(gate189inter7));
  inv1  gate2249(.a(G579), .O(gate189inter8));
  nand2 gate2250(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate2251(.a(s_243), .b(gate189inter3), .O(gate189inter10));
  nor2  gate2252(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate2253(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate2254(.a(gate189inter12), .b(gate189inter1), .O(G622));

  xor2  gate855(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate856(.a(gate190inter0), .b(s_44), .O(gate190inter1));
  and2  gate857(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate858(.a(s_44), .O(gate190inter3));
  inv1  gate859(.a(s_45), .O(gate190inter4));
  nand2 gate860(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate861(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate862(.a(G580), .O(gate190inter7));
  inv1  gate863(.a(G581), .O(gate190inter8));
  nand2 gate864(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate865(.a(s_45), .b(gate190inter3), .O(gate190inter10));
  nor2  gate866(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate867(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate868(.a(gate190inter12), .b(gate190inter1), .O(G627));

  xor2  gate575(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate576(.a(gate191inter0), .b(s_4), .O(gate191inter1));
  and2  gate577(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate578(.a(s_4), .O(gate191inter3));
  inv1  gate579(.a(s_5), .O(gate191inter4));
  nand2 gate580(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate581(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate582(.a(G582), .O(gate191inter7));
  inv1  gate583(.a(G583), .O(gate191inter8));
  nand2 gate584(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate585(.a(s_5), .b(gate191inter3), .O(gate191inter10));
  nor2  gate586(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate587(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate588(.a(gate191inter12), .b(gate191inter1), .O(G632));

  xor2  gate2129(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate2130(.a(gate192inter0), .b(s_226), .O(gate192inter1));
  and2  gate2131(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate2132(.a(s_226), .O(gate192inter3));
  inv1  gate2133(.a(s_227), .O(gate192inter4));
  nand2 gate2134(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate2135(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate2136(.a(G584), .O(gate192inter7));
  inv1  gate2137(.a(G585), .O(gate192inter8));
  nand2 gate2138(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate2139(.a(s_227), .b(gate192inter3), .O(gate192inter10));
  nor2  gate2140(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate2141(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate2142(.a(gate192inter12), .b(gate192inter1), .O(G637));

  xor2  gate1415(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate1416(.a(gate193inter0), .b(s_124), .O(gate193inter1));
  and2  gate1417(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate1418(.a(s_124), .O(gate193inter3));
  inv1  gate1419(.a(s_125), .O(gate193inter4));
  nand2 gate1420(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate1421(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate1422(.a(G586), .O(gate193inter7));
  inv1  gate1423(.a(G587), .O(gate193inter8));
  nand2 gate1424(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate1425(.a(s_125), .b(gate193inter3), .O(gate193inter10));
  nor2  gate1426(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate1427(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate1428(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate1513(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate1514(.a(gate195inter0), .b(s_138), .O(gate195inter1));
  and2  gate1515(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate1516(.a(s_138), .O(gate195inter3));
  inv1  gate1517(.a(s_139), .O(gate195inter4));
  nand2 gate1518(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate1519(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate1520(.a(G590), .O(gate195inter7));
  inv1  gate1521(.a(G591), .O(gate195inter8));
  nand2 gate1522(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate1523(.a(s_139), .b(gate195inter3), .O(gate195inter10));
  nor2  gate1524(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate1525(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate1526(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate1037(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate1038(.a(gate197inter0), .b(s_70), .O(gate197inter1));
  and2  gate1039(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate1040(.a(s_70), .O(gate197inter3));
  inv1  gate1041(.a(s_71), .O(gate197inter4));
  nand2 gate1042(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate1043(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate1044(.a(G594), .O(gate197inter7));
  inv1  gate1045(.a(G595), .O(gate197inter8));
  nand2 gate1046(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate1047(.a(s_71), .b(gate197inter3), .O(gate197inter10));
  nor2  gate1048(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate1049(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate1050(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );

  xor2  gate2213(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate2214(.a(gate200inter0), .b(s_238), .O(gate200inter1));
  and2  gate2215(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate2216(.a(s_238), .O(gate200inter3));
  inv1  gate2217(.a(s_239), .O(gate200inter4));
  nand2 gate2218(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate2219(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate2220(.a(G600), .O(gate200inter7));
  inv1  gate2221(.a(G601), .O(gate200inter8));
  nand2 gate2222(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate2223(.a(s_239), .b(gate200inter3), .O(gate200inter10));
  nor2  gate2224(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate2225(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate2226(.a(gate200inter12), .b(gate200inter1), .O(G663));
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );

  xor2  gate1135(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate1136(.a(gate209inter0), .b(s_84), .O(gate209inter1));
  and2  gate1137(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate1138(.a(s_84), .O(gate209inter3));
  inv1  gate1139(.a(s_85), .O(gate209inter4));
  nand2 gate1140(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate1141(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate1142(.a(G602), .O(gate209inter7));
  inv1  gate1143(.a(G666), .O(gate209inter8));
  nand2 gate1144(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate1145(.a(s_85), .b(gate209inter3), .O(gate209inter10));
  nor2  gate1146(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate1147(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate1148(.a(gate209inter12), .b(gate209inter1), .O(G690));
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );

  xor2  gate1485(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate1486(.a(gate212inter0), .b(s_134), .O(gate212inter1));
  and2  gate1487(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate1488(.a(s_134), .O(gate212inter3));
  inv1  gate1489(.a(s_135), .O(gate212inter4));
  nand2 gate1490(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate1491(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate1492(.a(G617), .O(gate212inter7));
  inv1  gate1493(.a(G669), .O(gate212inter8));
  nand2 gate1494(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate1495(.a(s_135), .b(gate212inter3), .O(gate212inter10));
  nor2  gate1496(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate1497(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate1498(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate659(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate660(.a(gate215inter0), .b(s_16), .O(gate215inter1));
  and2  gate661(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate662(.a(s_16), .O(gate215inter3));
  inv1  gate663(.a(s_17), .O(gate215inter4));
  nand2 gate664(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate665(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate666(.a(G607), .O(gate215inter7));
  inv1  gate667(.a(G675), .O(gate215inter8));
  nand2 gate668(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate669(.a(s_17), .b(gate215inter3), .O(gate215inter10));
  nor2  gate670(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate671(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate672(.a(gate215inter12), .b(gate215inter1), .O(G696));

  xor2  gate1191(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate1192(.a(gate216inter0), .b(s_92), .O(gate216inter1));
  and2  gate1193(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate1194(.a(s_92), .O(gate216inter3));
  inv1  gate1195(.a(s_93), .O(gate216inter4));
  nand2 gate1196(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate1197(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate1198(.a(G617), .O(gate216inter7));
  inv1  gate1199(.a(G675), .O(gate216inter8));
  nand2 gate1200(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate1201(.a(s_93), .b(gate216inter3), .O(gate216inter10));
  nor2  gate1202(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate1203(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate1204(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );

  xor2  gate925(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate926(.a(gate219inter0), .b(s_54), .O(gate219inter1));
  and2  gate927(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate928(.a(s_54), .O(gate219inter3));
  inv1  gate929(.a(s_55), .O(gate219inter4));
  nand2 gate930(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate931(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate932(.a(G632), .O(gate219inter7));
  inv1  gate933(.a(G681), .O(gate219inter8));
  nand2 gate934(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate935(.a(s_55), .b(gate219inter3), .O(gate219inter10));
  nor2  gate936(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate937(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate938(.a(gate219inter12), .b(gate219inter1), .O(G700));

  xor2  gate1261(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate1262(.a(gate220inter0), .b(s_102), .O(gate220inter1));
  and2  gate1263(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate1264(.a(s_102), .O(gate220inter3));
  inv1  gate1265(.a(s_103), .O(gate220inter4));
  nand2 gate1266(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate1267(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate1268(.a(G637), .O(gate220inter7));
  inv1  gate1269(.a(G681), .O(gate220inter8));
  nand2 gate1270(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate1271(.a(s_103), .b(gate220inter3), .O(gate220inter10));
  nor2  gate1272(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate1273(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate1274(.a(gate220inter12), .b(gate220inter1), .O(G701));

  xor2  gate1093(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate1094(.a(gate221inter0), .b(s_78), .O(gate221inter1));
  and2  gate1095(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate1096(.a(s_78), .O(gate221inter3));
  inv1  gate1097(.a(s_79), .O(gate221inter4));
  nand2 gate1098(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate1099(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate1100(.a(G622), .O(gate221inter7));
  inv1  gate1101(.a(G684), .O(gate221inter8));
  nand2 gate1102(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate1103(.a(s_79), .b(gate221inter3), .O(gate221inter10));
  nor2  gate1104(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate1105(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate1106(.a(gate221inter12), .b(gate221inter1), .O(G702));

  xor2  gate1401(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate1402(.a(gate222inter0), .b(s_122), .O(gate222inter1));
  and2  gate1403(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate1404(.a(s_122), .O(gate222inter3));
  inv1  gate1405(.a(s_123), .O(gate222inter4));
  nand2 gate1406(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate1407(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate1408(.a(G632), .O(gate222inter7));
  inv1  gate1409(.a(G684), .O(gate222inter8));
  nand2 gate1410(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate1411(.a(s_123), .b(gate222inter3), .O(gate222inter10));
  nor2  gate1412(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate1413(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate1414(.a(gate222inter12), .b(gate222inter1), .O(G703));

  xor2  gate2101(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate2102(.a(gate223inter0), .b(s_222), .O(gate223inter1));
  and2  gate2103(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate2104(.a(s_222), .O(gate223inter3));
  inv1  gate2105(.a(s_223), .O(gate223inter4));
  nand2 gate2106(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate2107(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate2108(.a(G627), .O(gate223inter7));
  inv1  gate2109(.a(G687), .O(gate223inter8));
  nand2 gate2110(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate2111(.a(s_223), .b(gate223inter3), .O(gate223inter10));
  nor2  gate2112(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate2113(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate2114(.a(gate223inter12), .b(gate223inter1), .O(G704));

  xor2  gate897(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate898(.a(gate224inter0), .b(s_50), .O(gate224inter1));
  and2  gate899(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate900(.a(s_50), .O(gate224inter3));
  inv1  gate901(.a(s_51), .O(gate224inter4));
  nand2 gate902(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate903(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate904(.a(G637), .O(gate224inter7));
  inv1  gate905(.a(G687), .O(gate224inter8));
  nand2 gate906(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate907(.a(s_51), .b(gate224inter3), .O(gate224inter10));
  nor2  gate908(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate909(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate910(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );

  xor2  gate2507(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate2508(.a(gate230inter0), .b(s_280), .O(gate230inter1));
  and2  gate2509(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate2510(.a(s_280), .O(gate230inter3));
  inv1  gate2511(.a(s_281), .O(gate230inter4));
  nand2 gate2512(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate2513(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate2514(.a(G700), .O(gate230inter7));
  inv1  gate2515(.a(G701), .O(gate230inter8));
  nand2 gate2516(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate2517(.a(s_281), .b(gate230inter3), .O(gate230inter10));
  nor2  gate2518(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate2519(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate2520(.a(gate230inter12), .b(gate230inter1), .O(G721));
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate2045(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate2046(.a(gate233inter0), .b(s_214), .O(gate233inter1));
  and2  gate2047(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate2048(.a(s_214), .O(gate233inter3));
  inv1  gate2049(.a(s_215), .O(gate233inter4));
  nand2 gate2050(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate2051(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate2052(.a(G242), .O(gate233inter7));
  inv1  gate2053(.a(G718), .O(gate233inter8));
  nand2 gate2054(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate2055(.a(s_215), .b(gate233inter3), .O(gate233inter10));
  nor2  gate2056(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate2057(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate2058(.a(gate233inter12), .b(gate233inter1), .O(G730));

  xor2  gate827(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate828(.a(gate234inter0), .b(s_40), .O(gate234inter1));
  and2  gate829(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate830(.a(s_40), .O(gate234inter3));
  inv1  gate831(.a(s_41), .O(gate234inter4));
  nand2 gate832(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate833(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate834(.a(G245), .O(gate234inter7));
  inv1  gate835(.a(G721), .O(gate234inter8));
  nand2 gate836(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate837(.a(s_41), .b(gate234inter3), .O(gate234inter10));
  nor2  gate838(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate839(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate840(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate1065(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate1066(.a(gate236inter0), .b(s_74), .O(gate236inter1));
  and2  gate1067(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate1068(.a(s_74), .O(gate236inter3));
  inv1  gate1069(.a(s_75), .O(gate236inter4));
  nand2 gate1070(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate1071(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate1072(.a(G251), .O(gate236inter7));
  inv1  gate1073(.a(G727), .O(gate236inter8));
  nand2 gate1074(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate1075(.a(s_75), .b(gate236inter3), .O(gate236inter10));
  nor2  gate1076(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate1077(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate1078(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate1793(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1794(.a(gate243inter0), .b(s_178), .O(gate243inter1));
  and2  gate1795(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1796(.a(s_178), .O(gate243inter3));
  inv1  gate1797(.a(s_179), .O(gate243inter4));
  nand2 gate1798(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1799(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1800(.a(G245), .O(gate243inter7));
  inv1  gate1801(.a(G733), .O(gate243inter8));
  nand2 gate1802(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1803(.a(s_179), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1804(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1805(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1806(.a(gate243inter12), .b(gate243inter1), .O(G756));

  xor2  gate1751(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate1752(.a(gate244inter0), .b(s_172), .O(gate244inter1));
  and2  gate1753(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate1754(.a(s_172), .O(gate244inter3));
  inv1  gate1755(.a(s_173), .O(gate244inter4));
  nand2 gate1756(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate1757(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate1758(.a(G721), .O(gate244inter7));
  inv1  gate1759(.a(G733), .O(gate244inter8));
  nand2 gate1760(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate1761(.a(s_173), .b(gate244inter3), .O(gate244inter10));
  nor2  gate1762(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate1763(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate1764(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );

  xor2  gate1891(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate1892(.a(gate247inter0), .b(s_192), .O(gate247inter1));
  and2  gate1893(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate1894(.a(s_192), .O(gate247inter3));
  inv1  gate1895(.a(s_193), .O(gate247inter4));
  nand2 gate1896(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate1897(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate1898(.a(G251), .O(gate247inter7));
  inv1  gate1899(.a(G739), .O(gate247inter8));
  nand2 gate1900(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate1901(.a(s_193), .b(gate247inter3), .O(gate247inter10));
  nor2  gate1902(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate1903(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate1904(.a(gate247inter12), .b(gate247inter1), .O(G760));
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate2311(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate2312(.a(gate249inter0), .b(s_252), .O(gate249inter1));
  and2  gate2313(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate2314(.a(s_252), .O(gate249inter3));
  inv1  gate2315(.a(s_253), .O(gate249inter4));
  nand2 gate2316(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate2317(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate2318(.a(G254), .O(gate249inter7));
  inv1  gate2319(.a(G742), .O(gate249inter8));
  nand2 gate2320(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate2321(.a(s_253), .b(gate249inter3), .O(gate249inter10));
  nor2  gate2322(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate2323(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate2324(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );

  xor2  gate2255(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate2256(.a(gate251inter0), .b(s_244), .O(gate251inter1));
  and2  gate2257(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate2258(.a(s_244), .O(gate251inter3));
  inv1  gate2259(.a(s_245), .O(gate251inter4));
  nand2 gate2260(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate2261(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate2262(.a(G257), .O(gate251inter7));
  inv1  gate2263(.a(G745), .O(gate251inter8));
  nand2 gate2264(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate2265(.a(s_245), .b(gate251inter3), .O(gate251inter10));
  nor2  gate2266(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate2267(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate2268(.a(gate251inter12), .b(gate251inter1), .O(G764));
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate953(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate954(.a(gate253inter0), .b(s_58), .O(gate253inter1));
  and2  gate955(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate956(.a(s_58), .O(gate253inter3));
  inv1  gate957(.a(s_59), .O(gate253inter4));
  nand2 gate958(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate959(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate960(.a(G260), .O(gate253inter7));
  inv1  gate961(.a(G748), .O(gate253inter8));
  nand2 gate962(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate963(.a(s_59), .b(gate253inter3), .O(gate253inter10));
  nor2  gate964(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate965(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate966(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );

  xor2  gate799(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate800(.a(gate255inter0), .b(s_36), .O(gate255inter1));
  and2  gate801(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate802(.a(s_36), .O(gate255inter3));
  inv1  gate803(.a(s_37), .O(gate255inter4));
  nand2 gate804(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate805(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate806(.a(G263), .O(gate255inter7));
  inv1  gate807(.a(G751), .O(gate255inter8));
  nand2 gate808(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate809(.a(s_37), .b(gate255inter3), .O(gate255inter10));
  nor2  gate810(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate811(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate812(.a(gate255inter12), .b(gate255inter1), .O(G768));

  xor2  gate2493(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate2494(.a(gate256inter0), .b(s_278), .O(gate256inter1));
  and2  gate2495(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate2496(.a(s_278), .O(gate256inter3));
  inv1  gate2497(.a(s_279), .O(gate256inter4));
  nand2 gate2498(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate2499(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate2500(.a(G715), .O(gate256inter7));
  inv1  gate2501(.a(G751), .O(gate256inter8));
  nand2 gate2502(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate2503(.a(s_279), .b(gate256inter3), .O(gate256inter10));
  nor2  gate2504(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate2505(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate2506(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );

  xor2  gate547(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate548(.a(gate264inter0), .b(s_0), .O(gate264inter1));
  and2  gate549(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate550(.a(s_0), .O(gate264inter3));
  inv1  gate551(.a(s_1), .O(gate264inter4));
  nand2 gate552(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate553(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate554(.a(G768), .O(gate264inter7));
  inv1  gate555(.a(G769), .O(gate264inter8));
  nand2 gate556(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate557(.a(s_1), .b(gate264inter3), .O(gate264inter10));
  nor2  gate558(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate559(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate560(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );

  xor2  gate1863(.a(G773), .b(G645), .O(gate266inter0));
  nand2 gate1864(.a(gate266inter0), .b(s_188), .O(gate266inter1));
  and2  gate1865(.a(G773), .b(G645), .O(gate266inter2));
  inv1  gate1866(.a(s_188), .O(gate266inter3));
  inv1  gate1867(.a(s_189), .O(gate266inter4));
  nand2 gate1868(.a(gate266inter4), .b(gate266inter3), .O(gate266inter5));
  nor2  gate1869(.a(gate266inter5), .b(gate266inter2), .O(gate266inter6));
  inv1  gate1870(.a(G645), .O(gate266inter7));
  inv1  gate1871(.a(G773), .O(gate266inter8));
  nand2 gate1872(.a(gate266inter8), .b(gate266inter7), .O(gate266inter9));
  nand2 gate1873(.a(s_189), .b(gate266inter3), .O(gate266inter10));
  nor2  gate1874(.a(gate266inter10), .b(gate266inter9), .O(gate266inter11));
  nor2  gate1875(.a(gate266inter11), .b(gate266inter6), .O(gate266inter12));
  nand2 gate1876(.a(gate266inter12), .b(gate266inter1), .O(G797));
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate841(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate842(.a(gate268inter0), .b(s_42), .O(gate268inter1));
  and2  gate843(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate844(.a(s_42), .O(gate268inter3));
  inv1  gate845(.a(s_43), .O(gate268inter4));
  nand2 gate846(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate847(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate848(.a(G651), .O(gate268inter7));
  inv1  gate849(.a(G779), .O(gate268inter8));
  nand2 gate850(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate851(.a(s_43), .b(gate268inter3), .O(gate268inter10));
  nor2  gate852(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate853(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate854(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate1499(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate1500(.a(gate270inter0), .b(s_136), .O(gate270inter1));
  and2  gate1501(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate1502(.a(s_136), .O(gate270inter3));
  inv1  gate1503(.a(s_137), .O(gate270inter4));
  nand2 gate1504(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate1505(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate1506(.a(G657), .O(gate270inter7));
  inv1  gate1507(.a(G785), .O(gate270inter8));
  nand2 gate1508(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate1509(.a(s_137), .b(gate270inter3), .O(gate270inter10));
  nor2  gate1510(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate1511(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate1512(.a(gate270inter12), .b(gate270inter1), .O(G809));
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate1107(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate1108(.a(gate272inter0), .b(s_80), .O(gate272inter1));
  and2  gate1109(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate1110(.a(s_80), .O(gate272inter3));
  inv1  gate1111(.a(s_81), .O(gate272inter4));
  nand2 gate1112(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate1113(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate1114(.a(G663), .O(gate272inter7));
  inv1  gate1115(.a(G791), .O(gate272inter8));
  nand2 gate1116(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate1117(.a(s_81), .b(gate272inter3), .O(gate272inter10));
  nor2  gate1118(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate1119(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate1120(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate2325(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate2326(.a(gate286inter0), .b(s_254), .O(gate286inter1));
  and2  gate2327(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate2328(.a(s_254), .O(gate286inter3));
  inv1  gate2329(.a(s_255), .O(gate286inter4));
  nand2 gate2330(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate2331(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate2332(.a(G788), .O(gate286inter7));
  inv1  gate2333(.a(G812), .O(gate286inter8));
  nand2 gate2334(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate2335(.a(s_255), .b(gate286inter3), .O(gate286inter10));
  nor2  gate2336(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate2337(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate2338(.a(gate286inter12), .b(gate286inter1), .O(G831));

  xor2  gate2465(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate2466(.a(gate287inter0), .b(s_274), .O(gate287inter1));
  and2  gate2467(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate2468(.a(s_274), .O(gate287inter3));
  inv1  gate2469(.a(s_275), .O(gate287inter4));
  nand2 gate2470(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate2471(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate2472(.a(G663), .O(gate287inter7));
  inv1  gate2473(.a(G815), .O(gate287inter8));
  nand2 gate2474(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate2475(.a(s_275), .b(gate287inter3), .O(gate287inter10));
  nor2  gate2476(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate2477(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate2478(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate1009(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate1010(.a(gate291inter0), .b(s_66), .O(gate291inter1));
  and2  gate1011(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate1012(.a(s_66), .O(gate291inter3));
  inv1  gate1013(.a(s_67), .O(gate291inter4));
  nand2 gate1014(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate1015(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate1016(.a(G822), .O(gate291inter7));
  inv1  gate1017(.a(G823), .O(gate291inter8));
  nand2 gate1018(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate1019(.a(s_67), .b(gate291inter3), .O(gate291inter10));
  nor2  gate1020(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate1021(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate1022(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate1429(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate1430(.a(gate293inter0), .b(s_126), .O(gate293inter1));
  and2  gate1431(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate1432(.a(s_126), .O(gate293inter3));
  inv1  gate1433(.a(s_127), .O(gate293inter4));
  nand2 gate1434(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate1435(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate1436(.a(G828), .O(gate293inter7));
  inv1  gate1437(.a(G829), .O(gate293inter8));
  nand2 gate1438(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate1439(.a(s_127), .b(gate293inter3), .O(gate293inter10));
  nor2  gate1440(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate1441(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate1442(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate1947(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate1948(.a(gate296inter0), .b(s_200), .O(gate296inter1));
  and2  gate1949(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate1950(.a(s_200), .O(gate296inter3));
  inv1  gate1951(.a(s_201), .O(gate296inter4));
  nand2 gate1952(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate1953(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate1954(.a(G826), .O(gate296inter7));
  inv1  gate1955(.a(G827), .O(gate296inter8));
  nand2 gate1956(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate1957(.a(s_201), .b(gate296inter3), .O(gate296inter10));
  nor2  gate1958(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate1959(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate1960(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate2437(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate2438(.a(gate387inter0), .b(s_270), .O(gate387inter1));
  and2  gate2439(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate2440(.a(s_270), .O(gate387inter3));
  inv1  gate2441(.a(s_271), .O(gate387inter4));
  nand2 gate2442(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate2443(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate2444(.a(G1), .O(gate387inter7));
  inv1  gate2445(.a(G1036), .O(gate387inter8));
  nand2 gate2446(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate2447(.a(s_271), .b(gate387inter3), .O(gate387inter10));
  nor2  gate2448(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate2449(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate2450(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate2535(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate2536(.a(gate395inter0), .b(s_284), .O(gate395inter1));
  and2  gate2537(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate2538(.a(s_284), .O(gate395inter3));
  inv1  gate2539(.a(s_285), .O(gate395inter4));
  nand2 gate2540(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate2541(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate2542(.a(G9), .O(gate395inter7));
  inv1  gate2543(.a(G1060), .O(gate395inter8));
  nand2 gate2544(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate2545(.a(s_285), .b(gate395inter3), .O(gate395inter10));
  nor2  gate2546(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate2547(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate2548(.a(gate395inter12), .b(gate395inter1), .O(G1156));

  xor2  gate2647(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate2648(.a(gate396inter0), .b(s_300), .O(gate396inter1));
  and2  gate2649(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate2650(.a(s_300), .O(gate396inter3));
  inv1  gate2651(.a(s_301), .O(gate396inter4));
  nand2 gate2652(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate2653(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate2654(.a(G10), .O(gate396inter7));
  inv1  gate2655(.a(G1063), .O(gate396inter8));
  nand2 gate2656(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate2657(.a(s_301), .b(gate396inter3), .O(gate396inter10));
  nor2  gate2658(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate2659(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate2660(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate1597(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate1598(.a(gate398inter0), .b(s_150), .O(gate398inter1));
  and2  gate1599(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate1600(.a(s_150), .O(gate398inter3));
  inv1  gate1601(.a(s_151), .O(gate398inter4));
  nand2 gate1602(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate1603(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate1604(.a(G12), .O(gate398inter7));
  inv1  gate1605(.a(G1069), .O(gate398inter8));
  nand2 gate1606(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate1607(.a(s_151), .b(gate398inter3), .O(gate398inter10));
  nor2  gate1608(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate1609(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate1610(.a(gate398inter12), .b(gate398inter1), .O(G1165));
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );

  xor2  gate2353(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate2354(.a(gate412inter0), .b(s_258), .O(gate412inter1));
  and2  gate2355(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate2356(.a(s_258), .O(gate412inter3));
  inv1  gate2357(.a(s_259), .O(gate412inter4));
  nand2 gate2358(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate2359(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate2360(.a(G26), .O(gate412inter7));
  inv1  gate2361(.a(G1111), .O(gate412inter8));
  nand2 gate2362(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate2363(.a(s_259), .b(gate412inter3), .O(gate412inter10));
  nor2  gate2364(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate2365(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate2366(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );

  xor2  gate1835(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate1836(.a(gate414inter0), .b(s_184), .O(gate414inter1));
  and2  gate1837(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate1838(.a(s_184), .O(gate414inter3));
  inv1  gate1839(.a(s_185), .O(gate414inter4));
  nand2 gate1840(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate1841(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate1842(.a(G28), .O(gate414inter7));
  inv1  gate1843(.a(G1117), .O(gate414inter8));
  nand2 gate1844(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate1845(.a(s_185), .b(gate414inter3), .O(gate414inter10));
  nor2  gate1846(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate1847(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate1848(.a(gate414inter12), .b(gate414inter1), .O(G1213));
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );

  xor2  gate1289(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate1290(.a(gate416inter0), .b(s_106), .O(gate416inter1));
  and2  gate1291(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate1292(.a(s_106), .O(gate416inter3));
  inv1  gate1293(.a(s_107), .O(gate416inter4));
  nand2 gate1294(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate1295(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate1296(.a(G30), .O(gate416inter7));
  inv1  gate1297(.a(G1123), .O(gate416inter8));
  nand2 gate1298(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate1299(.a(s_107), .b(gate416inter3), .O(gate416inter10));
  nor2  gate1300(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate1301(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate1302(.a(gate416inter12), .b(gate416inter1), .O(G1219));
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );

  xor2  gate2381(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate2382(.a(gate419inter0), .b(s_262), .O(gate419inter1));
  and2  gate2383(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate2384(.a(s_262), .O(gate419inter3));
  inv1  gate2385(.a(s_263), .O(gate419inter4));
  nand2 gate2386(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate2387(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate2388(.a(G1), .O(gate419inter7));
  inv1  gate2389(.a(G1132), .O(gate419inter8));
  nand2 gate2390(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate2391(.a(s_263), .b(gate419inter3), .O(gate419inter10));
  nor2  gate2392(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate2393(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate2394(.a(gate419inter12), .b(gate419inter1), .O(G1228));
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );

  xor2  gate1023(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate1024(.a(gate426inter0), .b(s_68), .O(gate426inter1));
  and2  gate1025(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate1026(.a(s_68), .O(gate426inter3));
  inv1  gate1027(.a(s_69), .O(gate426inter4));
  nand2 gate1028(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate1029(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate1030(.a(G1045), .O(gate426inter7));
  inv1  gate1031(.a(G1141), .O(gate426inter8));
  nand2 gate1032(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate1033(.a(s_69), .b(gate426inter3), .O(gate426inter10));
  nor2  gate1034(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate1035(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate1036(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate2451(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate2452(.a(gate430inter0), .b(s_272), .O(gate430inter1));
  and2  gate2453(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate2454(.a(s_272), .O(gate430inter3));
  inv1  gate2455(.a(s_273), .O(gate430inter4));
  nand2 gate2456(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate2457(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate2458(.a(G1051), .O(gate430inter7));
  inv1  gate2459(.a(G1147), .O(gate430inter8));
  nand2 gate2460(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate2461(.a(s_273), .b(gate430inter3), .O(gate430inter10));
  nor2  gate2462(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate2463(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate2464(.a(gate430inter12), .b(gate430inter1), .O(G1239));

  xor2  gate1233(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate1234(.a(gate431inter0), .b(s_98), .O(gate431inter1));
  and2  gate1235(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate1236(.a(s_98), .O(gate431inter3));
  inv1  gate1237(.a(s_99), .O(gate431inter4));
  nand2 gate1238(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate1239(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate1240(.a(G7), .O(gate431inter7));
  inv1  gate1241(.a(G1150), .O(gate431inter8));
  nand2 gate1242(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate1243(.a(s_99), .b(gate431inter3), .O(gate431inter10));
  nor2  gate1244(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate1245(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate1246(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate1471(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate1472(.a(gate433inter0), .b(s_132), .O(gate433inter1));
  and2  gate1473(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate1474(.a(s_132), .O(gate433inter3));
  inv1  gate1475(.a(s_133), .O(gate433inter4));
  nand2 gate1476(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate1477(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate1478(.a(G8), .O(gate433inter7));
  inv1  gate1479(.a(G1153), .O(gate433inter8));
  nand2 gate1480(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate1481(.a(s_133), .b(gate433inter3), .O(gate433inter10));
  nor2  gate1482(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate1483(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate1484(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate1919(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate1920(.a(gate435inter0), .b(s_196), .O(gate435inter1));
  and2  gate1921(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate1922(.a(s_196), .O(gate435inter3));
  inv1  gate1923(.a(s_197), .O(gate435inter4));
  nand2 gate1924(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate1925(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate1926(.a(G9), .O(gate435inter7));
  inv1  gate1927(.a(G1156), .O(gate435inter8));
  nand2 gate1928(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate1929(.a(s_197), .b(gate435inter3), .O(gate435inter10));
  nor2  gate1930(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate1931(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate1932(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );

  xor2  gate2409(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate2410(.a(gate438inter0), .b(s_266), .O(gate438inter1));
  and2  gate2411(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate2412(.a(s_266), .O(gate438inter3));
  inv1  gate2413(.a(s_267), .O(gate438inter4));
  nand2 gate2414(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate2415(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate2416(.a(G1063), .O(gate438inter7));
  inv1  gate2417(.a(G1159), .O(gate438inter8));
  nand2 gate2418(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate2419(.a(s_267), .b(gate438inter3), .O(gate438inter10));
  nor2  gate2420(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate2421(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate2422(.a(gate438inter12), .b(gate438inter1), .O(G1247));

  xor2  gate1163(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate1164(.a(gate439inter0), .b(s_88), .O(gate439inter1));
  and2  gate1165(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate1166(.a(s_88), .O(gate439inter3));
  inv1  gate1167(.a(s_89), .O(gate439inter4));
  nand2 gate1168(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate1169(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate1170(.a(G11), .O(gate439inter7));
  inv1  gate1171(.a(G1162), .O(gate439inter8));
  nand2 gate1172(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate1173(.a(s_89), .b(gate439inter3), .O(gate439inter10));
  nor2  gate1174(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate1175(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate1176(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate1205(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate1206(.a(gate445inter0), .b(s_94), .O(gate445inter1));
  and2  gate1207(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate1208(.a(s_94), .O(gate445inter3));
  inv1  gate1209(.a(s_95), .O(gate445inter4));
  nand2 gate1210(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate1211(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate1212(.a(G14), .O(gate445inter7));
  inv1  gate1213(.a(G1171), .O(gate445inter8));
  nand2 gate1214(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate1215(.a(s_95), .b(gate445inter3), .O(gate445inter10));
  nor2  gate1216(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate1217(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate1218(.a(gate445inter12), .b(gate445inter1), .O(G1254));
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );

  xor2  gate1359(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate1360(.a(gate449inter0), .b(s_116), .O(gate449inter1));
  and2  gate1361(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate1362(.a(s_116), .O(gate449inter3));
  inv1  gate1363(.a(s_117), .O(gate449inter4));
  nand2 gate1364(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate1365(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate1366(.a(G16), .O(gate449inter7));
  inv1  gate1367(.a(G1177), .O(gate449inter8));
  nand2 gate1368(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate1369(.a(s_117), .b(gate449inter3), .O(gate449inter10));
  nor2  gate1370(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate1371(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate1372(.a(gate449inter12), .b(gate449inter1), .O(G1258));

  xor2  gate715(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate716(.a(gate450inter0), .b(s_24), .O(gate450inter1));
  and2  gate717(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate718(.a(s_24), .O(gate450inter3));
  inv1  gate719(.a(s_25), .O(gate450inter4));
  nand2 gate720(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate721(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate722(.a(G1081), .O(gate450inter7));
  inv1  gate723(.a(G1177), .O(gate450inter8));
  nand2 gate724(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate725(.a(s_25), .b(gate450inter3), .O(gate450inter10));
  nor2  gate726(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate727(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate728(.a(gate450inter12), .b(gate450inter1), .O(G1259));
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );

  xor2  gate2185(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate2186(.a(gate452inter0), .b(s_234), .O(gate452inter1));
  and2  gate2187(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate2188(.a(s_234), .O(gate452inter3));
  inv1  gate2189(.a(s_235), .O(gate452inter4));
  nand2 gate2190(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate2191(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate2192(.a(G1084), .O(gate452inter7));
  inv1  gate2193(.a(G1180), .O(gate452inter8));
  nand2 gate2194(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate2195(.a(s_235), .b(gate452inter3), .O(gate452inter10));
  nor2  gate2196(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate2197(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate2198(.a(gate452inter12), .b(gate452inter1), .O(G1261));

  xor2  gate729(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate730(.a(gate453inter0), .b(s_26), .O(gate453inter1));
  and2  gate731(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate732(.a(s_26), .O(gate453inter3));
  inv1  gate733(.a(s_27), .O(gate453inter4));
  nand2 gate734(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate735(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate736(.a(G18), .O(gate453inter7));
  inv1  gate737(.a(G1183), .O(gate453inter8));
  nand2 gate738(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate739(.a(s_27), .b(gate453inter3), .O(gate453inter10));
  nor2  gate740(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate741(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate742(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );

  xor2  gate2367(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate2368(.a(gate458inter0), .b(s_260), .O(gate458inter1));
  and2  gate2369(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate2370(.a(s_260), .O(gate458inter3));
  inv1  gate2371(.a(s_261), .O(gate458inter4));
  nand2 gate2372(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate2373(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate2374(.a(G1093), .O(gate458inter7));
  inv1  gate2375(.a(G1189), .O(gate458inter8));
  nand2 gate2376(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate2377(.a(s_261), .b(gate458inter3), .O(gate458inter10));
  nor2  gate2378(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate2379(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate2380(.a(gate458inter12), .b(gate458inter1), .O(G1267));
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );

  xor2  gate939(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate940(.a(gate462inter0), .b(s_56), .O(gate462inter1));
  and2  gate941(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate942(.a(s_56), .O(gate462inter3));
  inv1  gate943(.a(s_57), .O(gate462inter4));
  nand2 gate944(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate945(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate946(.a(G1099), .O(gate462inter7));
  inv1  gate947(.a(G1195), .O(gate462inter8));
  nand2 gate948(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate949(.a(s_57), .b(gate462inter3), .O(gate462inter10));
  nor2  gate950(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate951(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate952(.a(gate462inter12), .b(gate462inter1), .O(G1271));

  xor2  gate1149(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate1150(.a(gate463inter0), .b(s_86), .O(gate463inter1));
  and2  gate1151(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate1152(.a(s_86), .O(gate463inter3));
  inv1  gate1153(.a(s_87), .O(gate463inter4));
  nand2 gate1154(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate1155(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate1156(.a(G23), .O(gate463inter7));
  inv1  gate1157(.a(G1198), .O(gate463inter8));
  nand2 gate1158(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate1159(.a(s_87), .b(gate463inter3), .O(gate463inter10));
  nor2  gate1160(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate1161(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate1162(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );

  xor2  gate1667(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate1668(.a(gate468inter0), .b(s_160), .O(gate468inter1));
  and2  gate1669(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate1670(.a(s_160), .O(gate468inter3));
  inv1  gate1671(.a(s_161), .O(gate468inter4));
  nand2 gate1672(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate1673(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate1674(.a(G1108), .O(gate468inter7));
  inv1  gate1675(.a(G1204), .O(gate468inter8));
  nand2 gate1676(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate1677(.a(s_161), .b(gate468inter3), .O(gate468inter10));
  nor2  gate1678(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate1679(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate1680(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate813(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate814(.a(gate471inter0), .b(s_38), .O(gate471inter1));
  and2  gate815(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate816(.a(s_38), .O(gate471inter3));
  inv1  gate817(.a(s_39), .O(gate471inter4));
  nand2 gate818(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate819(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate820(.a(G27), .O(gate471inter7));
  inv1  gate821(.a(G1210), .O(gate471inter8));
  nand2 gate822(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate823(.a(s_39), .b(gate471inter3), .O(gate471inter10));
  nor2  gate824(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate825(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate826(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate1989(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate1990(.a(gate474inter0), .b(s_206), .O(gate474inter1));
  and2  gate1991(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate1992(.a(s_206), .O(gate474inter3));
  inv1  gate1993(.a(s_207), .O(gate474inter4));
  nand2 gate1994(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate1995(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate1996(.a(G1117), .O(gate474inter7));
  inv1  gate1997(.a(G1213), .O(gate474inter8));
  nand2 gate1998(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate1999(.a(s_207), .b(gate474inter3), .O(gate474inter10));
  nor2  gate2000(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate2001(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate2002(.a(gate474inter12), .b(gate474inter1), .O(G1283));
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate1569(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate1570(.a(gate476inter0), .b(s_146), .O(gate476inter1));
  and2  gate1571(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate1572(.a(s_146), .O(gate476inter3));
  inv1  gate1573(.a(s_147), .O(gate476inter4));
  nand2 gate1574(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate1575(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate1576(.a(G1120), .O(gate476inter7));
  inv1  gate1577(.a(G1216), .O(gate476inter8));
  nand2 gate1578(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate1579(.a(s_147), .b(gate476inter3), .O(gate476inter10));
  nor2  gate1580(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate1581(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate1582(.a(gate476inter12), .b(gate476inter1), .O(G1285));
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );

  xor2  gate1611(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate1612(.a(gate478inter0), .b(s_152), .O(gate478inter1));
  and2  gate1613(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate1614(.a(s_152), .O(gate478inter3));
  inv1  gate1615(.a(s_153), .O(gate478inter4));
  nand2 gate1616(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate1617(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate1618(.a(G1123), .O(gate478inter7));
  inv1  gate1619(.a(G1219), .O(gate478inter8));
  nand2 gate1620(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate1621(.a(s_153), .b(gate478inter3), .O(gate478inter10));
  nor2  gate1622(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate1623(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate1624(.a(gate478inter12), .b(gate478inter1), .O(G1287));

  xor2  gate1905(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate1906(.a(gate479inter0), .b(s_194), .O(gate479inter1));
  and2  gate1907(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate1908(.a(s_194), .O(gate479inter3));
  inv1  gate1909(.a(s_195), .O(gate479inter4));
  nand2 gate1910(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate1911(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate1912(.a(G31), .O(gate479inter7));
  inv1  gate1913(.a(G1222), .O(gate479inter8));
  nand2 gate1914(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate1915(.a(s_195), .b(gate479inter3), .O(gate479inter10));
  nor2  gate1916(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate1917(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate1918(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate2017(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate2018(.a(gate482inter0), .b(s_210), .O(gate482inter1));
  and2  gate2019(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate2020(.a(s_210), .O(gate482inter3));
  inv1  gate2021(.a(s_211), .O(gate482inter4));
  nand2 gate2022(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate2023(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate2024(.a(G1129), .O(gate482inter7));
  inv1  gate2025(.a(G1225), .O(gate482inter8));
  nand2 gate2026(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate2027(.a(s_211), .b(gate482inter3), .O(gate482inter10));
  nor2  gate2028(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate2029(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate2030(.a(gate482inter12), .b(gate482inter1), .O(G1291));
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate2003(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate2004(.a(gate486inter0), .b(s_208), .O(gate486inter1));
  and2  gate2005(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate2006(.a(s_208), .O(gate486inter3));
  inv1  gate2007(.a(s_209), .O(gate486inter4));
  nand2 gate2008(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate2009(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate2010(.a(G1234), .O(gate486inter7));
  inv1  gate2011(.a(G1235), .O(gate486inter8));
  nand2 gate2012(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate2013(.a(s_209), .b(gate486inter3), .O(gate486inter10));
  nor2  gate2014(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate2015(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate2016(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );

  xor2  gate2521(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate2522(.a(gate488inter0), .b(s_282), .O(gate488inter1));
  and2  gate2523(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate2524(.a(s_282), .O(gate488inter3));
  inv1  gate2525(.a(s_283), .O(gate488inter4));
  nand2 gate2526(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate2527(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate2528(.a(G1238), .O(gate488inter7));
  inv1  gate2529(.a(G1239), .O(gate488inter8));
  nand2 gate2530(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate2531(.a(s_283), .b(gate488inter3), .O(gate488inter10));
  nor2  gate2532(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate2533(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate2534(.a(gate488inter12), .b(gate488inter1), .O(G1297));

  xor2  gate1051(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate1052(.a(gate489inter0), .b(s_72), .O(gate489inter1));
  and2  gate1053(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate1054(.a(s_72), .O(gate489inter3));
  inv1  gate1055(.a(s_73), .O(gate489inter4));
  nand2 gate1056(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate1057(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate1058(.a(G1240), .O(gate489inter7));
  inv1  gate1059(.a(G1241), .O(gate489inter8));
  nand2 gate1060(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate1061(.a(s_73), .b(gate489inter3), .O(gate489inter10));
  nor2  gate1062(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate1063(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate1064(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate1443(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate1444(.a(gate492inter0), .b(s_128), .O(gate492inter1));
  and2  gate1445(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate1446(.a(s_128), .O(gate492inter3));
  inv1  gate1447(.a(s_129), .O(gate492inter4));
  nand2 gate1448(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate1449(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate1450(.a(G1246), .O(gate492inter7));
  inv1  gate1451(.a(G1247), .O(gate492inter8));
  nand2 gate1452(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate1453(.a(s_129), .b(gate492inter3), .O(gate492inter10));
  nor2  gate1454(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate1455(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate1456(.a(gate492inter12), .b(gate492inter1), .O(G1301));
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate1723(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate1724(.a(gate494inter0), .b(s_168), .O(gate494inter1));
  and2  gate1725(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate1726(.a(s_168), .O(gate494inter3));
  inv1  gate1727(.a(s_169), .O(gate494inter4));
  nand2 gate1728(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate1729(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate1730(.a(G1250), .O(gate494inter7));
  inv1  gate1731(.a(G1251), .O(gate494inter8));
  nand2 gate1732(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate1733(.a(s_169), .b(gate494inter3), .O(gate494inter10));
  nor2  gate1734(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate1735(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate1736(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );

  xor2  gate1121(.a(G1261), .b(G1260), .O(gate499inter0));
  nand2 gate1122(.a(gate499inter0), .b(s_82), .O(gate499inter1));
  and2  gate1123(.a(G1261), .b(G1260), .O(gate499inter2));
  inv1  gate1124(.a(s_82), .O(gate499inter3));
  inv1  gate1125(.a(s_83), .O(gate499inter4));
  nand2 gate1126(.a(gate499inter4), .b(gate499inter3), .O(gate499inter5));
  nor2  gate1127(.a(gate499inter5), .b(gate499inter2), .O(gate499inter6));
  inv1  gate1128(.a(G1260), .O(gate499inter7));
  inv1  gate1129(.a(G1261), .O(gate499inter8));
  nand2 gate1130(.a(gate499inter8), .b(gate499inter7), .O(gate499inter9));
  nand2 gate1131(.a(s_83), .b(gate499inter3), .O(gate499inter10));
  nor2  gate1132(.a(gate499inter10), .b(gate499inter9), .O(gate499inter11));
  nor2  gate1133(.a(gate499inter11), .b(gate499inter6), .O(gate499inter12));
  nand2 gate1134(.a(gate499inter12), .b(gate499inter1), .O(G1308));

  xor2  gate981(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate982(.a(gate500inter0), .b(s_62), .O(gate500inter1));
  and2  gate983(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate984(.a(s_62), .O(gate500inter3));
  inv1  gate985(.a(s_63), .O(gate500inter4));
  nand2 gate986(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate987(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate988(.a(G1262), .O(gate500inter7));
  inv1  gate989(.a(G1263), .O(gate500inter8));
  nand2 gate990(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate991(.a(s_63), .b(gate500inter3), .O(gate500inter10));
  nor2  gate992(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate993(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate994(.a(gate500inter12), .b(gate500inter1), .O(G1309));
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate771(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate772(.a(gate503inter0), .b(s_32), .O(gate503inter1));
  and2  gate773(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate774(.a(s_32), .O(gate503inter3));
  inv1  gate775(.a(s_33), .O(gate503inter4));
  nand2 gate776(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate777(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate778(.a(G1268), .O(gate503inter7));
  inv1  gate779(.a(G1269), .O(gate503inter8));
  nand2 gate780(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate781(.a(s_33), .b(gate503inter3), .O(gate503inter10));
  nor2  gate782(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate783(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate784(.a(gate503inter12), .b(gate503inter1), .O(G1312));

  xor2  gate2031(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate2032(.a(gate504inter0), .b(s_212), .O(gate504inter1));
  and2  gate2033(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate2034(.a(s_212), .O(gate504inter3));
  inv1  gate2035(.a(s_213), .O(gate504inter4));
  nand2 gate2036(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate2037(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate2038(.a(G1270), .O(gate504inter7));
  inv1  gate2039(.a(G1271), .O(gate504inter8));
  nand2 gate2040(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate2041(.a(s_213), .b(gate504inter3), .O(gate504inter10));
  nor2  gate2042(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate2043(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate2044(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );

  xor2  gate1639(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate1640(.a(gate507inter0), .b(s_156), .O(gate507inter1));
  and2  gate1641(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate1642(.a(s_156), .O(gate507inter3));
  inv1  gate1643(.a(s_157), .O(gate507inter4));
  nand2 gate1644(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate1645(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate1646(.a(G1276), .O(gate507inter7));
  inv1  gate1647(.a(G1277), .O(gate507inter8));
  nand2 gate1648(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate1649(.a(s_157), .b(gate507inter3), .O(gate507inter10));
  nor2  gate1650(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate1651(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate1652(.a(gate507inter12), .b(gate507inter1), .O(G1316));
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate561(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate562(.a(gate509inter0), .b(s_2), .O(gate509inter1));
  and2  gate563(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate564(.a(s_2), .O(gate509inter3));
  inv1  gate565(.a(s_3), .O(gate509inter4));
  nand2 gate566(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate567(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate568(.a(G1280), .O(gate509inter7));
  inv1  gate569(.a(G1281), .O(gate509inter8));
  nand2 gate570(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate571(.a(s_3), .b(gate509inter3), .O(gate509inter10));
  nor2  gate572(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate573(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate574(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate2339(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate2340(.a(gate511inter0), .b(s_256), .O(gate511inter1));
  and2  gate2341(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate2342(.a(s_256), .O(gate511inter3));
  inv1  gate2343(.a(s_257), .O(gate511inter4));
  nand2 gate2344(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate2345(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate2346(.a(G1284), .O(gate511inter7));
  inv1  gate2347(.a(G1285), .O(gate511inter8));
  nand2 gate2348(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate2349(.a(s_257), .b(gate511inter3), .O(gate511inter10));
  nor2  gate2350(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate2351(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate2352(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );

  xor2  gate2479(.a(G1289), .b(G1288), .O(gate513inter0));
  nand2 gate2480(.a(gate513inter0), .b(s_276), .O(gate513inter1));
  and2  gate2481(.a(G1289), .b(G1288), .O(gate513inter2));
  inv1  gate2482(.a(s_276), .O(gate513inter3));
  inv1  gate2483(.a(s_277), .O(gate513inter4));
  nand2 gate2484(.a(gate513inter4), .b(gate513inter3), .O(gate513inter5));
  nor2  gate2485(.a(gate513inter5), .b(gate513inter2), .O(gate513inter6));
  inv1  gate2486(.a(G1288), .O(gate513inter7));
  inv1  gate2487(.a(G1289), .O(gate513inter8));
  nand2 gate2488(.a(gate513inter8), .b(gate513inter7), .O(gate513inter9));
  nand2 gate2489(.a(s_277), .b(gate513inter3), .O(gate513inter10));
  nor2  gate2490(.a(gate513inter10), .b(gate513inter9), .O(gate513inter11));
  nor2  gate2491(.a(gate513inter11), .b(gate513inter6), .O(gate513inter12));
  nand2 gate2492(.a(gate513inter12), .b(gate513inter1), .O(G1322));

  xor2  gate687(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate688(.a(gate514inter0), .b(s_20), .O(gate514inter1));
  and2  gate689(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate690(.a(s_20), .O(gate514inter3));
  inv1  gate691(.a(s_21), .O(gate514inter4));
  nand2 gate692(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate693(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate694(.a(G1290), .O(gate514inter7));
  inv1  gate695(.a(G1291), .O(gate514inter8));
  nand2 gate696(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate697(.a(s_21), .b(gate514inter3), .O(gate514inter10));
  nor2  gate698(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate699(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate700(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule