module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate209inter0, gate209inter1, gate209inter2, gate209inter3, gate209inter4, gate209inter5, gate209inter6, gate209inter7, gate209inter8, gate209inter9, gate209inter10, gate209inter11, gate209inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate289inter0, gate289inter1, gate289inter2, gate289inter3, gate289inter4, gate289inter5, gate289inter6, gate289inter7, gate289inter8, gate289inter9, gate289inter10, gate289inter11, gate289inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate493inter0, gate493inter1, gate493inter2, gate493inter3, gate493inter4, gate493inter5, gate493inter6, gate493inter7, gate493inter8, gate493inter9, gate493inter10, gate493inter11, gate493inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate396inter0, gate396inter1, gate396inter2, gate396inter3, gate396inter4, gate396inter5, gate396inter6, gate396inter7, gate396inter8, gate396inter9, gate396inter10, gate396inter11, gate396inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate194inter0, gate194inter1, gate194inter2, gate194inter3, gate194inter4, gate194inter5, gate194inter6, gate194inter7, gate194inter8, gate194inter9, gate194inter10, gate194inter11, gate194inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate134inter0, gate134inter1, gate134inter2, gate134inter3, gate134inter4, gate134inter5, gate134inter6, gate134inter7, gate134inter8, gate134inter9, gate134inter10, gate134inter11, gate134inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );

  xor2  gate1863(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate1864(.a(gate14inter0), .b(s_188), .O(gate14inter1));
  and2  gate1865(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate1866(.a(s_188), .O(gate14inter3));
  inv1  gate1867(.a(s_189), .O(gate14inter4));
  nand2 gate1868(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate1869(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate1870(.a(G11), .O(gate14inter7));
  inv1  gate1871(.a(G12), .O(gate14inter8));
  nand2 gate1872(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate1873(.a(s_189), .b(gate14inter3), .O(gate14inter10));
  nor2  gate1874(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate1875(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate1876(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate687(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate688(.a(gate21inter0), .b(s_20), .O(gate21inter1));
  and2  gate689(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate690(.a(s_20), .O(gate21inter3));
  inv1  gate691(.a(s_21), .O(gate21inter4));
  nand2 gate692(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate693(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate694(.a(G25), .O(gate21inter7));
  inv1  gate695(.a(G26), .O(gate21inter8));
  nand2 gate696(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate697(.a(s_21), .b(gate21inter3), .O(gate21inter10));
  nor2  gate698(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate699(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate700(.a(gate21inter12), .b(gate21inter1), .O(G302));

  xor2  gate1331(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate1332(.a(gate22inter0), .b(s_112), .O(gate22inter1));
  and2  gate1333(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate1334(.a(s_112), .O(gate22inter3));
  inv1  gate1335(.a(s_113), .O(gate22inter4));
  nand2 gate1336(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate1337(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate1338(.a(G27), .O(gate22inter7));
  inv1  gate1339(.a(G28), .O(gate22inter8));
  nand2 gate1340(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate1341(.a(s_113), .b(gate22inter3), .O(gate22inter10));
  nor2  gate1342(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate1343(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate1344(.a(gate22inter12), .b(gate22inter1), .O(G305));
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate673(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate674(.a(gate24inter0), .b(s_18), .O(gate24inter1));
  and2  gate675(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate676(.a(s_18), .O(gate24inter3));
  inv1  gate677(.a(s_19), .O(gate24inter4));
  nand2 gate678(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate679(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate680(.a(G31), .O(gate24inter7));
  inv1  gate681(.a(G32), .O(gate24inter8));
  nand2 gate682(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate683(.a(s_19), .b(gate24inter3), .O(gate24inter10));
  nor2  gate684(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate685(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate686(.a(gate24inter12), .b(gate24inter1), .O(G311));

  xor2  gate1961(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate1962(.a(gate25inter0), .b(s_202), .O(gate25inter1));
  and2  gate1963(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate1964(.a(s_202), .O(gate25inter3));
  inv1  gate1965(.a(s_203), .O(gate25inter4));
  nand2 gate1966(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate1967(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate1968(.a(G1), .O(gate25inter7));
  inv1  gate1969(.a(G5), .O(gate25inter8));
  nand2 gate1970(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate1971(.a(s_203), .b(gate25inter3), .O(gate25inter10));
  nor2  gate1972(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate1973(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate1974(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate1289(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate1290(.a(gate33inter0), .b(s_106), .O(gate33inter1));
  and2  gate1291(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate1292(.a(s_106), .O(gate33inter3));
  inv1  gate1293(.a(s_107), .O(gate33inter4));
  nand2 gate1294(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate1295(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate1296(.a(G17), .O(gate33inter7));
  inv1  gate1297(.a(G21), .O(gate33inter8));
  nand2 gate1298(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate1299(.a(s_107), .b(gate33inter3), .O(gate33inter10));
  nor2  gate1300(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate1301(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate1302(.a(gate33inter12), .b(gate33inter1), .O(G338));

  xor2  gate1681(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate1682(.a(gate34inter0), .b(s_162), .O(gate34inter1));
  and2  gate1683(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate1684(.a(s_162), .O(gate34inter3));
  inv1  gate1685(.a(s_163), .O(gate34inter4));
  nand2 gate1686(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate1687(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate1688(.a(G25), .O(gate34inter7));
  inv1  gate1689(.a(G29), .O(gate34inter8));
  nand2 gate1690(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate1691(.a(s_163), .b(gate34inter3), .O(gate34inter10));
  nor2  gate1692(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate1693(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate1694(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate1093(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate1094(.a(gate43inter0), .b(s_78), .O(gate43inter1));
  and2  gate1095(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate1096(.a(s_78), .O(gate43inter3));
  inv1  gate1097(.a(s_79), .O(gate43inter4));
  nand2 gate1098(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate1099(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate1100(.a(G3), .O(gate43inter7));
  inv1  gate1101(.a(G269), .O(gate43inter8));
  nand2 gate1102(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate1103(.a(s_79), .b(gate43inter3), .O(gate43inter10));
  nor2  gate1104(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate1105(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate1106(.a(gate43inter12), .b(gate43inter1), .O(G364));
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate561(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate562(.a(gate46inter0), .b(s_2), .O(gate46inter1));
  and2  gate563(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate564(.a(s_2), .O(gate46inter3));
  inv1  gate565(.a(s_3), .O(gate46inter4));
  nand2 gate566(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate567(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate568(.a(G6), .O(gate46inter7));
  inv1  gate569(.a(G272), .O(gate46inter8));
  nand2 gate570(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate571(.a(s_3), .b(gate46inter3), .O(gate46inter10));
  nor2  gate572(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate573(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate574(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );

  xor2  gate1569(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate1570(.a(gate50inter0), .b(s_146), .O(gate50inter1));
  and2  gate1571(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate1572(.a(s_146), .O(gate50inter3));
  inv1  gate1573(.a(s_147), .O(gate50inter4));
  nand2 gate1574(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate1575(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate1576(.a(G10), .O(gate50inter7));
  inv1  gate1577(.a(G278), .O(gate50inter8));
  nand2 gate1578(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate1579(.a(s_147), .b(gate50inter3), .O(gate50inter10));
  nor2  gate1580(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate1581(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate1582(.a(gate50inter12), .b(gate50inter1), .O(G371));

  xor2  gate1443(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate1444(.a(gate51inter0), .b(s_128), .O(gate51inter1));
  and2  gate1445(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate1446(.a(s_128), .O(gate51inter3));
  inv1  gate1447(.a(s_129), .O(gate51inter4));
  nand2 gate1448(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate1449(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate1450(.a(G11), .O(gate51inter7));
  inv1  gate1451(.a(G281), .O(gate51inter8));
  nand2 gate1452(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate1453(.a(s_129), .b(gate51inter3), .O(gate51inter10));
  nor2  gate1454(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate1455(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate1456(.a(gate51inter12), .b(gate51inter1), .O(G372));

  xor2  gate659(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate660(.a(gate52inter0), .b(s_16), .O(gate52inter1));
  and2  gate661(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate662(.a(s_16), .O(gate52inter3));
  inv1  gate663(.a(s_17), .O(gate52inter4));
  nand2 gate664(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate665(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate666(.a(G12), .O(gate52inter7));
  inv1  gate667(.a(G281), .O(gate52inter8));
  nand2 gate668(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate669(.a(s_17), .b(gate52inter3), .O(gate52inter10));
  nor2  gate670(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate671(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate672(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate1233(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate1234(.a(gate54inter0), .b(s_98), .O(gate54inter1));
  and2  gate1235(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate1236(.a(s_98), .O(gate54inter3));
  inv1  gate1237(.a(s_99), .O(gate54inter4));
  nand2 gate1238(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate1239(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate1240(.a(G14), .O(gate54inter7));
  inv1  gate1241(.a(G284), .O(gate54inter8));
  nand2 gate1242(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate1243(.a(s_99), .b(gate54inter3), .O(gate54inter10));
  nor2  gate1244(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate1245(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate1246(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate743(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate744(.a(gate57inter0), .b(s_28), .O(gate57inter1));
  and2  gate745(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate746(.a(s_28), .O(gate57inter3));
  inv1  gate747(.a(s_29), .O(gate57inter4));
  nand2 gate748(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate749(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate750(.a(G17), .O(gate57inter7));
  inv1  gate751(.a(G290), .O(gate57inter8));
  nand2 gate752(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate753(.a(s_29), .b(gate57inter3), .O(gate57inter10));
  nor2  gate754(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate755(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate756(.a(gate57inter12), .b(gate57inter1), .O(G378));
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );

  xor2  gate1653(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate1654(.a(gate68inter0), .b(s_158), .O(gate68inter1));
  and2  gate1655(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate1656(.a(s_158), .O(gate68inter3));
  inv1  gate1657(.a(s_159), .O(gate68inter4));
  nand2 gate1658(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate1659(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate1660(.a(G28), .O(gate68inter7));
  inv1  gate1661(.a(G305), .O(gate68inter8));
  nand2 gate1662(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate1663(.a(s_159), .b(gate68inter3), .O(gate68inter10));
  nor2  gate1664(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate1665(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate1666(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate1625(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate1626(.a(gate70inter0), .b(s_154), .O(gate70inter1));
  and2  gate1627(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate1628(.a(s_154), .O(gate70inter3));
  inv1  gate1629(.a(s_155), .O(gate70inter4));
  nand2 gate1630(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate1631(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate1632(.a(G30), .O(gate70inter7));
  inv1  gate1633(.a(G308), .O(gate70inter8));
  nand2 gate1634(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate1635(.a(s_155), .b(gate70inter3), .O(gate70inter10));
  nor2  gate1636(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate1637(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate1638(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );

  xor2  gate1919(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate1920(.a(gate72inter0), .b(s_196), .O(gate72inter1));
  and2  gate1921(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate1922(.a(s_196), .O(gate72inter3));
  inv1  gate1923(.a(s_197), .O(gate72inter4));
  nand2 gate1924(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate1925(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate1926(.a(G32), .O(gate72inter7));
  inv1  gate1927(.a(G311), .O(gate72inter8));
  nand2 gate1928(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate1929(.a(s_197), .b(gate72inter3), .O(gate72inter10));
  nor2  gate1930(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate1931(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate1932(.a(gate72inter12), .b(gate72inter1), .O(G393));
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate2101(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate2102(.a(gate82inter0), .b(s_222), .O(gate82inter1));
  and2  gate2103(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate2104(.a(s_222), .O(gate82inter3));
  inv1  gate2105(.a(s_223), .O(gate82inter4));
  nand2 gate2106(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate2107(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate2108(.a(G7), .O(gate82inter7));
  inv1  gate2109(.a(G326), .O(gate82inter8));
  nand2 gate2110(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate2111(.a(s_223), .b(gate82inter3), .O(gate82inter10));
  nor2  gate2112(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate2113(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate2114(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );

  xor2  gate953(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate954(.a(gate84inter0), .b(s_58), .O(gate84inter1));
  and2  gate955(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate956(.a(s_58), .O(gate84inter3));
  inv1  gate957(.a(s_59), .O(gate84inter4));
  nand2 gate958(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate959(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate960(.a(G15), .O(gate84inter7));
  inv1  gate961(.a(G329), .O(gate84inter8));
  nand2 gate962(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate963(.a(s_59), .b(gate84inter3), .O(gate84inter10));
  nor2  gate964(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate965(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate966(.a(gate84inter12), .b(gate84inter1), .O(G405));
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate1583(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate1584(.a(gate86inter0), .b(s_148), .O(gate86inter1));
  and2  gate1585(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate1586(.a(s_148), .O(gate86inter3));
  inv1  gate1587(.a(s_149), .O(gate86inter4));
  nand2 gate1588(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate1589(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate1590(.a(G8), .O(gate86inter7));
  inv1  gate1591(.a(G332), .O(gate86inter8));
  nand2 gate1592(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate1593(.a(s_149), .b(gate86inter3), .O(gate86inter10));
  nor2  gate1594(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate1595(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate1596(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );

  xor2  gate2283(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate2284(.a(gate103inter0), .b(s_248), .O(gate103inter1));
  and2  gate2285(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate2286(.a(s_248), .O(gate103inter3));
  inv1  gate2287(.a(s_249), .O(gate103inter4));
  nand2 gate2288(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate2289(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate2290(.a(G28), .O(gate103inter7));
  inv1  gate2291(.a(G359), .O(gate103inter8));
  nand2 gate2292(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate2293(.a(s_249), .b(gate103inter3), .O(gate103inter10));
  nor2  gate2294(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate2295(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate2296(.a(gate103inter12), .b(gate103inter1), .O(G424));
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate883(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate884(.a(gate106inter0), .b(s_48), .O(gate106inter1));
  and2  gate885(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate886(.a(s_48), .O(gate106inter3));
  inv1  gate887(.a(s_49), .O(gate106inter4));
  nand2 gate888(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate889(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate890(.a(G364), .O(gate106inter7));
  inv1  gate891(.a(G365), .O(gate106inter8));
  nand2 gate892(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate893(.a(s_49), .b(gate106inter3), .O(gate106inter10));
  nor2  gate894(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate895(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate896(.a(gate106inter12), .b(gate106inter1), .O(G429));

  xor2  gate1793(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate1794(.a(gate107inter0), .b(s_178), .O(gate107inter1));
  and2  gate1795(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate1796(.a(s_178), .O(gate107inter3));
  inv1  gate1797(.a(s_179), .O(gate107inter4));
  nand2 gate1798(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate1799(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate1800(.a(G366), .O(gate107inter7));
  inv1  gate1801(.a(G367), .O(gate107inter8));
  nand2 gate1802(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate1803(.a(s_179), .b(gate107inter3), .O(gate107inter10));
  nor2  gate1804(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate1805(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate1806(.a(gate107inter12), .b(gate107inter1), .O(G432));

  xor2  gate2087(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate2088(.a(gate108inter0), .b(s_220), .O(gate108inter1));
  and2  gate2089(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate2090(.a(s_220), .O(gate108inter3));
  inv1  gate2091(.a(s_221), .O(gate108inter4));
  nand2 gate2092(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate2093(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate2094(.a(G368), .O(gate108inter7));
  inv1  gate2095(.a(G369), .O(gate108inter8));
  nand2 gate2096(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate2097(.a(s_221), .b(gate108inter3), .O(gate108inter10));
  nor2  gate2098(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate2099(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate2100(.a(gate108inter12), .b(gate108inter1), .O(G435));
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate995(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate996(.a(gate110inter0), .b(s_64), .O(gate110inter1));
  and2  gate997(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate998(.a(s_64), .O(gate110inter3));
  inv1  gate999(.a(s_65), .O(gate110inter4));
  nand2 gate1000(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate1001(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate1002(.a(G372), .O(gate110inter7));
  inv1  gate1003(.a(G373), .O(gate110inter8));
  nand2 gate1004(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate1005(.a(s_65), .b(gate110inter3), .O(gate110inter10));
  nor2  gate1006(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate1007(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate1008(.a(gate110inter12), .b(gate110inter1), .O(G441));
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );

  xor2  gate617(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate618(.a(gate119inter0), .b(s_10), .O(gate119inter1));
  and2  gate619(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate620(.a(s_10), .O(gate119inter3));
  inv1  gate621(.a(s_11), .O(gate119inter4));
  nand2 gate622(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate623(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate624(.a(G390), .O(gate119inter7));
  inv1  gate625(.a(G391), .O(gate119inter8));
  nand2 gate626(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate627(.a(s_11), .b(gate119inter3), .O(gate119inter10));
  nor2  gate628(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate629(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate630(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate1471(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate1472(.a(gate132inter0), .b(s_132), .O(gate132inter1));
  and2  gate1473(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate1474(.a(s_132), .O(gate132inter3));
  inv1  gate1475(.a(s_133), .O(gate132inter4));
  nand2 gate1476(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate1477(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate1478(.a(G416), .O(gate132inter7));
  inv1  gate1479(.a(G417), .O(gate132inter8));
  nand2 gate1480(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate1481(.a(s_133), .b(gate132inter3), .O(gate132inter10));
  nor2  gate1482(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate1483(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate1484(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );

  xor2  gate2297(.a(G421), .b(G420), .O(gate134inter0));
  nand2 gate2298(.a(gate134inter0), .b(s_250), .O(gate134inter1));
  and2  gate2299(.a(G421), .b(G420), .O(gate134inter2));
  inv1  gate2300(.a(s_250), .O(gate134inter3));
  inv1  gate2301(.a(s_251), .O(gate134inter4));
  nand2 gate2302(.a(gate134inter4), .b(gate134inter3), .O(gate134inter5));
  nor2  gate2303(.a(gate134inter5), .b(gate134inter2), .O(gate134inter6));
  inv1  gate2304(.a(G420), .O(gate134inter7));
  inv1  gate2305(.a(G421), .O(gate134inter8));
  nand2 gate2306(.a(gate134inter8), .b(gate134inter7), .O(gate134inter9));
  nand2 gate2307(.a(s_251), .b(gate134inter3), .O(gate134inter10));
  nor2  gate2308(.a(gate134inter10), .b(gate134inter9), .O(gate134inter11));
  nor2  gate2309(.a(gate134inter11), .b(gate134inter6), .O(gate134inter12));
  nand2 gate2310(.a(gate134inter12), .b(gate134inter1), .O(G513));

  xor2  gate1541(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate1542(.a(gate135inter0), .b(s_142), .O(gate135inter1));
  and2  gate1543(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate1544(.a(s_142), .O(gate135inter3));
  inv1  gate1545(.a(s_143), .O(gate135inter4));
  nand2 gate1546(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate1547(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate1548(.a(G422), .O(gate135inter7));
  inv1  gate1549(.a(G423), .O(gate135inter8));
  nand2 gate1550(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate1551(.a(s_143), .b(gate135inter3), .O(gate135inter10));
  nor2  gate1552(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate1553(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate1554(.a(gate135inter12), .b(gate135inter1), .O(G516));

  xor2  gate1807(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate1808(.a(gate136inter0), .b(s_180), .O(gate136inter1));
  and2  gate1809(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate1810(.a(s_180), .O(gate136inter3));
  inv1  gate1811(.a(s_181), .O(gate136inter4));
  nand2 gate1812(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate1813(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate1814(.a(G424), .O(gate136inter7));
  inv1  gate1815(.a(G425), .O(gate136inter8));
  nand2 gate1816(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate1817(.a(s_181), .b(gate136inter3), .O(gate136inter10));
  nor2  gate1818(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate1819(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate1820(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate729(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate730(.a(gate138inter0), .b(s_26), .O(gate138inter1));
  and2  gate731(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate732(.a(s_26), .O(gate138inter3));
  inv1  gate733(.a(s_27), .O(gate138inter4));
  nand2 gate734(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate735(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate736(.a(G432), .O(gate138inter7));
  inv1  gate737(.a(G435), .O(gate138inter8));
  nand2 gate738(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate739(.a(s_27), .b(gate138inter3), .O(gate138inter10));
  nor2  gate740(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate741(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate742(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate1135(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate1136(.a(gate141inter0), .b(s_84), .O(gate141inter1));
  and2  gate1137(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate1138(.a(s_84), .O(gate141inter3));
  inv1  gate1139(.a(s_85), .O(gate141inter4));
  nand2 gate1140(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate1141(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate1142(.a(G450), .O(gate141inter7));
  inv1  gate1143(.a(G453), .O(gate141inter8));
  nand2 gate1144(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate1145(.a(s_85), .b(gate141inter3), .O(gate141inter10));
  nor2  gate1146(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate1147(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate1148(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate967(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate968(.a(gate144inter0), .b(s_60), .O(gate144inter1));
  and2  gate969(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate970(.a(s_60), .O(gate144inter3));
  inv1  gate971(.a(s_61), .O(gate144inter4));
  nand2 gate972(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate973(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate974(.a(G468), .O(gate144inter7));
  inv1  gate975(.a(G471), .O(gate144inter8));
  nand2 gate976(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate977(.a(s_61), .b(gate144inter3), .O(gate144inter10));
  nor2  gate978(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate979(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate980(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate1163(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate1164(.a(gate147inter0), .b(s_88), .O(gate147inter1));
  and2  gate1165(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate1166(.a(s_88), .O(gate147inter3));
  inv1  gate1167(.a(s_89), .O(gate147inter4));
  nand2 gate1168(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate1169(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate1170(.a(G486), .O(gate147inter7));
  inv1  gate1171(.a(G489), .O(gate147inter8));
  nand2 gate1172(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate1173(.a(s_89), .b(gate147inter3), .O(gate147inter10));
  nor2  gate1174(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate1175(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate1176(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate827(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate828(.a(gate151inter0), .b(s_40), .O(gate151inter1));
  and2  gate829(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate830(.a(s_40), .O(gate151inter3));
  inv1  gate831(.a(s_41), .O(gate151inter4));
  nand2 gate832(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate833(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate834(.a(G510), .O(gate151inter7));
  inv1  gate835(.a(G513), .O(gate151inter8));
  nand2 gate836(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate837(.a(s_41), .b(gate151inter3), .O(gate151inter10));
  nor2  gate838(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate839(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate840(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate1303(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate1304(.a(gate157inter0), .b(s_108), .O(gate157inter1));
  and2  gate1305(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate1306(.a(s_108), .O(gate157inter3));
  inv1  gate1307(.a(s_109), .O(gate157inter4));
  nand2 gate1308(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate1309(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate1310(.a(G438), .O(gate157inter7));
  inv1  gate1311(.a(G528), .O(gate157inter8));
  nand2 gate1312(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate1313(.a(s_109), .b(gate157inter3), .O(gate157inter10));
  nor2  gate1314(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate1315(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate1316(.a(gate157inter12), .b(gate157inter1), .O(G574));
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate813(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate814(.a(gate162inter0), .b(s_38), .O(gate162inter1));
  and2  gate815(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate816(.a(s_38), .O(gate162inter3));
  inv1  gate817(.a(s_39), .O(gate162inter4));
  nand2 gate818(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate819(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate820(.a(G453), .O(gate162inter7));
  inv1  gate821(.a(G534), .O(gate162inter8));
  nand2 gate822(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate823(.a(s_39), .b(gate162inter3), .O(gate162inter10));
  nor2  gate824(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate825(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate826(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate1639(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate1640(.a(gate165inter0), .b(s_156), .O(gate165inter1));
  and2  gate1641(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate1642(.a(s_156), .O(gate165inter3));
  inv1  gate1643(.a(s_157), .O(gate165inter4));
  nand2 gate1644(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate1645(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate1646(.a(G462), .O(gate165inter7));
  inv1  gate1647(.a(G540), .O(gate165inter8));
  nand2 gate1648(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate1649(.a(s_157), .b(gate165inter3), .O(gate165inter10));
  nor2  gate1650(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate1651(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate1652(.a(gate165inter12), .b(gate165inter1), .O(G582));

  xor2  gate1275(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate1276(.a(gate166inter0), .b(s_104), .O(gate166inter1));
  and2  gate1277(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate1278(.a(s_104), .O(gate166inter3));
  inv1  gate1279(.a(s_105), .O(gate166inter4));
  nand2 gate1280(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate1281(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate1282(.a(G465), .O(gate166inter7));
  inv1  gate1283(.a(G540), .O(gate166inter8));
  nand2 gate1284(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate1285(.a(s_105), .b(gate166inter3), .O(gate166inter10));
  nor2  gate1286(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate1287(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate1288(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );

  xor2  gate715(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate716(.a(gate168inter0), .b(s_24), .O(gate168inter1));
  and2  gate717(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate718(.a(s_24), .O(gate168inter3));
  inv1  gate719(.a(s_25), .O(gate168inter4));
  nand2 gate720(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate721(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate722(.a(G471), .O(gate168inter7));
  inv1  gate723(.a(G543), .O(gate168inter8));
  nand2 gate724(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate725(.a(s_25), .b(gate168inter3), .O(gate168inter10));
  nor2  gate726(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate727(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate728(.a(gate168inter12), .b(gate168inter1), .O(G585));

  xor2  gate1751(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate1752(.a(gate169inter0), .b(s_172), .O(gate169inter1));
  and2  gate1753(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate1754(.a(s_172), .O(gate169inter3));
  inv1  gate1755(.a(s_173), .O(gate169inter4));
  nand2 gate1756(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate1757(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate1758(.a(G474), .O(gate169inter7));
  inv1  gate1759(.a(G546), .O(gate169inter8));
  nand2 gate1760(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate1761(.a(s_173), .b(gate169inter3), .O(gate169inter10));
  nor2  gate1762(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate1763(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate1764(.a(gate169inter12), .b(gate169inter1), .O(G586));

  xor2  gate1345(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate1346(.a(gate170inter0), .b(s_114), .O(gate170inter1));
  and2  gate1347(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate1348(.a(s_114), .O(gate170inter3));
  inv1  gate1349(.a(s_115), .O(gate170inter4));
  nand2 gate1350(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate1351(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate1352(.a(G477), .O(gate170inter7));
  inv1  gate1353(.a(G546), .O(gate170inter8));
  nand2 gate1354(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate1355(.a(s_115), .b(gate170inter3), .O(gate170inter10));
  nor2  gate1356(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate1357(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate1358(.a(gate170inter12), .b(gate170inter1), .O(G587));

  xor2  gate1205(.a(G549), .b(G480), .O(gate171inter0));
  nand2 gate1206(.a(gate171inter0), .b(s_94), .O(gate171inter1));
  and2  gate1207(.a(G549), .b(G480), .O(gate171inter2));
  inv1  gate1208(.a(s_94), .O(gate171inter3));
  inv1  gate1209(.a(s_95), .O(gate171inter4));
  nand2 gate1210(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate1211(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate1212(.a(G480), .O(gate171inter7));
  inv1  gate1213(.a(G549), .O(gate171inter8));
  nand2 gate1214(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate1215(.a(s_95), .b(gate171inter3), .O(gate171inter10));
  nor2  gate1216(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate1217(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate1218(.a(gate171inter12), .b(gate171inter1), .O(G588));

  xor2  gate589(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate590(.a(gate172inter0), .b(s_6), .O(gate172inter1));
  and2  gate591(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate592(.a(s_6), .O(gate172inter3));
  inv1  gate593(.a(s_7), .O(gate172inter4));
  nand2 gate594(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate595(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate596(.a(G483), .O(gate172inter7));
  inv1  gate597(.a(G549), .O(gate172inter8));
  nand2 gate598(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate599(.a(s_7), .b(gate172inter3), .O(gate172inter10));
  nor2  gate600(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate601(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate602(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );

  xor2  gate785(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate786(.a(gate176inter0), .b(s_34), .O(gate176inter1));
  and2  gate787(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate788(.a(s_34), .O(gate176inter3));
  inv1  gate789(.a(s_35), .O(gate176inter4));
  nand2 gate790(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate791(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate792(.a(G495), .O(gate176inter7));
  inv1  gate793(.a(G555), .O(gate176inter8));
  nand2 gate794(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate795(.a(s_35), .b(gate176inter3), .O(gate176inter10));
  nor2  gate796(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate797(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate798(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );

  xor2  gate799(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate800(.a(gate184inter0), .b(s_36), .O(gate184inter1));
  and2  gate801(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate802(.a(s_36), .O(gate184inter3));
  inv1  gate803(.a(s_37), .O(gate184inter4));
  nand2 gate804(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate805(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate806(.a(G519), .O(gate184inter7));
  inv1  gate807(.a(G567), .O(gate184inter8));
  nand2 gate808(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate809(.a(s_37), .b(gate184inter3), .O(gate184inter10));
  nor2  gate810(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate811(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate812(.a(gate184inter12), .b(gate184inter1), .O(G601));
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate1555(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate1556(.a(gate193inter0), .b(s_144), .O(gate193inter1));
  and2  gate1557(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate1558(.a(s_144), .O(gate193inter3));
  inv1  gate1559(.a(s_145), .O(gate193inter4));
  nand2 gate1560(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate1561(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate1562(.a(G586), .O(gate193inter7));
  inv1  gate1563(.a(G587), .O(gate193inter8));
  nand2 gate1564(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate1565(.a(s_145), .b(gate193inter3), .O(gate193inter10));
  nor2  gate1566(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate1567(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate1568(.a(gate193inter12), .b(gate193inter1), .O(G642));

  xor2  gate2143(.a(G589), .b(G588), .O(gate194inter0));
  nand2 gate2144(.a(gate194inter0), .b(s_228), .O(gate194inter1));
  and2  gate2145(.a(G589), .b(G588), .O(gate194inter2));
  inv1  gate2146(.a(s_228), .O(gate194inter3));
  inv1  gate2147(.a(s_229), .O(gate194inter4));
  nand2 gate2148(.a(gate194inter4), .b(gate194inter3), .O(gate194inter5));
  nor2  gate2149(.a(gate194inter5), .b(gate194inter2), .O(gate194inter6));
  inv1  gate2150(.a(G588), .O(gate194inter7));
  inv1  gate2151(.a(G589), .O(gate194inter8));
  nand2 gate2152(.a(gate194inter8), .b(gate194inter7), .O(gate194inter9));
  nand2 gate2153(.a(s_229), .b(gate194inter3), .O(gate194inter10));
  nor2  gate2154(.a(gate194inter10), .b(gate194inter9), .O(gate194inter11));
  nor2  gate2155(.a(gate194inter11), .b(gate194inter6), .O(gate194inter12));
  nand2 gate2156(.a(gate194inter12), .b(gate194inter1), .O(G645));
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate1779(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate1780(.a(gate196inter0), .b(s_176), .O(gate196inter1));
  and2  gate1781(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate1782(.a(s_176), .O(gate196inter3));
  inv1  gate1783(.a(s_177), .O(gate196inter4));
  nand2 gate1784(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate1785(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate1786(.a(G592), .O(gate196inter7));
  inv1  gate1787(.a(G593), .O(gate196inter8));
  nand2 gate1788(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate1789(.a(s_177), .b(gate196inter3), .O(gate196inter10));
  nor2  gate1790(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate1791(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate1792(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate1527(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate1528(.a(gate198inter0), .b(s_140), .O(gate198inter1));
  and2  gate1529(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate1530(.a(s_140), .O(gate198inter3));
  inv1  gate1531(.a(s_141), .O(gate198inter4));
  nand2 gate1532(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate1533(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate1534(.a(G596), .O(gate198inter7));
  inv1  gate1535(.a(G597), .O(gate198inter8));
  nand2 gate1536(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate1537(.a(s_141), .b(gate198inter3), .O(gate198inter10));
  nor2  gate1538(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate1539(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate1540(.a(gate198inter12), .b(gate198inter1), .O(G657));

  xor2  gate911(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate912(.a(gate199inter0), .b(s_52), .O(gate199inter1));
  and2  gate913(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate914(.a(s_52), .O(gate199inter3));
  inv1  gate915(.a(s_53), .O(gate199inter4));
  nand2 gate916(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate917(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate918(.a(G598), .O(gate199inter7));
  inv1  gate919(.a(G599), .O(gate199inter8));
  nand2 gate920(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate921(.a(s_53), .b(gate199inter3), .O(gate199inter10));
  nor2  gate922(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate923(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate924(.a(gate199inter12), .b(gate199inter1), .O(G660));

  xor2  gate2241(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate2242(.a(gate200inter0), .b(s_242), .O(gate200inter1));
  and2  gate2243(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate2244(.a(s_242), .O(gate200inter3));
  inv1  gate2245(.a(s_243), .O(gate200inter4));
  nand2 gate2246(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate2247(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate2248(.a(G600), .O(gate200inter7));
  inv1  gate2249(.a(G601), .O(gate200inter8));
  nand2 gate2250(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate2251(.a(s_243), .b(gate200inter3), .O(gate200inter10));
  nor2  gate2252(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate2253(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate2254(.a(gate200inter12), .b(gate200inter1), .O(G663));
nand2 gate201( .a(G602), .b(G607), .O(G666) );

  xor2  gate1023(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate1024(.a(gate202inter0), .b(s_68), .O(gate202inter1));
  and2  gate1025(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate1026(.a(s_68), .O(gate202inter3));
  inv1  gate1027(.a(s_69), .O(gate202inter4));
  nand2 gate1028(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate1029(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate1030(.a(G612), .O(gate202inter7));
  inv1  gate1031(.a(G617), .O(gate202inter8));
  nand2 gate1032(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate1033(.a(s_69), .b(gate202inter3), .O(gate202inter10));
  nor2  gate1034(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate1035(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate1036(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate1821(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate1822(.a(gate205inter0), .b(s_182), .O(gate205inter1));
  and2  gate1823(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate1824(.a(s_182), .O(gate205inter3));
  inv1  gate1825(.a(s_183), .O(gate205inter4));
  nand2 gate1826(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate1827(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate1828(.a(G622), .O(gate205inter7));
  inv1  gate1829(.a(G627), .O(gate205inter8));
  nand2 gate1830(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate1831(.a(s_183), .b(gate205inter3), .O(gate205inter10));
  nor2  gate1832(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate1833(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate1834(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );

  xor2  gate897(.a(G666), .b(G602), .O(gate209inter0));
  nand2 gate898(.a(gate209inter0), .b(s_50), .O(gate209inter1));
  and2  gate899(.a(G666), .b(G602), .O(gate209inter2));
  inv1  gate900(.a(s_50), .O(gate209inter3));
  inv1  gate901(.a(s_51), .O(gate209inter4));
  nand2 gate902(.a(gate209inter4), .b(gate209inter3), .O(gate209inter5));
  nor2  gate903(.a(gate209inter5), .b(gate209inter2), .O(gate209inter6));
  inv1  gate904(.a(G602), .O(gate209inter7));
  inv1  gate905(.a(G666), .O(gate209inter8));
  nand2 gate906(.a(gate209inter8), .b(gate209inter7), .O(gate209inter9));
  nand2 gate907(.a(s_51), .b(gate209inter3), .O(gate209inter10));
  nor2  gate908(.a(gate209inter10), .b(gate209inter9), .O(gate209inter11));
  nor2  gate909(.a(gate209inter11), .b(gate209inter6), .O(gate209inter12));
  nand2 gate910(.a(gate209inter12), .b(gate209inter1), .O(G690));
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate2227(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate2228(.a(gate211inter0), .b(s_240), .O(gate211inter1));
  and2  gate2229(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate2230(.a(s_240), .O(gate211inter3));
  inv1  gate2231(.a(s_241), .O(gate211inter4));
  nand2 gate2232(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate2233(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate2234(.a(G612), .O(gate211inter7));
  inv1  gate2235(.a(G669), .O(gate211inter8));
  nand2 gate2236(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate2237(.a(s_241), .b(gate211inter3), .O(gate211inter10));
  nor2  gate2238(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate2239(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate2240(.a(gate211inter12), .b(gate211inter1), .O(G692));

  xor2  gate1611(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate1612(.a(gate212inter0), .b(s_152), .O(gate212inter1));
  and2  gate1613(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate1614(.a(s_152), .O(gate212inter3));
  inv1  gate1615(.a(s_153), .O(gate212inter4));
  nand2 gate1616(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate1617(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate1618(.a(G617), .O(gate212inter7));
  inv1  gate1619(.a(G669), .O(gate212inter8));
  nand2 gate1620(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate1621(.a(s_153), .b(gate212inter3), .O(gate212inter10));
  nor2  gate1622(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate1623(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate1624(.a(gate212inter12), .b(gate212inter1), .O(G693));

  xor2  gate1247(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate1248(.a(gate213inter0), .b(s_100), .O(gate213inter1));
  and2  gate1249(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate1250(.a(s_100), .O(gate213inter3));
  inv1  gate1251(.a(s_101), .O(gate213inter4));
  nand2 gate1252(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate1253(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate1254(.a(G602), .O(gate213inter7));
  inv1  gate1255(.a(G672), .O(gate213inter8));
  nand2 gate1256(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate1257(.a(s_101), .b(gate213inter3), .O(gate213inter10));
  nor2  gate1258(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate1259(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate1260(.a(gate213inter12), .b(gate213inter1), .O(G694));

  xor2  gate2199(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate2200(.a(gate214inter0), .b(s_236), .O(gate214inter1));
  and2  gate2201(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate2202(.a(s_236), .O(gate214inter3));
  inv1  gate2203(.a(s_237), .O(gate214inter4));
  nand2 gate2204(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate2205(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate2206(.a(G612), .O(gate214inter7));
  inv1  gate2207(.a(G672), .O(gate214inter8));
  nand2 gate2208(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate2209(.a(s_237), .b(gate214inter3), .O(gate214inter10));
  nor2  gate2210(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate2211(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate2212(.a(gate214inter12), .b(gate214inter1), .O(G695));

  xor2  gate2031(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate2032(.a(gate215inter0), .b(s_212), .O(gate215inter1));
  and2  gate2033(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate2034(.a(s_212), .O(gate215inter3));
  inv1  gate2035(.a(s_213), .O(gate215inter4));
  nand2 gate2036(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate2037(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate2038(.a(G607), .O(gate215inter7));
  inv1  gate2039(.a(G675), .O(gate215inter8));
  nand2 gate2040(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate2041(.a(s_213), .b(gate215inter3), .O(gate215inter10));
  nor2  gate2042(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate2043(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate2044(.a(gate215inter12), .b(gate215inter1), .O(G696));
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate771(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate772(.a(gate218inter0), .b(s_32), .O(gate218inter1));
  and2  gate773(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate774(.a(s_32), .O(gate218inter3));
  inv1  gate775(.a(s_33), .O(gate218inter4));
  nand2 gate776(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate777(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate778(.a(G627), .O(gate218inter7));
  inv1  gate779(.a(G678), .O(gate218inter8));
  nand2 gate780(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate781(.a(s_33), .b(gate218inter3), .O(gate218inter10));
  nor2  gate782(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate783(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate784(.a(gate218inter12), .b(gate218inter1), .O(G699));

  xor2  gate1695(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate1696(.a(gate219inter0), .b(s_164), .O(gate219inter1));
  and2  gate1697(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate1698(.a(s_164), .O(gate219inter3));
  inv1  gate1699(.a(s_165), .O(gate219inter4));
  nand2 gate1700(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate1701(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate1702(.a(G632), .O(gate219inter7));
  inv1  gate1703(.a(G681), .O(gate219inter8));
  nand2 gate1704(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate1705(.a(s_165), .b(gate219inter3), .O(gate219inter10));
  nor2  gate1706(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate1707(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate1708(.a(gate219inter12), .b(gate219inter1), .O(G700));

  xor2  gate1177(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate1178(.a(gate220inter0), .b(s_90), .O(gate220inter1));
  and2  gate1179(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate1180(.a(s_90), .O(gate220inter3));
  inv1  gate1181(.a(s_91), .O(gate220inter4));
  nand2 gate1182(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate1183(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate1184(.a(G637), .O(gate220inter7));
  inv1  gate1185(.a(G681), .O(gate220inter8));
  nand2 gate1186(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate1187(.a(s_91), .b(gate220inter3), .O(gate220inter10));
  nor2  gate1188(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate1189(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate1190(.a(gate220inter12), .b(gate220inter1), .O(G701));

  xor2  gate1401(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate1402(.a(gate221inter0), .b(s_122), .O(gate221inter1));
  and2  gate1403(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate1404(.a(s_122), .O(gate221inter3));
  inv1  gate1405(.a(s_123), .O(gate221inter4));
  nand2 gate1406(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate1407(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate1408(.a(G622), .O(gate221inter7));
  inv1  gate1409(.a(G684), .O(gate221inter8));
  nand2 gate1410(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate1411(.a(s_123), .b(gate221inter3), .O(gate221inter10));
  nor2  gate1412(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate1413(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate1414(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );

  xor2  gate1513(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate1514(.a(gate226inter0), .b(s_138), .O(gate226inter1));
  and2  gate1515(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate1516(.a(s_138), .O(gate226inter3));
  inv1  gate1517(.a(s_139), .O(gate226inter4));
  nand2 gate1518(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate1519(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate1520(.a(G692), .O(gate226inter7));
  inv1  gate1521(.a(G693), .O(gate226inter8));
  nand2 gate1522(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate1523(.a(s_139), .b(gate226inter3), .O(gate226inter10));
  nor2  gate1524(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate1525(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate1526(.a(gate226inter12), .b(gate226inter1), .O(G709));

  xor2  gate1051(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate1052(.a(gate227inter0), .b(s_72), .O(gate227inter1));
  and2  gate1053(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate1054(.a(s_72), .O(gate227inter3));
  inv1  gate1055(.a(s_73), .O(gate227inter4));
  nand2 gate1056(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate1057(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate1058(.a(G694), .O(gate227inter7));
  inv1  gate1059(.a(G695), .O(gate227inter8));
  nand2 gate1060(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate1061(.a(s_73), .b(gate227inter3), .O(gate227inter10));
  nor2  gate1062(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate1063(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate1064(.a(gate227inter12), .b(gate227inter1), .O(G712));
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate1485(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate1486(.a(gate233inter0), .b(s_134), .O(gate233inter1));
  and2  gate1487(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate1488(.a(s_134), .O(gate233inter3));
  inv1  gate1489(.a(s_135), .O(gate233inter4));
  nand2 gate1490(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate1491(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate1492(.a(G242), .O(gate233inter7));
  inv1  gate1493(.a(G718), .O(gate233inter8));
  nand2 gate1494(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate1495(.a(s_135), .b(gate233inter3), .O(gate233inter10));
  nor2  gate1496(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate1497(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate1498(.a(gate233inter12), .b(gate233inter1), .O(G730));

  xor2  gate1387(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate1388(.a(gate234inter0), .b(s_120), .O(gate234inter1));
  and2  gate1389(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate1390(.a(s_120), .O(gate234inter3));
  inv1  gate1391(.a(s_121), .O(gate234inter4));
  nand2 gate1392(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1393(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1394(.a(G245), .O(gate234inter7));
  inv1  gate1395(.a(G721), .O(gate234inter8));
  nand2 gate1396(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1397(.a(s_121), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1398(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1399(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1400(.a(gate234inter12), .b(gate234inter1), .O(G733));

  xor2  gate1947(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate1948(.a(gate235inter0), .b(s_200), .O(gate235inter1));
  and2  gate1949(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate1950(.a(s_200), .O(gate235inter3));
  inv1  gate1951(.a(s_201), .O(gate235inter4));
  nand2 gate1952(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate1953(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate1954(.a(G248), .O(gate235inter7));
  inv1  gate1955(.a(G724), .O(gate235inter8));
  nand2 gate1956(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate1957(.a(s_201), .b(gate235inter3), .O(gate235inter10));
  nor2  gate1958(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate1959(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate1960(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate1891(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate1892(.a(gate237inter0), .b(s_192), .O(gate237inter1));
  and2  gate1893(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate1894(.a(s_192), .O(gate237inter3));
  inv1  gate1895(.a(s_193), .O(gate237inter4));
  nand2 gate1896(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1897(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1898(.a(G254), .O(gate237inter7));
  inv1  gate1899(.a(G706), .O(gate237inter8));
  nand2 gate1900(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1901(.a(s_193), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1902(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1903(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1904(.a(gate237inter12), .b(gate237inter1), .O(G742));

  xor2  gate645(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate646(.a(gate238inter0), .b(s_14), .O(gate238inter1));
  and2  gate647(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate648(.a(s_14), .O(gate238inter3));
  inv1  gate649(.a(s_15), .O(gate238inter4));
  nand2 gate650(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate651(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate652(.a(G257), .O(gate238inter7));
  inv1  gate653(.a(G709), .O(gate238inter8));
  nand2 gate654(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate655(.a(s_15), .b(gate238inter3), .O(gate238inter10));
  nor2  gate656(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate657(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate658(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate869(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate870(.a(gate241inter0), .b(s_46), .O(gate241inter1));
  and2  gate871(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate872(.a(s_46), .O(gate241inter3));
  inv1  gate873(.a(s_47), .O(gate241inter4));
  nand2 gate874(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate875(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate876(.a(G242), .O(gate241inter7));
  inv1  gate877(.a(G730), .O(gate241inter8));
  nand2 gate878(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate879(.a(s_47), .b(gate241inter3), .O(gate241inter10));
  nor2  gate880(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate881(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate882(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate1667(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate1668(.a(gate245inter0), .b(s_160), .O(gate245inter1));
  and2  gate1669(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate1670(.a(s_160), .O(gate245inter3));
  inv1  gate1671(.a(s_161), .O(gate245inter4));
  nand2 gate1672(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate1673(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate1674(.a(G248), .O(gate245inter7));
  inv1  gate1675(.a(G736), .O(gate245inter8));
  nand2 gate1676(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate1677(.a(s_161), .b(gate245inter3), .O(gate245inter10));
  nor2  gate1678(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate1679(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate1680(.a(gate245inter12), .b(gate245inter1), .O(G758));
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );

  xor2  gate1191(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate1192(.a(gate259inter0), .b(s_92), .O(gate259inter1));
  and2  gate1193(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate1194(.a(s_92), .O(gate259inter3));
  inv1  gate1195(.a(s_93), .O(gate259inter4));
  nand2 gate1196(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate1197(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate1198(.a(G758), .O(gate259inter7));
  inv1  gate1199(.a(G759), .O(gate259inter8));
  nand2 gate1200(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate1201(.a(s_93), .b(gate259inter3), .O(gate259inter10));
  nor2  gate1202(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate1203(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate1204(.a(gate259inter12), .b(gate259inter1), .O(G776));

  xor2  gate1499(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate1500(.a(gate260inter0), .b(s_136), .O(gate260inter1));
  and2  gate1501(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate1502(.a(s_136), .O(gate260inter3));
  inv1  gate1503(.a(s_137), .O(gate260inter4));
  nand2 gate1504(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate1505(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate1506(.a(G760), .O(gate260inter7));
  inv1  gate1507(.a(G761), .O(gate260inter8));
  nand2 gate1508(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate1509(.a(s_137), .b(gate260inter3), .O(gate260inter10));
  nor2  gate1510(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate1511(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate1512(.a(gate260inter12), .b(gate260inter1), .O(G779));
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate2157(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate2158(.a(gate262inter0), .b(s_230), .O(gate262inter1));
  and2  gate2159(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate2160(.a(s_230), .O(gate262inter3));
  inv1  gate2161(.a(s_231), .O(gate262inter4));
  nand2 gate2162(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate2163(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate2164(.a(G764), .O(gate262inter7));
  inv1  gate2165(.a(G765), .O(gate262inter8));
  nand2 gate2166(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate2167(.a(s_231), .b(gate262inter3), .O(gate262inter10));
  nor2  gate2168(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate2169(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate2170(.a(gate262inter12), .b(gate262inter1), .O(G785));

  xor2  gate1149(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate1150(.a(gate263inter0), .b(s_86), .O(gate263inter1));
  and2  gate1151(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate1152(.a(s_86), .O(gate263inter3));
  inv1  gate1153(.a(s_87), .O(gate263inter4));
  nand2 gate1154(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate1155(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate1156(.a(G766), .O(gate263inter7));
  inv1  gate1157(.a(G767), .O(gate263inter8));
  nand2 gate1158(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate1159(.a(s_87), .b(gate263inter3), .O(gate263inter10));
  nor2  gate1160(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate1161(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate1162(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate855(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate856(.a(gate272inter0), .b(s_44), .O(gate272inter1));
  and2  gate857(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate858(.a(s_44), .O(gate272inter3));
  inv1  gate859(.a(s_45), .O(gate272inter4));
  nand2 gate860(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate861(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate862(.a(G663), .O(gate272inter7));
  inv1  gate863(.a(G791), .O(gate272inter8));
  nand2 gate864(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate865(.a(s_45), .b(gate272inter3), .O(gate272inter10));
  nor2  gate866(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate867(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate868(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );

  xor2  gate631(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate632(.a(gate276inter0), .b(s_12), .O(gate276inter1));
  and2  gate633(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate634(.a(s_12), .O(gate276inter3));
  inv1  gate635(.a(s_13), .O(gate276inter4));
  nand2 gate636(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate637(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate638(.a(G773), .O(gate276inter7));
  inv1  gate639(.a(G797), .O(gate276inter8));
  nand2 gate640(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate641(.a(s_13), .b(gate276inter3), .O(gate276inter10));
  nor2  gate642(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate643(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate644(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate1415(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate1416(.a(gate280inter0), .b(s_124), .O(gate280inter1));
  and2  gate1417(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate1418(.a(s_124), .O(gate280inter3));
  inv1  gate1419(.a(s_125), .O(gate280inter4));
  nand2 gate1420(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate1421(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate1422(.a(G779), .O(gate280inter7));
  inv1  gate1423(.a(G803), .O(gate280inter8));
  nand2 gate1424(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate1425(.a(s_125), .b(gate280inter3), .O(gate280inter10));
  nor2  gate1426(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate1427(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate1428(.a(gate280inter12), .b(gate280inter1), .O(G825));

  xor2  gate1009(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate1010(.a(gate281inter0), .b(s_66), .O(gate281inter1));
  and2  gate1011(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate1012(.a(s_66), .O(gate281inter3));
  inv1  gate1013(.a(s_67), .O(gate281inter4));
  nand2 gate1014(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate1015(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate1016(.a(G654), .O(gate281inter7));
  inv1  gate1017(.a(G806), .O(gate281inter8));
  nand2 gate1018(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate1019(.a(s_67), .b(gate281inter3), .O(gate281inter10));
  nor2  gate1020(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate1021(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate1022(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );

  xor2  gate2129(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate2130(.a(gate284inter0), .b(s_226), .O(gate284inter1));
  and2  gate2131(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate2132(.a(s_226), .O(gate284inter3));
  inv1  gate2133(.a(s_227), .O(gate284inter4));
  nand2 gate2134(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate2135(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate2136(.a(G785), .O(gate284inter7));
  inv1  gate2137(.a(G809), .O(gate284inter8));
  nand2 gate2138(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate2139(.a(s_227), .b(gate284inter3), .O(gate284inter10));
  nor2  gate2140(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate2141(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate2142(.a(gate284inter12), .b(gate284inter1), .O(G829));
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate1737(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate1738(.a(gate286inter0), .b(s_170), .O(gate286inter1));
  and2  gate1739(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate1740(.a(s_170), .O(gate286inter3));
  inv1  gate1741(.a(s_171), .O(gate286inter4));
  nand2 gate1742(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate1743(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate1744(.a(G788), .O(gate286inter7));
  inv1  gate1745(.a(G812), .O(gate286inter8));
  nand2 gate1746(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate1747(.a(s_171), .b(gate286inter3), .O(gate286inter10));
  nor2  gate1748(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate1749(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate1750(.a(gate286inter12), .b(gate286inter1), .O(G831));
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate2269(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate2270(.a(gate288inter0), .b(s_246), .O(gate288inter1));
  and2  gate2271(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate2272(.a(s_246), .O(gate288inter3));
  inv1  gate2273(.a(s_247), .O(gate288inter4));
  nand2 gate2274(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate2275(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate2276(.a(G791), .O(gate288inter7));
  inv1  gate2277(.a(G815), .O(gate288inter8));
  nand2 gate2278(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate2279(.a(s_247), .b(gate288inter3), .O(gate288inter10));
  nor2  gate2280(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate2281(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate2282(.a(gate288inter12), .b(gate288inter1), .O(G833));

  xor2  gate925(.a(G819), .b(G818), .O(gate289inter0));
  nand2 gate926(.a(gate289inter0), .b(s_54), .O(gate289inter1));
  and2  gate927(.a(G819), .b(G818), .O(gate289inter2));
  inv1  gate928(.a(s_54), .O(gate289inter3));
  inv1  gate929(.a(s_55), .O(gate289inter4));
  nand2 gate930(.a(gate289inter4), .b(gate289inter3), .O(gate289inter5));
  nor2  gate931(.a(gate289inter5), .b(gate289inter2), .O(gate289inter6));
  inv1  gate932(.a(G818), .O(gate289inter7));
  inv1  gate933(.a(G819), .O(gate289inter8));
  nand2 gate934(.a(gate289inter8), .b(gate289inter7), .O(gate289inter9));
  nand2 gate935(.a(s_55), .b(gate289inter3), .O(gate289inter10));
  nor2  gate936(.a(gate289inter10), .b(gate289inter9), .O(gate289inter11));
  nor2  gate937(.a(gate289inter11), .b(gate289inter6), .O(gate289inter12));
  nand2 gate938(.a(gate289inter12), .b(gate289inter1), .O(G834));
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate1877(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate1878(.a(gate292inter0), .b(s_190), .O(gate292inter1));
  and2  gate1879(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate1880(.a(s_190), .O(gate292inter3));
  inv1  gate1881(.a(s_191), .O(gate292inter4));
  nand2 gate1882(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate1883(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate1884(.a(G824), .O(gate292inter7));
  inv1  gate1885(.a(G825), .O(gate292inter8));
  nand2 gate1886(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate1887(.a(s_191), .b(gate292inter3), .O(gate292inter10));
  nor2  gate1888(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate1889(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate1890(.a(gate292inter12), .b(gate292inter1), .O(G873));

  xor2  gate1317(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate1318(.a(gate293inter0), .b(s_110), .O(gate293inter1));
  and2  gate1319(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate1320(.a(s_110), .O(gate293inter3));
  inv1  gate1321(.a(s_111), .O(gate293inter4));
  nand2 gate1322(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate1323(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate1324(.a(G828), .O(gate293inter7));
  inv1  gate1325(.a(G829), .O(gate293inter8));
  nand2 gate1326(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate1327(.a(s_111), .b(gate293inter3), .O(gate293inter10));
  nor2  gate1328(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate1329(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate1330(.a(gate293inter12), .b(gate293inter1), .O(G886));

  xor2  gate1429(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate1430(.a(gate294inter0), .b(s_126), .O(gate294inter1));
  and2  gate1431(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate1432(.a(s_126), .O(gate294inter3));
  inv1  gate1433(.a(s_127), .O(gate294inter4));
  nand2 gate1434(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate1435(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate1436(.a(G832), .O(gate294inter7));
  inv1  gate1437(.a(G833), .O(gate294inter8));
  nand2 gate1438(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate1439(.a(s_127), .b(gate294inter3), .O(gate294inter10));
  nor2  gate1440(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate1441(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate1442(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate2185(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate2186(.a(gate296inter0), .b(s_234), .O(gate296inter1));
  and2  gate2187(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate2188(.a(s_234), .O(gate296inter3));
  inv1  gate2189(.a(s_235), .O(gate296inter4));
  nand2 gate2190(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate2191(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate2192(.a(G826), .O(gate296inter7));
  inv1  gate2193(.a(G827), .O(gate296inter8));
  nand2 gate2194(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate2195(.a(s_235), .b(gate296inter3), .O(gate296inter10));
  nor2  gate2196(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate2197(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate2198(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate1835(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate1836(.a(gate389inter0), .b(s_184), .O(gate389inter1));
  and2  gate1837(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate1838(.a(s_184), .O(gate389inter3));
  inv1  gate1839(.a(s_185), .O(gate389inter4));
  nand2 gate1840(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate1841(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate1842(.a(G3), .O(gate389inter7));
  inv1  gate1843(.a(G1042), .O(gate389inter8));
  nand2 gate1844(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate1845(.a(s_185), .b(gate389inter3), .O(gate389inter10));
  nor2  gate1846(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate1847(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate1848(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );

  xor2  gate2059(.a(G1063), .b(G10), .O(gate396inter0));
  nand2 gate2060(.a(gate396inter0), .b(s_216), .O(gate396inter1));
  and2  gate2061(.a(G1063), .b(G10), .O(gate396inter2));
  inv1  gate2062(.a(s_216), .O(gate396inter3));
  inv1  gate2063(.a(s_217), .O(gate396inter4));
  nand2 gate2064(.a(gate396inter4), .b(gate396inter3), .O(gate396inter5));
  nor2  gate2065(.a(gate396inter5), .b(gate396inter2), .O(gate396inter6));
  inv1  gate2066(.a(G10), .O(gate396inter7));
  inv1  gate2067(.a(G1063), .O(gate396inter8));
  nand2 gate2068(.a(gate396inter8), .b(gate396inter7), .O(gate396inter9));
  nand2 gate2069(.a(s_217), .b(gate396inter3), .O(gate396inter10));
  nor2  gate2070(.a(gate396inter10), .b(gate396inter9), .O(gate396inter11));
  nor2  gate2071(.a(gate396inter11), .b(gate396inter6), .O(gate396inter12));
  nand2 gate2072(.a(gate396inter12), .b(gate396inter1), .O(G1159));
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate1709(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate1710(.a(gate399inter0), .b(s_166), .O(gate399inter1));
  and2  gate1711(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate1712(.a(s_166), .O(gate399inter3));
  inv1  gate1713(.a(s_167), .O(gate399inter4));
  nand2 gate1714(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate1715(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate1716(.a(G13), .O(gate399inter7));
  inv1  gate1717(.a(G1072), .O(gate399inter8));
  nand2 gate1718(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate1719(.a(s_167), .b(gate399inter3), .O(gate399inter10));
  nor2  gate1720(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate1721(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate1722(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );

  xor2  gate2045(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate2046(.a(gate401inter0), .b(s_214), .O(gate401inter1));
  and2  gate2047(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate2048(.a(s_214), .O(gate401inter3));
  inv1  gate2049(.a(s_215), .O(gate401inter4));
  nand2 gate2050(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate2051(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate2052(.a(G15), .O(gate401inter7));
  inv1  gate2053(.a(G1078), .O(gate401inter8));
  nand2 gate2054(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate2055(.a(s_215), .b(gate401inter3), .O(gate401inter10));
  nor2  gate2056(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate2057(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate2058(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate2017(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate2018(.a(gate403inter0), .b(s_210), .O(gate403inter1));
  and2  gate2019(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate2020(.a(s_210), .O(gate403inter3));
  inv1  gate2021(.a(s_211), .O(gate403inter4));
  nand2 gate2022(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate2023(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate2024(.a(G17), .O(gate403inter7));
  inv1  gate2025(.a(G1084), .O(gate403inter8));
  nand2 gate2026(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate2027(.a(s_211), .b(gate403inter3), .O(gate403inter10));
  nor2  gate2028(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate2029(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate2030(.a(gate403inter12), .b(gate403inter1), .O(G1180));
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );

  xor2  gate1933(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate1934(.a(gate405inter0), .b(s_198), .O(gate405inter1));
  and2  gate1935(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate1936(.a(s_198), .O(gate405inter3));
  inv1  gate1937(.a(s_199), .O(gate405inter4));
  nand2 gate1938(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate1939(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate1940(.a(G19), .O(gate405inter7));
  inv1  gate1941(.a(G1090), .O(gate405inter8));
  nand2 gate1942(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate1943(.a(s_199), .b(gate405inter3), .O(gate405inter10));
  nor2  gate1944(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate1945(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate1946(.a(gate405inter12), .b(gate405inter1), .O(G1186));
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );

  xor2  gate2213(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate2214(.a(gate416inter0), .b(s_238), .O(gate416inter1));
  and2  gate2215(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate2216(.a(s_238), .O(gate416inter3));
  inv1  gate2217(.a(s_239), .O(gate416inter4));
  nand2 gate2218(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate2219(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate2220(.a(G30), .O(gate416inter7));
  inv1  gate2221(.a(G1123), .O(gate416inter8));
  nand2 gate2222(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate2223(.a(s_239), .b(gate416inter3), .O(gate416inter10));
  nor2  gate2224(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate2225(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate2226(.a(gate416inter12), .b(gate416inter1), .O(G1219));
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );

  xor2  gate575(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate576(.a(gate424inter0), .b(s_4), .O(gate424inter1));
  and2  gate577(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate578(.a(s_4), .O(gate424inter3));
  inv1  gate579(.a(s_5), .O(gate424inter4));
  nand2 gate580(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate581(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate582(.a(G1042), .O(gate424inter7));
  inv1  gate583(.a(G1138), .O(gate424inter8));
  nand2 gate584(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate585(.a(s_5), .b(gate424inter3), .O(gate424inter10));
  nor2  gate586(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate587(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate588(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );

  xor2  gate1359(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate1360(.a(gate427inter0), .b(s_116), .O(gate427inter1));
  and2  gate1361(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate1362(.a(s_116), .O(gate427inter3));
  inv1  gate1363(.a(s_117), .O(gate427inter4));
  nand2 gate1364(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate1365(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate1366(.a(G5), .O(gate427inter7));
  inv1  gate1367(.a(G1144), .O(gate427inter8));
  nand2 gate1368(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate1369(.a(s_117), .b(gate427inter3), .O(gate427inter10));
  nor2  gate1370(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate1371(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate1372(.a(gate427inter12), .b(gate427inter1), .O(G1236));

  xor2  gate1373(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate1374(.a(gate428inter0), .b(s_118), .O(gate428inter1));
  and2  gate1375(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate1376(.a(s_118), .O(gate428inter3));
  inv1  gate1377(.a(s_119), .O(gate428inter4));
  nand2 gate1378(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate1379(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate1380(.a(G1048), .O(gate428inter7));
  inv1  gate1381(.a(G1144), .O(gate428inter8));
  nand2 gate1382(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate1383(.a(s_119), .b(gate428inter3), .O(gate428inter10));
  nor2  gate1384(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate1385(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate1386(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate1121(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate1122(.a(gate435inter0), .b(s_82), .O(gate435inter1));
  and2  gate1123(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate1124(.a(s_82), .O(gate435inter3));
  inv1  gate1125(.a(s_83), .O(gate435inter4));
  nand2 gate1126(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate1127(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate1128(.a(G9), .O(gate435inter7));
  inv1  gate1129(.a(G1156), .O(gate435inter8));
  nand2 gate1130(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate1131(.a(s_83), .b(gate435inter3), .O(gate435inter10));
  nor2  gate1132(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate1133(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate1134(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );

  xor2  gate1765(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate1766(.a(gate440inter0), .b(s_174), .O(gate440inter1));
  and2  gate1767(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate1768(.a(s_174), .O(gate440inter3));
  inv1  gate1769(.a(s_175), .O(gate440inter4));
  nand2 gate1770(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate1771(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate1772(.a(G1066), .O(gate440inter7));
  inv1  gate1773(.a(G1162), .O(gate440inter8));
  nand2 gate1774(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate1775(.a(s_175), .b(gate440inter3), .O(gate440inter10));
  nor2  gate1776(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate1777(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate1778(.a(gate440inter12), .b(gate440inter1), .O(G1249));
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate1989(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate1990(.a(gate442inter0), .b(s_206), .O(gate442inter1));
  and2  gate1991(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate1992(.a(s_206), .O(gate442inter3));
  inv1  gate1993(.a(s_207), .O(gate442inter4));
  nand2 gate1994(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate1995(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate1996(.a(G1069), .O(gate442inter7));
  inv1  gate1997(.a(G1165), .O(gate442inter8));
  nand2 gate1998(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate1999(.a(s_207), .b(gate442inter3), .O(gate442inter10));
  nor2  gate2000(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate2001(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate2002(.a(gate442inter12), .b(gate442inter1), .O(G1251));

  xor2  gate701(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate702(.a(gate443inter0), .b(s_22), .O(gate443inter1));
  and2  gate703(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate704(.a(s_22), .O(gate443inter3));
  inv1  gate705(.a(s_23), .O(gate443inter4));
  nand2 gate706(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate707(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate708(.a(G13), .O(gate443inter7));
  inv1  gate709(.a(G1168), .O(gate443inter8));
  nand2 gate710(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate711(.a(s_23), .b(gate443inter3), .O(gate443inter10));
  nor2  gate712(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate713(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate714(.a(gate443inter12), .b(gate443inter1), .O(G1252));

  xor2  gate1065(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate1066(.a(gate444inter0), .b(s_74), .O(gate444inter1));
  and2  gate1067(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate1068(.a(s_74), .O(gate444inter3));
  inv1  gate1069(.a(s_75), .O(gate444inter4));
  nand2 gate1070(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate1071(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate1072(.a(G1072), .O(gate444inter7));
  inv1  gate1073(.a(G1168), .O(gate444inter8));
  nand2 gate1074(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate1075(.a(s_75), .b(gate444inter3), .O(gate444inter10));
  nor2  gate1076(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate1077(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate1078(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );

  xor2  gate1849(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate1850(.a(gate449inter0), .b(s_186), .O(gate449inter1));
  and2  gate1851(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate1852(.a(s_186), .O(gate449inter3));
  inv1  gate1853(.a(s_187), .O(gate449inter4));
  nand2 gate1854(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate1855(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate1856(.a(G16), .O(gate449inter7));
  inv1  gate1857(.a(G1177), .O(gate449inter8));
  nand2 gate1858(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate1859(.a(s_187), .b(gate449inter3), .O(gate449inter10));
  nor2  gate1860(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate1861(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate1862(.a(gate449inter12), .b(gate449inter1), .O(G1258));

  xor2  gate1079(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate1080(.a(gate450inter0), .b(s_76), .O(gate450inter1));
  and2  gate1081(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate1082(.a(s_76), .O(gate450inter3));
  inv1  gate1083(.a(s_77), .O(gate450inter4));
  nand2 gate1084(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate1085(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate1086(.a(G1081), .O(gate450inter7));
  inv1  gate1087(.a(G1177), .O(gate450inter8));
  nand2 gate1088(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate1089(.a(s_77), .b(gate450inter3), .O(gate450inter10));
  nor2  gate1090(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate1091(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate1092(.a(gate450inter12), .b(gate450inter1), .O(G1259));

  xor2  gate1905(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate1906(.a(gate451inter0), .b(s_194), .O(gate451inter1));
  and2  gate1907(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate1908(.a(s_194), .O(gate451inter3));
  inv1  gate1909(.a(s_195), .O(gate451inter4));
  nand2 gate1910(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate1911(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate1912(.a(G17), .O(gate451inter7));
  inv1  gate1913(.a(G1180), .O(gate451inter8));
  nand2 gate1914(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate1915(.a(s_195), .b(gate451inter3), .O(gate451inter10));
  nor2  gate1916(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate1917(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate1918(.a(gate451inter12), .b(gate451inter1), .O(G1260));

  xor2  gate603(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate604(.a(gate452inter0), .b(s_8), .O(gate452inter1));
  and2  gate605(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate606(.a(s_8), .O(gate452inter3));
  inv1  gate607(.a(s_9), .O(gate452inter4));
  nand2 gate608(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate609(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate610(.a(G1084), .O(gate452inter7));
  inv1  gate611(.a(G1180), .O(gate452inter8));
  nand2 gate612(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate613(.a(s_9), .b(gate452inter3), .O(gate452inter10));
  nor2  gate614(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate615(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate616(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate1107(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate1108(.a(gate456inter0), .b(s_80), .O(gate456inter1));
  and2  gate1109(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate1110(.a(s_80), .O(gate456inter3));
  inv1  gate1111(.a(s_81), .O(gate456inter4));
  nand2 gate1112(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate1113(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate1114(.a(G1090), .O(gate456inter7));
  inv1  gate1115(.a(G1186), .O(gate456inter8));
  nand2 gate1116(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate1117(.a(s_81), .b(gate456inter3), .O(gate456inter10));
  nor2  gate1118(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate1119(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate1120(.a(gate456inter12), .b(gate456inter1), .O(G1265));

  xor2  gate1037(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate1038(.a(gate457inter0), .b(s_70), .O(gate457inter1));
  and2  gate1039(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate1040(.a(s_70), .O(gate457inter3));
  inv1  gate1041(.a(s_71), .O(gate457inter4));
  nand2 gate1042(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate1043(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate1044(.a(G20), .O(gate457inter7));
  inv1  gate1045(.a(G1189), .O(gate457inter8));
  nand2 gate1046(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate1047(.a(s_71), .b(gate457inter3), .O(gate457inter10));
  nor2  gate1048(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate1049(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate1050(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate1219(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate1220(.a(gate461inter0), .b(s_96), .O(gate461inter1));
  and2  gate1221(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate1222(.a(s_96), .O(gate461inter3));
  inv1  gate1223(.a(s_97), .O(gate461inter4));
  nand2 gate1224(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate1225(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate1226(.a(G22), .O(gate461inter7));
  inv1  gate1227(.a(G1195), .O(gate461inter8));
  nand2 gate1228(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate1229(.a(s_97), .b(gate461inter3), .O(gate461inter10));
  nor2  gate1230(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate1231(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate1232(.a(gate461inter12), .b(gate461inter1), .O(G1270));
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate841(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate842(.a(gate463inter0), .b(s_42), .O(gate463inter1));
  and2  gate843(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate844(.a(s_42), .O(gate463inter3));
  inv1  gate845(.a(s_43), .O(gate463inter4));
  nand2 gate846(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate847(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate848(.a(G23), .O(gate463inter7));
  inv1  gate849(.a(G1198), .O(gate463inter8));
  nand2 gate850(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate851(.a(s_43), .b(gate463inter3), .O(gate463inter10));
  nor2  gate852(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate853(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate854(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate2171(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate2172(.a(gate466inter0), .b(s_232), .O(gate466inter1));
  and2  gate2173(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate2174(.a(s_232), .O(gate466inter3));
  inv1  gate2175(.a(s_233), .O(gate466inter4));
  nand2 gate2176(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate2177(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate2178(.a(G1105), .O(gate466inter7));
  inv1  gate2179(.a(G1201), .O(gate466inter8));
  nand2 gate2180(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate2181(.a(s_233), .b(gate466inter3), .O(gate466inter10));
  nor2  gate2182(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate2183(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate2184(.a(gate466inter12), .b(gate466inter1), .O(G1275));

  xor2  gate2003(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate2004(.a(gate467inter0), .b(s_208), .O(gate467inter1));
  and2  gate2005(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate2006(.a(s_208), .O(gate467inter3));
  inv1  gate2007(.a(s_209), .O(gate467inter4));
  nand2 gate2008(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate2009(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate2010(.a(G25), .O(gate467inter7));
  inv1  gate2011(.a(G1204), .O(gate467inter8));
  nand2 gate2012(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate2013(.a(s_209), .b(gate467inter3), .O(gate467inter10));
  nor2  gate2014(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate2015(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate2016(.a(gate467inter12), .b(gate467inter1), .O(G1276));

  xor2  gate2255(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate2256(.a(gate468inter0), .b(s_244), .O(gate468inter1));
  and2  gate2257(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate2258(.a(s_244), .O(gate468inter3));
  inv1  gate2259(.a(s_245), .O(gate468inter4));
  nand2 gate2260(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate2261(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate2262(.a(G1108), .O(gate468inter7));
  inv1  gate2263(.a(G1204), .O(gate468inter8));
  nand2 gate2264(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate2265(.a(s_245), .b(gate468inter3), .O(gate468inter10));
  nor2  gate2266(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate2267(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate2268(.a(gate468inter12), .b(gate468inter1), .O(G1277));

  xor2  gate1597(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate1598(.a(gate469inter0), .b(s_150), .O(gate469inter1));
  and2  gate1599(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate1600(.a(s_150), .O(gate469inter3));
  inv1  gate1601(.a(s_151), .O(gate469inter4));
  nand2 gate1602(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate1603(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate1604(.a(G26), .O(gate469inter7));
  inv1  gate1605(.a(G1207), .O(gate469inter8));
  nand2 gate1606(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate1607(.a(s_151), .b(gate469inter3), .O(gate469inter10));
  nor2  gate1608(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate1609(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate1610(.a(gate469inter12), .b(gate469inter1), .O(G1278));

  xor2  gate1723(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate1724(.a(gate470inter0), .b(s_168), .O(gate470inter1));
  and2  gate1725(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate1726(.a(s_168), .O(gate470inter3));
  inv1  gate1727(.a(s_169), .O(gate470inter4));
  nand2 gate1728(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate1729(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate1730(.a(G1111), .O(gate470inter7));
  inv1  gate1731(.a(G1207), .O(gate470inter8));
  nand2 gate1732(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate1733(.a(s_169), .b(gate470inter3), .O(gate470inter10));
  nor2  gate1734(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate1735(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate1736(.a(gate470inter12), .b(gate470inter1), .O(G1279));

  xor2  gate2073(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate2074(.a(gate471inter0), .b(s_218), .O(gate471inter1));
  and2  gate2075(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate2076(.a(s_218), .O(gate471inter3));
  inv1  gate2077(.a(s_219), .O(gate471inter4));
  nand2 gate2078(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate2079(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate2080(.a(G27), .O(gate471inter7));
  inv1  gate2081(.a(G1210), .O(gate471inter8));
  nand2 gate2082(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate2083(.a(s_219), .b(gate471inter3), .O(gate471inter10));
  nor2  gate2084(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate2085(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate2086(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate547(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate548(.a(gate475inter0), .b(s_0), .O(gate475inter1));
  and2  gate549(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate550(.a(s_0), .O(gate475inter3));
  inv1  gate551(.a(s_1), .O(gate475inter4));
  nand2 gate552(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate553(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate554(.a(G29), .O(gate475inter7));
  inv1  gate555(.a(G1216), .O(gate475inter8));
  nand2 gate556(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate557(.a(s_1), .b(gate475inter3), .O(gate475inter10));
  nor2  gate558(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate559(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate560(.a(gate475inter12), .b(gate475inter1), .O(G1284));
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate2115(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate2116(.a(gate477inter0), .b(s_224), .O(gate477inter1));
  and2  gate2117(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate2118(.a(s_224), .O(gate477inter3));
  inv1  gate2119(.a(s_225), .O(gate477inter4));
  nand2 gate2120(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate2121(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate2122(.a(G30), .O(gate477inter7));
  inv1  gate2123(.a(G1219), .O(gate477inter8));
  nand2 gate2124(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate2125(.a(s_225), .b(gate477inter3), .O(gate477inter10));
  nor2  gate2126(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate2127(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate2128(.a(gate477inter12), .b(gate477inter1), .O(G1286));

  xor2  gate1457(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate1458(.a(gate478inter0), .b(s_130), .O(gate478inter1));
  and2  gate1459(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate1460(.a(s_130), .O(gate478inter3));
  inv1  gate1461(.a(s_131), .O(gate478inter4));
  nand2 gate1462(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate1463(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate1464(.a(G1123), .O(gate478inter7));
  inv1  gate1465(.a(G1219), .O(gate478inter8));
  nand2 gate1466(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate1467(.a(s_131), .b(gate478inter3), .O(gate478inter10));
  nor2  gate1468(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate1469(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate1470(.a(gate478inter12), .b(gate478inter1), .O(G1287));
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );

  xor2  gate757(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate758(.a(gate483inter0), .b(s_30), .O(gate483inter1));
  and2  gate759(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate760(.a(s_30), .O(gate483inter3));
  inv1  gate761(.a(s_31), .O(gate483inter4));
  nand2 gate762(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate763(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate764(.a(G1228), .O(gate483inter7));
  inv1  gate765(.a(G1229), .O(gate483inter8));
  nand2 gate766(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate767(.a(s_31), .b(gate483inter3), .O(gate483inter10));
  nor2  gate768(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate769(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate770(.a(gate483inter12), .b(gate483inter1), .O(G1292));

  xor2  gate939(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate940(.a(gate484inter0), .b(s_56), .O(gate484inter1));
  and2  gate941(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate942(.a(s_56), .O(gate484inter3));
  inv1  gate943(.a(s_57), .O(gate484inter4));
  nand2 gate944(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate945(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate946(.a(G1230), .O(gate484inter7));
  inv1  gate947(.a(G1231), .O(gate484inter8));
  nand2 gate948(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate949(.a(s_57), .b(gate484inter3), .O(gate484inter10));
  nor2  gate950(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate951(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate952(.a(gate484inter12), .b(gate484inter1), .O(G1293));
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );

  xor2  gate1261(.a(G1249), .b(G1248), .O(gate493inter0));
  nand2 gate1262(.a(gate493inter0), .b(s_102), .O(gate493inter1));
  and2  gate1263(.a(G1249), .b(G1248), .O(gate493inter2));
  inv1  gate1264(.a(s_102), .O(gate493inter3));
  inv1  gate1265(.a(s_103), .O(gate493inter4));
  nand2 gate1266(.a(gate493inter4), .b(gate493inter3), .O(gate493inter5));
  nor2  gate1267(.a(gate493inter5), .b(gate493inter2), .O(gate493inter6));
  inv1  gate1268(.a(G1248), .O(gate493inter7));
  inv1  gate1269(.a(G1249), .O(gate493inter8));
  nand2 gate1270(.a(gate493inter8), .b(gate493inter7), .O(gate493inter9));
  nand2 gate1271(.a(s_103), .b(gate493inter3), .O(gate493inter10));
  nor2  gate1272(.a(gate493inter10), .b(gate493inter9), .O(gate493inter11));
  nor2  gate1273(.a(gate493inter11), .b(gate493inter6), .O(gate493inter12));
  nand2 gate1274(.a(gate493inter12), .b(gate493inter1), .O(G1302));
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate981(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate982(.a(gate510inter0), .b(s_62), .O(gate510inter1));
  and2  gate983(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate984(.a(s_62), .O(gate510inter3));
  inv1  gate985(.a(s_63), .O(gate510inter4));
  nand2 gate986(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate987(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate988(.a(G1282), .O(gate510inter7));
  inv1  gate989(.a(G1283), .O(gate510inter8));
  nand2 gate990(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate991(.a(s_63), .b(gate510inter3), .O(gate510inter10));
  nor2  gate992(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate993(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate994(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );

  xor2  gate1975(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate1976(.a(gate512inter0), .b(s_204), .O(gate512inter1));
  and2  gate1977(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate1978(.a(s_204), .O(gate512inter3));
  inv1  gate1979(.a(s_205), .O(gate512inter4));
  nand2 gate1980(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate1981(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate1982(.a(G1286), .O(gate512inter7));
  inv1  gate1983(.a(G1287), .O(gate512inter8));
  nand2 gate1984(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate1985(.a(s_205), .b(gate512inter3), .O(gate512inter10));
  nor2  gate1986(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate1987(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate1988(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule