module c432 (N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
             N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
             N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
             N99,N102,N105,N108,N112,N115,N223,N329,N370,N421,
             N430,N431,N432);
input N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
      N99,N102,N105,N108,N112,N115;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51;
output N223,N329,N370,N421,N430,N431,N432;
wire N118,N119,N122,N123,N126,N127,N130,N131,N134,N135,
     N138,N139,N142,N143,N146,N147,N150,N151,N154,N157,
     N158,N159,N162,N165,N168,N171,N174,N177,N180,N183,
     N184,N185,N186,N187,N188,N189,N190,N191,N192,N193,
     N194,N195,N196,N197,N198,N199,N203,N213,N224,N227,
     N230,N233,N236,N239,N242,N243,N246,N247,N250,N251,
     N254,N255,N256,N257,N258,N259,N260,N263,N264,N267,
     N270,N273,N276,N279,N282,N285,N288,N289,N290,N291,
     N292,N293,N294,N295,N296,N300,N301,N302,N303,N304,
     N305,N306,N307,N308,N309,N319,N330,N331,N332,N333,
     N334,N335,N336,N337,N338,N339,N340,N341,N342,N343,
     N344,N345,N346,N347,N348,N349,N350,N351,N352,N353,
     N354,N355,N356,N357,N360,N371,N372,N373,N374,N375,
     N376,N377,N378,N379,N380,N381,N386,N393,N399,N404,
     N407,N411,N414,N415,N416,N417,N418,N419,N420,N422,
     N425,N428,N429, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate28inter0, gate28inter1, gate28inter2, gate28inter3, gate28inter4, gate28inter5, gate28inter6, gate28inter7, gate28inter8, gate28inter9, gate28inter10, gate28inter11, gate28inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate30inter0, gate30inter1, gate30inter2, gate30inter3, gate30inter4, gate30inter5, gate30inter6, gate30inter7, gate30inter8, gate30inter9, gate30inter10, gate30inter11, gate30inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12;


inv1 gate1( .a(N1), .O(N118) );
inv1 gate2( .a(N4), .O(N119) );
inv1 gate3( .a(N11), .O(N122) );
inv1 gate4( .a(N17), .O(N123) );
inv1 gate5( .a(N24), .O(N126) );
inv1 gate6( .a(N30), .O(N127) );
inv1 gate7( .a(N37), .O(N130) );
inv1 gate8( .a(N43), .O(N131) );
inv1 gate9( .a(N50), .O(N134) );
inv1 gate10( .a(N56), .O(N135) );
inv1 gate11( .a(N63), .O(N138) );
inv1 gate12( .a(N69), .O(N139) );
inv1 gate13( .a(N76), .O(N142) );
inv1 gate14( .a(N82), .O(N143) );
inv1 gate15( .a(N89), .O(N146) );
inv1 gate16( .a(N95), .O(N147) );
inv1 gate17( .a(N102), .O(N150) );
inv1 gate18( .a(N108), .O(N151) );

  xor2  gate357(.a(N4), .b(N118), .O(gate19inter0));
  nand2 gate358(.a(gate19inter0), .b(s_28), .O(gate19inter1));
  and2  gate359(.a(N4), .b(N118), .O(gate19inter2));
  inv1  gate360(.a(s_28), .O(gate19inter3));
  inv1  gate361(.a(s_29), .O(gate19inter4));
  nand2 gate362(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate363(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate364(.a(N118), .O(gate19inter7));
  inv1  gate365(.a(N4), .O(gate19inter8));
  nand2 gate366(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate367(.a(s_29), .b(gate19inter3), .O(gate19inter10));
  nor2  gate368(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate369(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate370(.a(gate19inter12), .b(gate19inter1), .O(N154));

  xor2  gate245(.a(N119), .b(N8), .O(gate20inter0));
  nand2 gate246(.a(gate20inter0), .b(s_12), .O(gate20inter1));
  and2  gate247(.a(N119), .b(N8), .O(gate20inter2));
  inv1  gate248(.a(s_12), .O(gate20inter3));
  inv1  gate249(.a(s_13), .O(gate20inter4));
  nand2 gate250(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate251(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate252(.a(N8), .O(gate20inter7));
  inv1  gate253(.a(N119), .O(gate20inter8));
  nand2 gate254(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate255(.a(s_13), .b(gate20inter3), .O(gate20inter10));
  nor2  gate256(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate257(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate258(.a(gate20inter12), .b(gate20inter1), .O(N157));
nor2 gate21( .a(N14), .b(N119), .O(N158) );
nand2 gate22( .a(N122), .b(N17), .O(N159) );
nand2 gate23( .a(N126), .b(N30), .O(N162) );
nand2 gate24( .a(N130), .b(N43), .O(N165) );
nand2 gate25( .a(N134), .b(N56), .O(N168) );

  xor2  gate441(.a(N69), .b(N138), .O(gate26inter0));
  nand2 gate442(.a(gate26inter0), .b(s_40), .O(gate26inter1));
  and2  gate443(.a(N69), .b(N138), .O(gate26inter2));
  inv1  gate444(.a(s_40), .O(gate26inter3));
  inv1  gate445(.a(s_41), .O(gate26inter4));
  nand2 gate446(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate447(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate448(.a(N138), .O(gate26inter7));
  inv1  gate449(.a(N69), .O(gate26inter8));
  nand2 gate450(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate451(.a(s_41), .b(gate26inter3), .O(gate26inter10));
  nor2  gate452(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate453(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate454(.a(gate26inter12), .b(gate26inter1), .O(N171));
nand2 gate27( .a(N142), .b(N82), .O(N174) );

  xor2  gate203(.a(N95), .b(N146), .O(gate28inter0));
  nand2 gate204(.a(gate28inter0), .b(s_6), .O(gate28inter1));
  and2  gate205(.a(N95), .b(N146), .O(gate28inter2));
  inv1  gate206(.a(s_6), .O(gate28inter3));
  inv1  gate207(.a(s_7), .O(gate28inter4));
  nand2 gate208(.a(gate28inter4), .b(gate28inter3), .O(gate28inter5));
  nor2  gate209(.a(gate28inter5), .b(gate28inter2), .O(gate28inter6));
  inv1  gate210(.a(N146), .O(gate28inter7));
  inv1  gate211(.a(N95), .O(gate28inter8));
  nand2 gate212(.a(gate28inter8), .b(gate28inter7), .O(gate28inter9));
  nand2 gate213(.a(s_7), .b(gate28inter3), .O(gate28inter10));
  nor2  gate214(.a(gate28inter10), .b(gate28inter9), .O(gate28inter11));
  nor2  gate215(.a(gate28inter11), .b(gate28inter6), .O(gate28inter12));
  nand2 gate216(.a(gate28inter12), .b(gate28inter1), .O(N177));
nand2 gate29( .a(N150), .b(N108), .O(N180) );

  xor2  gate343(.a(N123), .b(N21), .O(gate30inter0));
  nand2 gate344(.a(gate30inter0), .b(s_26), .O(gate30inter1));
  and2  gate345(.a(N123), .b(N21), .O(gate30inter2));
  inv1  gate346(.a(s_26), .O(gate30inter3));
  inv1  gate347(.a(s_27), .O(gate30inter4));
  nand2 gate348(.a(gate30inter4), .b(gate30inter3), .O(gate30inter5));
  nor2  gate349(.a(gate30inter5), .b(gate30inter2), .O(gate30inter6));
  inv1  gate350(.a(N21), .O(gate30inter7));
  inv1  gate351(.a(N123), .O(gate30inter8));
  nand2 gate352(.a(gate30inter8), .b(gate30inter7), .O(gate30inter9));
  nand2 gate353(.a(s_27), .b(gate30inter3), .O(gate30inter10));
  nor2  gate354(.a(gate30inter10), .b(gate30inter9), .O(gate30inter11));
  nor2  gate355(.a(gate30inter11), .b(gate30inter6), .O(gate30inter12));
  nand2 gate356(.a(gate30inter12), .b(gate30inter1), .O(N183));

  xor2  gate259(.a(N123), .b(N27), .O(gate31inter0));
  nand2 gate260(.a(gate31inter0), .b(s_14), .O(gate31inter1));
  and2  gate261(.a(N123), .b(N27), .O(gate31inter2));
  inv1  gate262(.a(s_14), .O(gate31inter3));
  inv1  gate263(.a(s_15), .O(gate31inter4));
  nand2 gate264(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate265(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate266(.a(N27), .O(gate31inter7));
  inv1  gate267(.a(N123), .O(gate31inter8));
  nand2 gate268(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate269(.a(s_15), .b(gate31inter3), .O(gate31inter10));
  nor2  gate270(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate271(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate272(.a(gate31inter12), .b(gate31inter1), .O(N184));
nor2 gate32( .a(N34), .b(N127), .O(N185) );
nor2 gate33( .a(N40), .b(N127), .O(N186) );
nor2 gate34( .a(N47), .b(N131), .O(N187) );
nor2 gate35( .a(N53), .b(N131), .O(N188) );
nor2 gate36( .a(N60), .b(N135), .O(N189) );
nor2 gate37( .a(N66), .b(N135), .O(N190) );
nor2 gate38( .a(N73), .b(N139), .O(N191) );
nor2 gate39( .a(N79), .b(N139), .O(N192) );
nor2 gate40( .a(N86), .b(N143), .O(N193) );
nor2 gate41( .a(N92), .b(N143), .O(N194) );
nor2 gate42( .a(N99), .b(N147), .O(N195) );

  xor2  gate497(.a(N147), .b(N105), .O(gate43inter0));
  nand2 gate498(.a(gate43inter0), .b(s_48), .O(gate43inter1));
  and2  gate499(.a(N147), .b(N105), .O(gate43inter2));
  inv1  gate500(.a(s_48), .O(gate43inter3));
  inv1  gate501(.a(s_49), .O(gate43inter4));
  nand2 gate502(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate503(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate504(.a(N105), .O(gate43inter7));
  inv1  gate505(.a(N147), .O(gate43inter8));
  nand2 gate506(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate507(.a(s_49), .b(gate43inter3), .O(gate43inter10));
  nor2  gate508(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate509(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate510(.a(gate43inter12), .b(gate43inter1), .O(N196));
nor2 gate44( .a(N112), .b(N151), .O(N197) );
nor2 gate45( .a(N115), .b(N151), .O(N198) );
and9 gate46( .a(N154), .b(N159), .c(N162), .d(N165), .e(N168), .f(N171), .g(N174), .h(N177), .i(N180), .O(N199) );
inv1 gate47( .a(N199), .O(N203) );
inv1 gate48( .a(N199), .O(N213) );
inv1 gate49( .a(N199), .O(N223) );

  xor2  gate511(.a(N154), .b(N203), .O(gate50inter0));
  nand2 gate512(.a(gate50inter0), .b(s_50), .O(gate50inter1));
  and2  gate513(.a(N154), .b(N203), .O(gate50inter2));
  inv1  gate514(.a(s_50), .O(gate50inter3));
  inv1  gate515(.a(s_51), .O(gate50inter4));
  nand2 gate516(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate517(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate518(.a(N203), .O(gate50inter7));
  inv1  gate519(.a(N154), .O(gate50inter8));
  nand2 gate520(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate521(.a(s_51), .b(gate50inter3), .O(gate50inter10));
  nor2  gate522(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate523(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate524(.a(gate50inter12), .b(gate50inter1), .O(N224));

  xor2  gate175(.a(N159), .b(N203), .O(gate51inter0));
  nand2 gate176(.a(gate51inter0), .b(s_2), .O(gate51inter1));
  and2  gate177(.a(N159), .b(N203), .O(gate51inter2));
  inv1  gate178(.a(s_2), .O(gate51inter3));
  inv1  gate179(.a(s_3), .O(gate51inter4));
  nand2 gate180(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate181(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate182(.a(N203), .O(gate51inter7));
  inv1  gate183(.a(N159), .O(gate51inter8));
  nand2 gate184(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate185(.a(s_3), .b(gate51inter3), .O(gate51inter10));
  nor2  gate186(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate187(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate188(.a(gate51inter12), .b(gate51inter1), .O(N227));
xor2 gate52( .a(N203), .b(N162), .O(N230) );
xor2 gate53( .a(N203), .b(N165), .O(N233) );
xor2 gate54( .a(N203), .b(N168), .O(N236) );
xor2 gate55( .a(N203), .b(N171), .O(N239) );

  xor2  gate469(.a(N213), .b(N1), .O(gate56inter0));
  nand2 gate470(.a(gate56inter0), .b(s_44), .O(gate56inter1));
  and2  gate471(.a(N213), .b(N1), .O(gate56inter2));
  inv1  gate472(.a(s_44), .O(gate56inter3));
  inv1  gate473(.a(s_45), .O(gate56inter4));
  nand2 gate474(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate475(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate476(.a(N1), .O(gate56inter7));
  inv1  gate477(.a(N213), .O(gate56inter8));
  nand2 gate478(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate479(.a(s_45), .b(gate56inter3), .O(gate56inter10));
  nor2  gate480(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate481(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate482(.a(gate56inter12), .b(gate56inter1), .O(N242));
xor2 gate57( .a(N203), .b(N174), .O(N243) );

  xor2  gate399(.a(N11), .b(N213), .O(gate58inter0));
  nand2 gate400(.a(gate58inter0), .b(s_34), .O(gate58inter1));
  and2  gate401(.a(N11), .b(N213), .O(gate58inter2));
  inv1  gate402(.a(s_34), .O(gate58inter3));
  inv1  gate403(.a(s_35), .O(gate58inter4));
  nand2 gate404(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate405(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate406(.a(N213), .O(gate58inter7));
  inv1  gate407(.a(N11), .O(gate58inter8));
  nand2 gate408(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate409(.a(s_35), .b(gate58inter3), .O(gate58inter10));
  nor2  gate410(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate411(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate412(.a(gate58inter12), .b(gate58inter1), .O(N246));

  xor2  gate455(.a(N177), .b(N203), .O(gate59inter0));
  nand2 gate456(.a(gate59inter0), .b(s_42), .O(gate59inter1));
  and2  gate457(.a(N177), .b(N203), .O(gate59inter2));
  inv1  gate458(.a(s_42), .O(gate59inter3));
  inv1  gate459(.a(s_43), .O(gate59inter4));
  nand2 gate460(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate461(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate462(.a(N203), .O(gate59inter7));
  inv1  gate463(.a(N177), .O(gate59inter8));
  nand2 gate464(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate465(.a(s_43), .b(gate59inter3), .O(gate59inter10));
  nor2  gate466(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate467(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate468(.a(gate59inter12), .b(gate59inter1), .O(N247));
nand2 gate60( .a(N213), .b(N24), .O(N250) );
xor2 gate61( .a(N203), .b(N180), .O(N251) );
nand2 gate62( .a(N213), .b(N37), .O(N254) );
nand2 gate63( .a(N213), .b(N50), .O(N255) );
nand2 gate64( .a(N213), .b(N63), .O(N256) );
nand2 gate65( .a(N213), .b(N76), .O(N257) );

  xor2  gate371(.a(N89), .b(N213), .O(gate66inter0));
  nand2 gate372(.a(gate66inter0), .b(s_30), .O(gate66inter1));
  and2  gate373(.a(N89), .b(N213), .O(gate66inter2));
  inv1  gate374(.a(s_30), .O(gate66inter3));
  inv1  gate375(.a(s_31), .O(gate66inter4));
  nand2 gate376(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate377(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate378(.a(N213), .O(gate66inter7));
  inv1  gate379(.a(N89), .O(gate66inter8));
  nand2 gate380(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate381(.a(s_31), .b(gate66inter3), .O(gate66inter10));
  nor2  gate382(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate383(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate384(.a(gate66inter12), .b(gate66inter1), .O(N258));
nand2 gate67( .a(N213), .b(N102), .O(N259) );
nand2 gate68( .a(N224), .b(N157), .O(N260) );
nand2 gate69( .a(N224), .b(N158), .O(N263) );
nand2 gate70( .a(N227), .b(N183), .O(N264) );

  xor2  gate315(.a(N185), .b(N230), .O(gate71inter0));
  nand2 gate316(.a(gate71inter0), .b(s_22), .O(gate71inter1));
  and2  gate317(.a(N185), .b(N230), .O(gate71inter2));
  inv1  gate318(.a(s_22), .O(gate71inter3));
  inv1  gate319(.a(s_23), .O(gate71inter4));
  nand2 gate320(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate321(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate322(.a(N230), .O(gate71inter7));
  inv1  gate323(.a(N185), .O(gate71inter8));
  nand2 gate324(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate325(.a(s_23), .b(gate71inter3), .O(gate71inter10));
  nor2  gate326(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate327(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate328(.a(gate71inter12), .b(gate71inter1), .O(N267));
nand2 gate72( .a(N233), .b(N187), .O(N270) );

  xor2  gate385(.a(N189), .b(N236), .O(gate73inter0));
  nand2 gate386(.a(gate73inter0), .b(s_32), .O(gate73inter1));
  and2  gate387(.a(N189), .b(N236), .O(gate73inter2));
  inv1  gate388(.a(s_32), .O(gate73inter3));
  inv1  gate389(.a(s_33), .O(gate73inter4));
  nand2 gate390(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate391(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate392(.a(N236), .O(gate73inter7));
  inv1  gate393(.a(N189), .O(gate73inter8));
  nand2 gate394(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate395(.a(s_33), .b(gate73inter3), .O(gate73inter10));
  nor2  gate396(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate397(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate398(.a(gate73inter12), .b(gate73inter1), .O(N273));
nand2 gate74( .a(N239), .b(N191), .O(N276) );
nand2 gate75( .a(N243), .b(N193), .O(N279) );
nand2 gate76( .a(N247), .b(N195), .O(N282) );
nand2 gate77( .a(N251), .b(N197), .O(N285) );

  xor2  gate329(.a(N184), .b(N227), .O(gate78inter0));
  nand2 gate330(.a(gate78inter0), .b(s_24), .O(gate78inter1));
  and2  gate331(.a(N184), .b(N227), .O(gate78inter2));
  inv1  gate332(.a(s_24), .O(gate78inter3));
  inv1  gate333(.a(s_25), .O(gate78inter4));
  nand2 gate334(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate335(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate336(.a(N227), .O(gate78inter7));
  inv1  gate337(.a(N184), .O(gate78inter8));
  nand2 gate338(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate339(.a(s_25), .b(gate78inter3), .O(gate78inter10));
  nor2  gate340(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate341(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate342(.a(gate78inter12), .b(gate78inter1), .O(N288));
nand2 gate79( .a(N230), .b(N186), .O(N289) );
nand2 gate80( .a(N233), .b(N188), .O(N290) );
nand2 gate81( .a(N236), .b(N190), .O(N291) );
nand2 gate82( .a(N239), .b(N192), .O(N292) );
nand2 gate83( .a(N243), .b(N194), .O(N293) );

  xor2  gate217(.a(N196), .b(N247), .O(gate84inter0));
  nand2 gate218(.a(gate84inter0), .b(s_8), .O(gate84inter1));
  and2  gate219(.a(N196), .b(N247), .O(gate84inter2));
  inv1  gate220(.a(s_8), .O(gate84inter3));
  inv1  gate221(.a(s_9), .O(gate84inter4));
  nand2 gate222(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate223(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate224(.a(N247), .O(gate84inter7));
  inv1  gate225(.a(N196), .O(gate84inter8));
  nand2 gate226(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate227(.a(s_9), .b(gate84inter3), .O(gate84inter10));
  nor2  gate228(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate229(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate230(.a(gate84inter12), .b(gate84inter1), .O(N294));
nand2 gate85( .a(N251), .b(N198), .O(N295) );
and9 gate86( .a(N260), .b(N264), .c(N267), .d(N270), .e(N273), .f(N276), .g(N279), .h(N282), .i(N285), .O(N296) );
inv1 gate87( .a(N263), .O(N300) );
inv1 gate88( .a(N288), .O(N301) );
inv1 gate89( .a(N289), .O(N302) );
inv1 gate90( .a(N290), .O(N303) );
inv1 gate91( .a(N291), .O(N304) );
inv1 gate92( .a(N292), .O(N305) );
inv1 gate93( .a(N293), .O(N306) );
inv1 gate94( .a(N294), .O(N307) );
inv1 gate95( .a(N295), .O(N308) );
inv1 gate96( .a(N296), .O(N309) );
inv1 gate97( .a(N296), .O(N319) );
inv1 gate98( .a(N296), .O(N329) );
xor2 gate99( .a(N309), .b(N260), .O(N330) );
xor2 gate100( .a(N309), .b(N264), .O(N331) );
xor2 gate101( .a(N309), .b(N267), .O(N332) );
xor2 gate102( .a(N309), .b(N270), .O(N333) );
nand2 gate103( .a(N8), .b(N319), .O(N334) );
xor2 gate104( .a(N309), .b(N273), .O(N335) );
nand2 gate105( .a(N319), .b(N21), .O(N336) );
xor2 gate106( .a(N309), .b(N276), .O(N337) );
nand2 gate107( .a(N319), .b(N34), .O(N338) );
xor2 gate108( .a(N309), .b(N279), .O(N339) );
nand2 gate109( .a(N319), .b(N47), .O(N340) );
xor2 gate110( .a(N309), .b(N282), .O(N341) );

  xor2  gate427(.a(N60), .b(N319), .O(gate111inter0));
  nand2 gate428(.a(gate111inter0), .b(s_38), .O(gate111inter1));
  and2  gate429(.a(N60), .b(N319), .O(gate111inter2));
  inv1  gate430(.a(s_38), .O(gate111inter3));
  inv1  gate431(.a(s_39), .O(gate111inter4));
  nand2 gate432(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate433(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate434(.a(N319), .O(gate111inter7));
  inv1  gate435(.a(N60), .O(gate111inter8));
  nand2 gate436(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate437(.a(s_39), .b(gate111inter3), .O(gate111inter10));
  nor2  gate438(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate439(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate440(.a(gate111inter12), .b(gate111inter1), .O(N342));
xor2 gate112( .a(N309), .b(N285), .O(N343) );

  xor2  gate189(.a(N73), .b(N319), .O(gate113inter0));
  nand2 gate190(.a(gate113inter0), .b(s_4), .O(gate113inter1));
  and2  gate191(.a(N73), .b(N319), .O(gate113inter2));
  inv1  gate192(.a(s_4), .O(gate113inter3));
  inv1  gate193(.a(s_5), .O(gate113inter4));
  nand2 gate194(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate195(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate196(.a(N319), .O(gate113inter7));
  inv1  gate197(.a(N73), .O(gate113inter8));
  nand2 gate198(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate199(.a(s_5), .b(gate113inter3), .O(gate113inter10));
  nor2  gate200(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate201(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate202(.a(gate113inter12), .b(gate113inter1), .O(N344));
nand2 gate114( .a(N319), .b(N86), .O(N345) );
nand2 gate115( .a(N319), .b(N99), .O(N346) );
nand2 gate116( .a(N319), .b(N112), .O(N347) );
nand2 gate117( .a(N330), .b(N300), .O(N348) );
nand2 gate118( .a(N331), .b(N301), .O(N349) );

  xor2  gate483(.a(N302), .b(N332), .O(gate119inter0));
  nand2 gate484(.a(gate119inter0), .b(s_46), .O(gate119inter1));
  and2  gate485(.a(N302), .b(N332), .O(gate119inter2));
  inv1  gate486(.a(s_46), .O(gate119inter3));
  inv1  gate487(.a(s_47), .O(gate119inter4));
  nand2 gate488(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate489(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate490(.a(N332), .O(gate119inter7));
  inv1  gate491(.a(N302), .O(gate119inter8));
  nand2 gate492(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate493(.a(s_47), .b(gate119inter3), .O(gate119inter10));
  nor2  gate494(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate495(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate496(.a(gate119inter12), .b(gate119inter1), .O(N350));

  xor2  gate161(.a(N303), .b(N333), .O(gate120inter0));
  nand2 gate162(.a(gate120inter0), .b(s_0), .O(gate120inter1));
  and2  gate163(.a(N303), .b(N333), .O(gate120inter2));
  inv1  gate164(.a(s_0), .O(gate120inter3));
  inv1  gate165(.a(s_1), .O(gate120inter4));
  nand2 gate166(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate167(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate168(.a(N333), .O(gate120inter7));
  inv1  gate169(.a(N303), .O(gate120inter8));
  nand2 gate170(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate171(.a(s_1), .b(gate120inter3), .O(gate120inter10));
  nor2  gate172(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate173(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate174(.a(gate120inter12), .b(gate120inter1), .O(N351));
nand2 gate121( .a(N335), .b(N304), .O(N352) );
nand2 gate122( .a(N337), .b(N305), .O(N353) );
nand2 gate123( .a(N339), .b(N306), .O(N354) );
nand2 gate124( .a(N341), .b(N307), .O(N355) );

  xor2  gate231(.a(N308), .b(N343), .O(gate125inter0));
  nand2 gate232(.a(gate125inter0), .b(s_10), .O(gate125inter1));
  and2  gate233(.a(N308), .b(N343), .O(gate125inter2));
  inv1  gate234(.a(s_10), .O(gate125inter3));
  inv1  gate235(.a(s_11), .O(gate125inter4));
  nand2 gate236(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate237(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate238(.a(N343), .O(gate125inter7));
  inv1  gate239(.a(N308), .O(gate125inter8));
  nand2 gate240(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate241(.a(s_11), .b(gate125inter3), .O(gate125inter10));
  nor2  gate242(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate243(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate244(.a(gate125inter12), .b(gate125inter1), .O(N356));
and9 gate126( .a(N348), .b(N349), .c(N350), .d(N351), .e(N352), .f(N353), .g(N354), .h(N355), .i(N356), .O(N357) );
inv1 gate127( .a(N357), .O(N360) );
inv1 gate128( .a(N357), .O(N370) );
nand2 gate129( .a(N14), .b(N360), .O(N371) );
nand2 gate130( .a(N360), .b(N27), .O(N372) );

  xor2  gate273(.a(N40), .b(N360), .O(gate131inter0));
  nand2 gate274(.a(gate131inter0), .b(s_16), .O(gate131inter1));
  and2  gate275(.a(N40), .b(N360), .O(gate131inter2));
  inv1  gate276(.a(s_16), .O(gate131inter3));
  inv1  gate277(.a(s_17), .O(gate131inter4));
  nand2 gate278(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate279(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate280(.a(N360), .O(gate131inter7));
  inv1  gate281(.a(N40), .O(gate131inter8));
  nand2 gate282(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate283(.a(s_17), .b(gate131inter3), .O(gate131inter10));
  nor2  gate284(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate285(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate286(.a(gate131inter12), .b(gate131inter1), .O(N373));

  xor2  gate301(.a(N53), .b(N360), .O(gate132inter0));
  nand2 gate302(.a(gate132inter0), .b(s_20), .O(gate132inter1));
  and2  gate303(.a(N53), .b(N360), .O(gate132inter2));
  inv1  gate304(.a(s_20), .O(gate132inter3));
  inv1  gate305(.a(s_21), .O(gate132inter4));
  nand2 gate306(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate307(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate308(.a(N360), .O(gate132inter7));
  inv1  gate309(.a(N53), .O(gate132inter8));
  nand2 gate310(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate311(.a(s_21), .b(gate132inter3), .O(gate132inter10));
  nor2  gate312(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate313(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate314(.a(gate132inter12), .b(gate132inter1), .O(N374));
nand2 gate133( .a(N360), .b(N66), .O(N375) );
nand2 gate134( .a(N360), .b(N79), .O(N376) );

  xor2  gate413(.a(N92), .b(N360), .O(gate135inter0));
  nand2 gate414(.a(gate135inter0), .b(s_36), .O(gate135inter1));
  and2  gate415(.a(N92), .b(N360), .O(gate135inter2));
  inv1  gate416(.a(s_36), .O(gate135inter3));
  inv1  gate417(.a(s_37), .O(gate135inter4));
  nand2 gate418(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate419(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate420(.a(N360), .O(gate135inter7));
  inv1  gate421(.a(N92), .O(gate135inter8));
  nand2 gate422(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate423(.a(s_37), .b(gate135inter3), .O(gate135inter10));
  nor2  gate424(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate425(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate426(.a(gate135inter12), .b(gate135inter1), .O(N377));
nand2 gate136( .a(N360), .b(N105), .O(N378) );
nand2 gate137( .a(N360), .b(N115), .O(N379) );
nand4 gate138( .a(N4), .b(N242), .c(N334), .d(N371), .O(N380) );
nand4 gate139( .a(N246), .b(N336), .c(N372), .d(N17), .O(N381) );
nand4 gate140( .a(N250), .b(N338), .c(N373), .d(N30), .O(N386) );
nand4 gate141( .a(N254), .b(N340), .c(N374), .d(N43), .O(N393) );
nand4 gate142( .a(N255), .b(N342), .c(N375), .d(N56), .O(N399) );
nand4 gate143( .a(N256), .b(N344), .c(N376), .d(N69), .O(N404) );
nand4 gate144( .a(N257), .b(N345), .c(N377), .d(N82), .O(N407) );
nand4 gate145( .a(N258), .b(N346), .c(N378), .d(N95), .O(N411) );
nand4 gate146( .a(N259), .b(N347), .c(N379), .d(N108), .O(N414) );
inv1 gate147( .a(N380), .O(N415) );
and8 gate148( .a(N381), .b(N386), .c(N393), .d(N399), .e(N404), .f(N407), .g(N411), .h(N414), .O(N416) );
inv1 gate149( .a(N393), .O(N417) );
inv1 gate150( .a(N404), .O(N418) );
inv1 gate151( .a(N407), .O(N419) );
inv1 gate152( .a(N411), .O(N420) );
nor2 gate153( .a(N415), .b(N416), .O(N421) );

  xor2  gate287(.a(N417), .b(N386), .O(gate154inter0));
  nand2 gate288(.a(gate154inter0), .b(s_18), .O(gate154inter1));
  and2  gate289(.a(N417), .b(N386), .O(gate154inter2));
  inv1  gate290(.a(s_18), .O(gate154inter3));
  inv1  gate291(.a(s_19), .O(gate154inter4));
  nand2 gate292(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate293(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate294(.a(N386), .O(gate154inter7));
  inv1  gate295(.a(N417), .O(gate154inter8));
  nand2 gate296(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate297(.a(s_19), .b(gate154inter3), .O(gate154inter10));
  nor2  gate298(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate299(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate300(.a(gate154inter12), .b(gate154inter1), .O(N422));
nand4 gate155( .a(N386), .b(N393), .c(N418), .d(N399), .O(N425) );
nand3 gate156( .a(N399), .b(N393), .c(N419), .O(N428) );
nand4 gate157( .a(N386), .b(N393), .c(N407), .d(N420), .O(N429) );
nand4 gate158( .a(N381), .b(N386), .c(N422), .d(N399), .O(N430) );
nand4 gate159( .a(N381), .b(N386), .c(N425), .d(N428), .O(N431) );
nand4 gate160( .a(N381), .b(N422), .c(N425), .d(N429), .O(N432) );

endmodule