module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate259inter0, gate259inter1, gate259inter2, gate259inter3, gate259inter4, gate259inter5, gate259inter6, gate259inter7, gate259inter8, gate259inter9, gate259inter10, gate259inter11, gate259inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate1079(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate1080(.a(gate17inter0), .b(s_76), .O(gate17inter1));
  and2  gate1081(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate1082(.a(s_76), .O(gate17inter3));
  inv1  gate1083(.a(s_77), .O(gate17inter4));
  nand2 gate1084(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate1085(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate1086(.a(G17), .O(gate17inter7));
  inv1  gate1087(.a(G18), .O(gate17inter8));
  nand2 gate1088(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate1089(.a(s_77), .b(gate17inter3), .O(gate17inter10));
  nor2  gate1090(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate1091(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate1092(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );

  xor2  gate1233(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate1234(.a(gate32inter0), .b(s_98), .O(gate32inter1));
  and2  gate1235(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate1236(.a(s_98), .O(gate32inter3));
  inv1  gate1237(.a(s_99), .O(gate32inter4));
  nand2 gate1238(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate1239(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate1240(.a(G12), .O(gate32inter7));
  inv1  gate1241(.a(G16), .O(gate32inter8));
  nand2 gate1242(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate1243(.a(s_99), .b(gate32inter3), .O(gate32inter10));
  nor2  gate1244(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate1245(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate1246(.a(gate32inter12), .b(gate32inter1), .O(G335));
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );

  xor2  gate1135(.a(G22), .b(G18), .O(gate35inter0));
  nand2 gate1136(.a(gate35inter0), .b(s_84), .O(gate35inter1));
  and2  gate1137(.a(G22), .b(G18), .O(gate35inter2));
  inv1  gate1138(.a(s_84), .O(gate35inter3));
  inv1  gate1139(.a(s_85), .O(gate35inter4));
  nand2 gate1140(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate1141(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate1142(.a(G18), .O(gate35inter7));
  inv1  gate1143(.a(G22), .O(gate35inter8));
  nand2 gate1144(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate1145(.a(s_85), .b(gate35inter3), .O(gate35inter10));
  nor2  gate1146(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate1147(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate1148(.a(gate35inter12), .b(gate35inter1), .O(G344));
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );

  xor2  gate1317(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate1318(.a(gate40inter0), .b(s_110), .O(gate40inter1));
  and2  gate1319(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate1320(.a(s_110), .O(gate40inter3));
  inv1  gate1321(.a(s_111), .O(gate40inter4));
  nand2 gate1322(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate1323(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate1324(.a(G28), .O(gate40inter7));
  inv1  gate1325(.a(G32), .O(gate40inter8));
  nand2 gate1326(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate1327(.a(s_111), .b(gate40inter3), .O(gate40inter10));
  nor2  gate1328(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate1329(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate1330(.a(gate40inter12), .b(gate40inter1), .O(G359));
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );

  xor2  gate729(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate730(.a(gate47inter0), .b(s_26), .O(gate47inter1));
  and2  gate731(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate732(.a(s_26), .O(gate47inter3));
  inv1  gate733(.a(s_27), .O(gate47inter4));
  nand2 gate734(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate735(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate736(.a(G7), .O(gate47inter7));
  inv1  gate737(.a(G275), .O(gate47inter8));
  nand2 gate738(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate739(.a(s_27), .b(gate47inter3), .O(gate47inter10));
  nor2  gate740(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate741(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate742(.a(gate47inter12), .b(gate47inter1), .O(G368));
nand2 gate48( .a(G8), .b(G275), .O(G369) );

  xor2  gate1177(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate1178(.a(gate49inter0), .b(s_90), .O(gate49inter1));
  and2  gate1179(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate1180(.a(s_90), .O(gate49inter3));
  inv1  gate1181(.a(s_91), .O(gate49inter4));
  nand2 gate1182(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate1183(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate1184(.a(G9), .O(gate49inter7));
  inv1  gate1185(.a(G278), .O(gate49inter8));
  nand2 gate1186(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate1187(.a(s_91), .b(gate49inter3), .O(gate49inter10));
  nor2  gate1188(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate1189(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate1190(.a(gate49inter12), .b(gate49inter1), .O(G370));
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate1429(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate1430(.a(gate57inter0), .b(s_126), .O(gate57inter1));
  and2  gate1431(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate1432(.a(s_126), .O(gate57inter3));
  inv1  gate1433(.a(s_127), .O(gate57inter4));
  nand2 gate1434(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate1435(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate1436(.a(G17), .O(gate57inter7));
  inv1  gate1437(.a(G290), .O(gate57inter8));
  nand2 gate1438(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate1439(.a(s_127), .b(gate57inter3), .O(gate57inter10));
  nor2  gate1440(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate1441(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate1442(.a(gate57inter12), .b(gate57inter1), .O(G378));
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate911(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate912(.a(gate63inter0), .b(s_52), .O(gate63inter1));
  and2  gate913(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate914(.a(s_52), .O(gate63inter3));
  inv1  gate915(.a(s_53), .O(gate63inter4));
  nand2 gate916(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate917(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate918(.a(G23), .O(gate63inter7));
  inv1  gate919(.a(G299), .O(gate63inter8));
  nand2 gate920(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate921(.a(s_53), .b(gate63inter3), .O(gate63inter10));
  nor2  gate922(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate923(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate924(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );

  xor2  gate1527(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate1528(.a(gate68inter0), .b(s_140), .O(gate68inter1));
  and2  gate1529(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate1530(.a(s_140), .O(gate68inter3));
  inv1  gate1531(.a(s_141), .O(gate68inter4));
  nand2 gate1532(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate1533(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate1534(.a(G28), .O(gate68inter7));
  inv1  gate1535(.a(G305), .O(gate68inter8));
  nand2 gate1536(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate1537(.a(s_141), .b(gate68inter3), .O(gate68inter10));
  nor2  gate1538(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate1539(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate1540(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );

  xor2  gate631(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate632(.a(gate70inter0), .b(s_12), .O(gate70inter1));
  and2  gate633(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate634(.a(s_12), .O(gate70inter3));
  inv1  gate635(.a(s_13), .O(gate70inter4));
  nand2 gate636(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate637(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate638(.a(G30), .O(gate70inter7));
  inv1  gate639(.a(G308), .O(gate70inter8));
  nand2 gate640(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate641(.a(s_13), .b(gate70inter3), .O(gate70inter10));
  nor2  gate642(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate643(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate644(.a(gate70inter12), .b(gate70inter1), .O(G391));

  xor2  gate1121(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate1122(.a(gate71inter0), .b(s_82), .O(gate71inter1));
  and2  gate1123(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate1124(.a(s_82), .O(gate71inter3));
  inv1  gate1125(.a(s_83), .O(gate71inter4));
  nand2 gate1126(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate1127(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate1128(.a(G31), .O(gate71inter7));
  inv1  gate1129(.a(G311), .O(gate71inter8));
  nand2 gate1130(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate1131(.a(s_83), .b(gate71inter3), .O(gate71inter10));
  nor2  gate1132(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate1133(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate1134(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );

  xor2  gate547(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate548(.a(gate73inter0), .b(s_0), .O(gate73inter1));
  and2  gate549(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate550(.a(s_0), .O(gate73inter3));
  inv1  gate551(.a(s_1), .O(gate73inter4));
  nand2 gate552(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate553(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate554(.a(G1), .O(gate73inter7));
  inv1  gate555(.a(G314), .O(gate73inter8));
  nand2 gate556(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate557(.a(s_1), .b(gate73inter3), .O(gate73inter10));
  nor2  gate558(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate559(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate560(.a(gate73inter12), .b(gate73inter1), .O(G394));

  xor2  gate1009(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate1010(.a(gate74inter0), .b(s_66), .O(gate74inter1));
  and2  gate1011(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate1012(.a(s_66), .O(gate74inter3));
  inv1  gate1013(.a(s_67), .O(gate74inter4));
  nand2 gate1014(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate1015(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate1016(.a(G5), .O(gate74inter7));
  inv1  gate1017(.a(G314), .O(gate74inter8));
  nand2 gate1018(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate1019(.a(s_67), .b(gate74inter3), .O(gate74inter10));
  nor2  gate1020(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate1021(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate1022(.a(gate74inter12), .b(gate74inter1), .O(G395));
nand2 gate75( .a(G9), .b(G317), .O(G396) );

  xor2  gate1443(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate1444(.a(gate76inter0), .b(s_128), .O(gate76inter1));
  and2  gate1445(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate1446(.a(s_128), .O(gate76inter3));
  inv1  gate1447(.a(s_129), .O(gate76inter4));
  nand2 gate1448(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate1449(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate1450(.a(G13), .O(gate76inter7));
  inv1  gate1451(.a(G317), .O(gate76inter8));
  nand2 gate1452(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate1453(.a(s_129), .b(gate76inter3), .O(gate76inter10));
  nor2  gate1454(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate1455(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate1456(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );

  xor2  gate1345(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate1346(.a(gate79inter0), .b(s_114), .O(gate79inter1));
  and2  gate1347(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate1348(.a(s_114), .O(gate79inter3));
  inv1  gate1349(.a(s_115), .O(gate79inter4));
  nand2 gate1350(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate1351(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate1352(.a(G10), .O(gate79inter7));
  inv1  gate1353(.a(G323), .O(gate79inter8));
  nand2 gate1354(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate1355(.a(s_115), .b(gate79inter3), .O(gate79inter10));
  nor2  gate1356(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate1357(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate1358(.a(gate79inter12), .b(gate79inter1), .O(G400));
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );

  xor2  gate673(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate674(.a(gate84inter0), .b(s_18), .O(gate84inter1));
  and2  gate675(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate676(.a(s_18), .O(gate84inter3));
  inv1  gate677(.a(s_19), .O(gate84inter4));
  nand2 gate678(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate679(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate680(.a(G15), .O(gate84inter7));
  inv1  gate681(.a(G329), .O(gate84inter8));
  nand2 gate682(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate683(.a(s_19), .b(gate84inter3), .O(gate84inter10));
  nor2  gate684(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate685(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate686(.a(gate84inter12), .b(gate84inter1), .O(G405));
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate981(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate982(.a(gate86inter0), .b(s_62), .O(gate86inter1));
  and2  gate983(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate984(.a(s_62), .O(gate86inter3));
  inv1  gate985(.a(s_63), .O(gate86inter4));
  nand2 gate986(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate987(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate988(.a(G8), .O(gate86inter7));
  inv1  gate989(.a(G332), .O(gate86inter8));
  nand2 gate990(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate991(.a(s_63), .b(gate86inter3), .O(gate86inter10));
  nor2  gate992(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate993(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate994(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate785(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate786(.a(gate88inter0), .b(s_34), .O(gate88inter1));
  and2  gate787(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate788(.a(s_34), .O(gate88inter3));
  inv1  gate789(.a(s_35), .O(gate88inter4));
  nand2 gate790(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate791(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate792(.a(G16), .O(gate88inter7));
  inv1  gate793(.a(G335), .O(gate88inter8));
  nand2 gate794(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate795(.a(s_35), .b(gate88inter3), .O(gate88inter10));
  nor2  gate796(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate797(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate798(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate1261(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate1262(.a(gate91inter0), .b(s_102), .O(gate91inter1));
  and2  gate1263(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate1264(.a(s_102), .O(gate91inter3));
  inv1  gate1265(.a(s_103), .O(gate91inter4));
  nand2 gate1266(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate1267(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate1268(.a(G25), .O(gate91inter7));
  inv1  gate1269(.a(G341), .O(gate91inter8));
  nand2 gate1270(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate1271(.a(s_103), .b(gate91inter3), .O(gate91inter10));
  nor2  gate1272(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate1273(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate1274(.a(gate91inter12), .b(gate91inter1), .O(G412));

  xor2  gate897(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate898(.a(gate92inter0), .b(s_50), .O(gate92inter1));
  and2  gate899(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate900(.a(s_50), .O(gate92inter3));
  inv1  gate901(.a(s_51), .O(gate92inter4));
  nand2 gate902(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate903(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate904(.a(G29), .O(gate92inter7));
  inv1  gate905(.a(G341), .O(gate92inter8));
  nand2 gate906(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate907(.a(s_51), .b(gate92inter3), .O(gate92inter10));
  nor2  gate908(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate909(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate910(.a(gate92inter12), .b(gate92inter1), .O(G413));

  xor2  gate645(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate646(.a(gate93inter0), .b(s_14), .O(gate93inter1));
  and2  gate647(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate648(.a(s_14), .O(gate93inter3));
  inv1  gate649(.a(s_15), .O(gate93inter4));
  nand2 gate650(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate651(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate652(.a(G18), .O(gate93inter7));
  inv1  gate653(.a(G344), .O(gate93inter8));
  nand2 gate654(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate655(.a(s_15), .b(gate93inter3), .O(gate93inter10));
  nor2  gate656(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate657(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate658(.a(gate93inter12), .b(gate93inter1), .O(G414));
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate1373(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate1374(.a(gate99inter0), .b(s_118), .O(gate99inter1));
  and2  gate1375(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate1376(.a(s_118), .O(gate99inter3));
  inv1  gate1377(.a(s_119), .O(gate99inter4));
  nand2 gate1378(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate1379(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate1380(.a(G27), .O(gate99inter7));
  inv1  gate1381(.a(G353), .O(gate99inter8));
  nand2 gate1382(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate1383(.a(s_119), .b(gate99inter3), .O(gate99inter10));
  nor2  gate1384(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate1385(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate1386(.a(gate99inter12), .b(gate99inter1), .O(G420));

  xor2  gate561(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate562(.a(gate100inter0), .b(s_2), .O(gate100inter1));
  and2  gate563(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate564(.a(s_2), .O(gate100inter3));
  inv1  gate565(.a(s_3), .O(gate100inter4));
  nand2 gate566(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate567(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate568(.a(G31), .O(gate100inter7));
  inv1  gate569(.a(G353), .O(gate100inter8));
  nand2 gate570(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate571(.a(s_3), .b(gate100inter3), .O(gate100inter10));
  nor2  gate572(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate573(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate574(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );

  xor2  gate939(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate940(.a(gate109inter0), .b(s_56), .O(gate109inter1));
  and2  gate941(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate942(.a(s_56), .O(gate109inter3));
  inv1  gate943(.a(s_57), .O(gate109inter4));
  nand2 gate944(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate945(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate946(.a(G370), .O(gate109inter7));
  inv1  gate947(.a(G371), .O(gate109inter8));
  nand2 gate948(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate949(.a(s_57), .b(gate109inter3), .O(gate109inter10));
  nor2  gate950(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate951(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate952(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );

  xor2  gate1107(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate1108(.a(gate111inter0), .b(s_80), .O(gate111inter1));
  and2  gate1109(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate1110(.a(s_80), .O(gate111inter3));
  inv1  gate1111(.a(s_81), .O(gate111inter4));
  nand2 gate1112(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate1113(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate1114(.a(G374), .O(gate111inter7));
  inv1  gate1115(.a(G375), .O(gate111inter8));
  nand2 gate1116(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate1117(.a(s_81), .b(gate111inter3), .O(gate111inter10));
  nor2  gate1118(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate1119(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate1120(.a(gate111inter12), .b(gate111inter1), .O(G444));
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );

  xor2  gate967(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate968(.a(gate114inter0), .b(s_60), .O(gate114inter1));
  and2  gate969(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate970(.a(s_60), .O(gate114inter3));
  inv1  gate971(.a(s_61), .O(gate114inter4));
  nand2 gate972(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate973(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate974(.a(G380), .O(gate114inter7));
  inv1  gate975(.a(G381), .O(gate114inter8));
  nand2 gate976(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate977(.a(s_61), .b(gate114inter3), .O(gate114inter10));
  nor2  gate978(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate979(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate980(.a(gate114inter12), .b(gate114inter1), .O(G453));

  xor2  gate757(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate758(.a(gate115inter0), .b(s_30), .O(gate115inter1));
  and2  gate759(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate760(.a(s_30), .O(gate115inter3));
  inv1  gate761(.a(s_31), .O(gate115inter4));
  nand2 gate762(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate763(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate764(.a(G382), .O(gate115inter7));
  inv1  gate765(.a(G383), .O(gate115inter8));
  nand2 gate766(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate767(.a(s_31), .b(gate115inter3), .O(gate115inter10));
  nor2  gate768(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate769(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate770(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate659(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate660(.a(gate126inter0), .b(s_16), .O(gate126inter1));
  and2  gate661(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate662(.a(s_16), .O(gate126inter3));
  inv1  gate663(.a(s_17), .O(gate126inter4));
  nand2 gate664(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate665(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate666(.a(G404), .O(gate126inter7));
  inv1  gate667(.a(G405), .O(gate126inter8));
  nand2 gate668(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate669(.a(s_17), .b(gate126inter3), .O(gate126inter10));
  nor2  gate670(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate671(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate672(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );

  xor2  gate603(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate604(.a(gate129inter0), .b(s_8), .O(gate129inter1));
  and2  gate605(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate606(.a(s_8), .O(gate129inter3));
  inv1  gate607(.a(s_9), .O(gate129inter4));
  nand2 gate608(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate609(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate610(.a(G410), .O(gate129inter7));
  inv1  gate611(.a(G411), .O(gate129inter8));
  nand2 gate612(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate613(.a(s_9), .b(gate129inter3), .O(gate129inter10));
  nor2  gate614(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate615(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate616(.a(gate129inter12), .b(gate129inter1), .O(G498));
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate1163(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate1164(.a(gate132inter0), .b(s_88), .O(gate132inter1));
  and2  gate1165(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate1166(.a(s_88), .O(gate132inter3));
  inv1  gate1167(.a(s_89), .O(gate132inter4));
  nand2 gate1168(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate1169(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate1170(.a(G416), .O(gate132inter7));
  inv1  gate1171(.a(G417), .O(gate132inter8));
  nand2 gate1172(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate1173(.a(s_89), .b(gate132inter3), .O(gate132inter10));
  nor2  gate1174(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate1175(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate1176(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );

  xor2  gate1471(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate1472(.a(gate139inter0), .b(s_132), .O(gate139inter1));
  and2  gate1473(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate1474(.a(s_132), .O(gate139inter3));
  inv1  gate1475(.a(s_133), .O(gate139inter4));
  nand2 gate1476(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate1477(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate1478(.a(G438), .O(gate139inter7));
  inv1  gate1479(.a(G441), .O(gate139inter8));
  nand2 gate1480(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate1481(.a(s_133), .b(gate139inter3), .O(gate139inter10));
  nor2  gate1482(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate1483(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate1484(.a(gate139inter12), .b(gate139inter1), .O(G528));

  xor2  gate1415(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate1416(.a(gate140inter0), .b(s_124), .O(gate140inter1));
  and2  gate1417(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate1418(.a(s_124), .O(gate140inter3));
  inv1  gate1419(.a(s_125), .O(gate140inter4));
  nand2 gate1420(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate1421(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate1422(.a(G444), .O(gate140inter7));
  inv1  gate1423(.a(G447), .O(gate140inter8));
  nand2 gate1424(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate1425(.a(s_125), .b(gate140inter3), .O(gate140inter10));
  nor2  gate1426(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate1427(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate1428(.a(gate140inter12), .b(gate140inter1), .O(G531));
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate1023(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1024(.a(gate148inter0), .b(s_68), .O(gate148inter1));
  and2  gate1025(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1026(.a(s_68), .O(gate148inter3));
  inv1  gate1027(.a(s_69), .O(gate148inter4));
  nand2 gate1028(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1029(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1030(.a(G492), .O(gate148inter7));
  inv1  gate1031(.a(G495), .O(gate148inter8));
  nand2 gate1032(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1033(.a(s_69), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1034(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1035(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1036(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate827(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate828(.a(gate153inter0), .b(s_40), .O(gate153inter1));
  and2  gate829(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate830(.a(s_40), .O(gate153inter3));
  inv1  gate831(.a(s_41), .O(gate153inter4));
  nand2 gate832(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate833(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate834(.a(G426), .O(gate153inter7));
  inv1  gate835(.a(G522), .O(gate153inter8));
  nand2 gate836(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate837(.a(s_41), .b(gate153inter3), .O(gate153inter10));
  nor2  gate838(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate839(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate840(.a(gate153inter12), .b(gate153inter1), .O(G570));

  xor2  gate1289(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate1290(.a(gate154inter0), .b(s_106), .O(gate154inter1));
  and2  gate1291(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate1292(.a(s_106), .O(gate154inter3));
  inv1  gate1293(.a(s_107), .O(gate154inter4));
  nand2 gate1294(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate1295(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate1296(.a(G429), .O(gate154inter7));
  inv1  gate1297(.a(G522), .O(gate154inter8));
  nand2 gate1298(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate1299(.a(s_107), .b(gate154inter3), .O(gate154inter10));
  nor2  gate1300(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate1301(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate1302(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate1205(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate1206(.a(gate156inter0), .b(s_94), .O(gate156inter1));
  and2  gate1207(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate1208(.a(s_94), .O(gate156inter3));
  inv1  gate1209(.a(s_95), .O(gate156inter4));
  nand2 gate1210(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate1211(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate1212(.a(G435), .O(gate156inter7));
  inv1  gate1213(.a(G525), .O(gate156inter8));
  nand2 gate1214(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate1215(.a(s_95), .b(gate156inter3), .O(gate156inter10));
  nor2  gate1216(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate1217(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate1218(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate841(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate842(.a(gate165inter0), .b(s_42), .O(gate165inter1));
  and2  gate843(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate844(.a(s_42), .O(gate165inter3));
  inv1  gate845(.a(s_43), .O(gate165inter4));
  nand2 gate846(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate847(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate848(.a(G462), .O(gate165inter7));
  inv1  gate849(.a(G540), .O(gate165inter8));
  nand2 gate850(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate851(.a(s_43), .b(gate165inter3), .O(gate165inter10));
  nor2  gate852(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate853(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate854(.a(gate165inter12), .b(gate165inter1), .O(G582));

  xor2  gate1387(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate1388(.a(gate166inter0), .b(s_120), .O(gate166inter1));
  and2  gate1389(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate1390(.a(s_120), .O(gate166inter3));
  inv1  gate1391(.a(s_121), .O(gate166inter4));
  nand2 gate1392(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate1393(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate1394(.a(G465), .O(gate166inter7));
  inv1  gate1395(.a(G540), .O(gate166inter8));
  nand2 gate1396(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate1397(.a(s_121), .b(gate166inter3), .O(gate166inter10));
  nor2  gate1398(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate1399(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate1400(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate1303(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate1304(.a(gate198inter0), .b(s_108), .O(gate198inter1));
  and2  gate1305(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate1306(.a(s_108), .O(gate198inter3));
  inv1  gate1307(.a(s_109), .O(gate198inter4));
  nand2 gate1308(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate1309(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate1310(.a(G596), .O(gate198inter7));
  inv1  gate1311(.a(G597), .O(gate198inter8));
  nand2 gate1312(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate1313(.a(s_109), .b(gate198inter3), .O(gate198inter10));
  nor2  gate1314(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate1315(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate1316(.a(gate198inter12), .b(gate198inter1), .O(G657));
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );

  xor2  gate813(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate814(.a(gate221inter0), .b(s_38), .O(gate221inter1));
  and2  gate815(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate816(.a(s_38), .O(gate221inter3));
  inv1  gate817(.a(s_39), .O(gate221inter4));
  nand2 gate818(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate819(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate820(.a(G622), .O(gate221inter7));
  inv1  gate821(.a(G684), .O(gate221inter8));
  nand2 gate822(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate823(.a(s_39), .b(gate221inter3), .O(gate221inter10));
  nor2  gate824(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate825(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate826(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate855(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate856(.a(gate227inter0), .b(s_44), .O(gate227inter1));
  and2  gate857(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate858(.a(s_44), .O(gate227inter3));
  inv1  gate859(.a(s_45), .O(gate227inter4));
  nand2 gate860(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate861(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate862(.a(G694), .O(gate227inter7));
  inv1  gate863(.a(G695), .O(gate227inter8));
  nand2 gate864(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate865(.a(s_45), .b(gate227inter3), .O(gate227inter10));
  nor2  gate866(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate867(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate868(.a(gate227inter12), .b(gate227inter1), .O(G712));
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate771(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate772(.a(gate258inter0), .b(s_32), .O(gate258inter1));
  and2  gate773(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate774(.a(s_32), .O(gate258inter3));
  inv1  gate775(.a(s_33), .O(gate258inter4));
  nand2 gate776(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate777(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate778(.a(G756), .O(gate258inter7));
  inv1  gate779(.a(G757), .O(gate258inter8));
  nand2 gate780(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate781(.a(s_33), .b(gate258inter3), .O(gate258inter10));
  nor2  gate782(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate783(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate784(.a(gate258inter12), .b(gate258inter1), .O(G773));

  xor2  gate1247(.a(G759), .b(G758), .O(gate259inter0));
  nand2 gate1248(.a(gate259inter0), .b(s_100), .O(gate259inter1));
  and2  gate1249(.a(G759), .b(G758), .O(gate259inter2));
  inv1  gate1250(.a(s_100), .O(gate259inter3));
  inv1  gate1251(.a(s_101), .O(gate259inter4));
  nand2 gate1252(.a(gate259inter4), .b(gate259inter3), .O(gate259inter5));
  nor2  gate1253(.a(gate259inter5), .b(gate259inter2), .O(gate259inter6));
  inv1  gate1254(.a(G758), .O(gate259inter7));
  inv1  gate1255(.a(G759), .O(gate259inter8));
  nand2 gate1256(.a(gate259inter8), .b(gate259inter7), .O(gate259inter9));
  nand2 gate1257(.a(s_101), .b(gate259inter3), .O(gate259inter10));
  nor2  gate1258(.a(gate259inter10), .b(gate259inter9), .O(gate259inter11));
  nor2  gate1259(.a(gate259inter11), .b(gate259inter6), .O(gate259inter12));
  nand2 gate1260(.a(gate259inter12), .b(gate259inter1), .O(G776));
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate1275(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate1276(.a(gate271inter0), .b(s_104), .O(gate271inter1));
  and2  gate1277(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate1278(.a(s_104), .O(gate271inter3));
  inv1  gate1279(.a(s_105), .O(gate271inter4));
  nand2 gate1280(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate1281(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate1282(.a(G660), .O(gate271inter7));
  inv1  gate1283(.a(G788), .O(gate271inter8));
  nand2 gate1284(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate1285(.a(s_105), .b(gate271inter3), .O(gate271inter10));
  nor2  gate1286(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate1287(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate1288(.a(gate271inter12), .b(gate271inter1), .O(G812));

  xor2  gate1457(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate1458(.a(gate272inter0), .b(s_130), .O(gate272inter1));
  and2  gate1459(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate1460(.a(s_130), .O(gate272inter3));
  inv1  gate1461(.a(s_131), .O(gate272inter4));
  nand2 gate1462(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate1463(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate1464(.a(G663), .O(gate272inter7));
  inv1  gate1465(.a(G791), .O(gate272inter8));
  nand2 gate1466(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate1467(.a(s_131), .b(gate272inter3), .O(gate272inter10));
  nor2  gate1468(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate1469(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate1470(.a(gate272inter12), .b(gate272inter1), .O(G815));
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );

  xor2  gate1037(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate1038(.a(gate281inter0), .b(s_70), .O(gate281inter1));
  and2  gate1039(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate1040(.a(s_70), .O(gate281inter3));
  inv1  gate1041(.a(s_71), .O(gate281inter4));
  nand2 gate1042(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate1043(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate1044(.a(G654), .O(gate281inter7));
  inv1  gate1045(.a(G806), .O(gate281inter8));
  nand2 gate1046(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate1047(.a(s_71), .b(gate281inter3), .O(gate281inter10));
  nor2  gate1048(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate1049(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate1050(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );

  xor2  gate1513(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate1514(.a(gate288inter0), .b(s_138), .O(gate288inter1));
  and2  gate1515(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate1516(.a(s_138), .O(gate288inter3));
  inv1  gate1517(.a(s_139), .O(gate288inter4));
  nand2 gate1518(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate1519(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate1520(.a(G791), .O(gate288inter7));
  inv1  gate1521(.a(G815), .O(gate288inter8));
  nand2 gate1522(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate1523(.a(s_139), .b(gate288inter3), .O(gate288inter10));
  nor2  gate1524(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate1525(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate1526(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate925(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate926(.a(gate389inter0), .b(s_54), .O(gate389inter1));
  and2  gate927(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate928(.a(s_54), .O(gate389inter3));
  inv1  gate929(.a(s_55), .O(gate389inter4));
  nand2 gate930(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate931(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate932(.a(G3), .O(gate389inter7));
  inv1  gate933(.a(G1042), .O(gate389inter8));
  nand2 gate934(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate935(.a(s_55), .b(gate389inter3), .O(gate389inter10));
  nor2  gate936(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate937(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate938(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate883(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate884(.a(gate391inter0), .b(s_48), .O(gate391inter1));
  and2  gate885(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate886(.a(s_48), .O(gate391inter3));
  inv1  gate887(.a(s_49), .O(gate391inter4));
  nand2 gate888(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate889(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate890(.a(G5), .O(gate391inter7));
  inv1  gate891(.a(G1048), .O(gate391inter8));
  nand2 gate892(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate893(.a(s_49), .b(gate391inter3), .O(gate391inter10));
  nor2  gate894(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate895(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate896(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );

  xor2  gate1093(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate1094(.a(gate405inter0), .b(s_78), .O(gate405inter1));
  and2  gate1095(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate1096(.a(s_78), .O(gate405inter3));
  inv1  gate1097(.a(s_79), .O(gate405inter4));
  nand2 gate1098(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate1099(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate1100(.a(G19), .O(gate405inter7));
  inv1  gate1101(.a(G1090), .O(gate405inter8));
  nand2 gate1102(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate1103(.a(s_79), .b(gate405inter3), .O(gate405inter10));
  nor2  gate1104(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate1105(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate1106(.a(gate405inter12), .b(gate405inter1), .O(G1186));
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate1219(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate1220(.a(gate407inter0), .b(s_96), .O(gate407inter1));
  and2  gate1221(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate1222(.a(s_96), .O(gate407inter3));
  inv1  gate1223(.a(s_97), .O(gate407inter4));
  nand2 gate1224(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate1225(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate1226(.a(G21), .O(gate407inter7));
  inv1  gate1227(.a(G1096), .O(gate407inter8));
  nand2 gate1228(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate1229(.a(s_97), .b(gate407inter3), .O(gate407inter10));
  nor2  gate1230(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate1231(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate1232(.a(gate407inter12), .b(gate407inter1), .O(G1192));

  xor2  gate715(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate716(.a(gate408inter0), .b(s_24), .O(gate408inter1));
  and2  gate717(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate718(.a(s_24), .O(gate408inter3));
  inv1  gate719(.a(s_25), .O(gate408inter4));
  nand2 gate720(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate721(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate722(.a(G22), .O(gate408inter7));
  inv1  gate723(.a(G1099), .O(gate408inter8));
  nand2 gate724(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate725(.a(s_25), .b(gate408inter3), .O(gate408inter10));
  nor2  gate726(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate727(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate728(.a(gate408inter12), .b(gate408inter1), .O(G1195));
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );

  xor2  gate617(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate618(.a(gate412inter0), .b(s_10), .O(gate412inter1));
  and2  gate619(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate620(.a(s_10), .O(gate412inter3));
  inv1  gate621(.a(s_11), .O(gate412inter4));
  nand2 gate622(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate623(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate624(.a(G26), .O(gate412inter7));
  inv1  gate625(.a(G1111), .O(gate412inter8));
  nand2 gate626(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate627(.a(s_11), .b(gate412inter3), .O(gate412inter10));
  nor2  gate628(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate629(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate630(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate589(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate590(.a(gate415inter0), .b(s_6), .O(gate415inter1));
  and2  gate591(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate592(.a(s_6), .O(gate415inter3));
  inv1  gate593(.a(s_7), .O(gate415inter4));
  nand2 gate594(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate595(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate596(.a(G29), .O(gate415inter7));
  inv1  gate597(.a(G1120), .O(gate415inter8));
  nand2 gate598(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate599(.a(s_7), .b(gate415inter3), .O(gate415inter10));
  nor2  gate600(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate601(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate602(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );

  xor2  gate1149(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate1150(.a(gate426inter0), .b(s_86), .O(gate426inter1));
  and2  gate1151(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate1152(.a(s_86), .O(gate426inter3));
  inv1  gate1153(.a(s_87), .O(gate426inter4));
  nand2 gate1154(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate1155(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate1156(.a(G1045), .O(gate426inter7));
  inv1  gate1157(.a(G1141), .O(gate426inter8));
  nand2 gate1158(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate1159(.a(s_87), .b(gate426inter3), .O(gate426inter10));
  nor2  gate1160(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate1161(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate1162(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );

  xor2  gate1499(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate1500(.a(gate428inter0), .b(s_136), .O(gate428inter1));
  and2  gate1501(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate1502(.a(s_136), .O(gate428inter3));
  inv1  gate1503(.a(s_137), .O(gate428inter4));
  nand2 gate1504(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate1505(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate1506(.a(G1048), .O(gate428inter7));
  inv1  gate1507(.a(G1144), .O(gate428inter8));
  nand2 gate1508(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate1509(.a(s_137), .b(gate428inter3), .O(gate428inter10));
  nor2  gate1510(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate1511(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate1512(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );

  xor2  gate1401(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate1402(.a(gate431inter0), .b(s_122), .O(gate431inter1));
  and2  gate1403(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate1404(.a(s_122), .O(gate431inter3));
  inv1  gate1405(.a(s_123), .O(gate431inter4));
  nand2 gate1406(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate1407(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate1408(.a(G7), .O(gate431inter7));
  inv1  gate1409(.a(G1150), .O(gate431inter8));
  nand2 gate1410(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate1411(.a(s_123), .b(gate431inter3), .O(gate431inter10));
  nor2  gate1412(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate1413(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate1414(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate1065(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate1066(.a(gate439inter0), .b(s_74), .O(gate439inter1));
  and2  gate1067(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate1068(.a(s_74), .O(gate439inter3));
  inv1  gate1069(.a(s_75), .O(gate439inter4));
  nand2 gate1070(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate1071(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate1072(.a(G11), .O(gate439inter7));
  inv1  gate1073(.a(G1162), .O(gate439inter8));
  nand2 gate1074(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate1075(.a(s_75), .b(gate439inter3), .O(gate439inter10));
  nor2  gate1076(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate1077(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate1078(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate953(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate954(.a(gate444inter0), .b(s_58), .O(gate444inter1));
  and2  gate955(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate956(.a(s_58), .O(gate444inter3));
  inv1  gate957(.a(s_59), .O(gate444inter4));
  nand2 gate958(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate959(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate960(.a(G1072), .O(gate444inter7));
  inv1  gate961(.a(G1168), .O(gate444inter8));
  nand2 gate962(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate963(.a(s_59), .b(gate444inter3), .O(gate444inter10));
  nor2  gate964(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate965(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate966(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );

  xor2  gate869(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate870(.a(gate446inter0), .b(s_46), .O(gate446inter1));
  and2  gate871(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate872(.a(s_46), .O(gate446inter3));
  inv1  gate873(.a(s_47), .O(gate446inter4));
  nand2 gate874(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate875(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate876(.a(G1075), .O(gate446inter7));
  inv1  gate877(.a(G1171), .O(gate446inter8));
  nand2 gate878(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate879(.a(s_47), .b(gate446inter3), .O(gate446inter10));
  nor2  gate880(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate881(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate882(.a(gate446inter12), .b(gate446inter1), .O(G1255));
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate575(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate576(.a(gate448inter0), .b(s_4), .O(gate448inter1));
  and2  gate577(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate578(.a(s_4), .O(gate448inter3));
  inv1  gate579(.a(s_5), .O(gate448inter4));
  nand2 gate580(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate581(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate582(.a(G1078), .O(gate448inter7));
  inv1  gate583(.a(G1174), .O(gate448inter8));
  nand2 gate584(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate585(.a(s_5), .b(gate448inter3), .O(gate448inter10));
  nor2  gate586(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate587(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate588(.a(gate448inter12), .b(gate448inter1), .O(G1257));
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate799(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate800(.a(gate453inter0), .b(s_36), .O(gate453inter1));
  and2  gate801(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate802(.a(s_36), .O(gate453inter3));
  inv1  gate803(.a(s_37), .O(gate453inter4));
  nand2 gate804(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate805(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate806(.a(G18), .O(gate453inter7));
  inv1  gate807(.a(G1183), .O(gate453inter8));
  nand2 gate808(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate809(.a(s_37), .b(gate453inter3), .O(gate453inter10));
  nor2  gate810(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate811(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate812(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate743(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate744(.a(gate464inter0), .b(s_28), .O(gate464inter1));
  and2  gate745(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate746(.a(s_28), .O(gate464inter3));
  inv1  gate747(.a(s_29), .O(gate464inter4));
  nand2 gate748(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate749(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate750(.a(G1102), .O(gate464inter7));
  inv1  gate751(.a(G1198), .O(gate464inter8));
  nand2 gate752(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate753(.a(s_29), .b(gate464inter3), .O(gate464inter10));
  nor2  gate754(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate755(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate756(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );

  xor2  gate1191(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate1192(.a(gate476inter0), .b(s_92), .O(gate476inter1));
  and2  gate1193(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate1194(.a(s_92), .O(gate476inter3));
  inv1  gate1195(.a(s_93), .O(gate476inter4));
  nand2 gate1196(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate1197(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate1198(.a(G1120), .O(gate476inter7));
  inv1  gate1199(.a(G1216), .O(gate476inter8));
  nand2 gate1200(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate1201(.a(s_93), .b(gate476inter3), .O(gate476inter10));
  nor2  gate1202(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate1203(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate1204(.a(gate476inter12), .b(gate476inter1), .O(G1285));

  xor2  gate1359(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate1360(.a(gate477inter0), .b(s_116), .O(gate477inter1));
  and2  gate1361(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate1362(.a(s_116), .O(gate477inter3));
  inv1  gate1363(.a(s_117), .O(gate477inter4));
  nand2 gate1364(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate1365(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate1366(.a(G30), .O(gate477inter7));
  inv1  gate1367(.a(G1219), .O(gate477inter8));
  nand2 gate1368(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate1369(.a(s_117), .b(gate477inter3), .O(gate477inter10));
  nor2  gate1370(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate1371(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate1372(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );

  xor2  gate1051(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate1052(.a(gate486inter0), .b(s_72), .O(gate486inter1));
  and2  gate1053(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate1054(.a(s_72), .O(gate486inter3));
  inv1  gate1055(.a(s_73), .O(gate486inter4));
  nand2 gate1056(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate1057(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate1058(.a(G1234), .O(gate486inter7));
  inv1  gate1059(.a(G1235), .O(gate486inter8));
  nand2 gate1060(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate1061(.a(s_73), .b(gate486inter3), .O(gate486inter10));
  nor2  gate1062(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate1063(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate1064(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate995(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate996(.a(gate490inter0), .b(s_64), .O(gate490inter1));
  and2  gate997(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate998(.a(s_64), .O(gate490inter3));
  inv1  gate999(.a(s_65), .O(gate490inter4));
  nand2 gate1000(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate1001(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate1002(.a(G1242), .O(gate490inter7));
  inv1  gate1003(.a(G1243), .O(gate490inter8));
  nand2 gate1004(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate1005(.a(s_65), .b(gate490inter3), .O(gate490inter10));
  nor2  gate1006(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate1007(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate1008(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate1485(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate1486(.a(gate496inter0), .b(s_134), .O(gate496inter1));
  and2  gate1487(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate1488(.a(s_134), .O(gate496inter3));
  inv1  gate1489(.a(s_135), .O(gate496inter4));
  nand2 gate1490(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate1491(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate1492(.a(G1254), .O(gate496inter7));
  inv1  gate1493(.a(G1255), .O(gate496inter8));
  nand2 gate1494(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate1495(.a(s_135), .b(gate496inter3), .O(gate496inter10));
  nor2  gate1496(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate1497(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate1498(.a(gate496inter12), .b(gate496inter1), .O(G1305));
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );

  xor2  gate701(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate702(.a(gate498inter0), .b(s_22), .O(gate498inter1));
  and2  gate703(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate704(.a(s_22), .O(gate498inter3));
  inv1  gate705(.a(s_23), .O(gate498inter4));
  nand2 gate706(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate707(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate708(.a(G1258), .O(gate498inter7));
  inv1  gate709(.a(G1259), .O(gate498inter8));
  nand2 gate710(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate711(.a(s_23), .b(gate498inter3), .O(gate498inter10));
  nor2  gate712(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate713(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate714(.a(gate498inter12), .b(gate498inter1), .O(G1307));
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate687(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate688(.a(gate504inter0), .b(s_20), .O(gate504inter1));
  and2  gate689(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate690(.a(s_20), .O(gate504inter3));
  inv1  gate691(.a(s_21), .O(gate504inter4));
  nand2 gate692(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate693(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate694(.a(G1270), .O(gate504inter7));
  inv1  gate695(.a(G1271), .O(gate504inter8));
  nand2 gate696(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate697(.a(s_21), .b(gate504inter3), .O(gate504inter10));
  nor2  gate698(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate699(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate700(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate1331(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate1332(.a(gate509inter0), .b(s_112), .O(gate509inter1));
  and2  gate1333(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate1334(.a(s_112), .O(gate509inter3));
  inv1  gate1335(.a(s_113), .O(gate509inter4));
  nand2 gate1336(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate1337(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate1338(.a(G1280), .O(gate509inter7));
  inv1  gate1339(.a(G1281), .O(gate509inter8));
  nand2 gate1340(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate1341(.a(s_113), .b(gate509inter3), .O(gate509inter10));
  nor2  gate1342(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate1343(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate1344(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule