module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281, s_282, s_283, s_284, s_285, s_286, s_287, s_288, s_289, s_290, s_291, s_292, s_293, s_294, s_295, s_296, s_297, s_298, s_299, s_300, s_301, s_302, s_303, s_304, s_305, s_306, s_307, s_308, s_309, s_310, s_311, s_312, s_313, s_314, s_315, s_316, s_317, s_318, s_319, s_320, s_321, s_322, s_323, s_324, s_325, s_326, s_327, s_328, s_329, s_330, s_331;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate176inter0, gate176inter1, gate176inter2, gate176inter3, gate176inter4, gate176inter5, gate176inter6, gate176inter7, gate176inter8, gate176inter9, gate176inter10, gate176inter11, gate176inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate476inter0, gate476inter1, gate476inter2, gate476inter3, gate476inter4, gate476inter5, gate476inter6, gate476inter7, gate476inter8, gate476inter9, gate476inter10, gate476inter11, gate476inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate108inter0, gate108inter1, gate108inter2, gate108inter3, gate108inter4, gate108inter5, gate108inter6, gate108inter7, gate108inter8, gate108inter9, gate108inter10, gate108inter11, gate108inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate481inter0, gate481inter1, gate481inter2, gate481inter3, gate481inter4, gate481inter5, gate481inter6, gate481inter7, gate481inter8, gate481inter9, gate481inter10, gate481inter11, gate481inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate445inter0, gate445inter1, gate445inter2, gate445inter3, gate445inter4, gate445inter5, gate445inter6, gate445inter7, gate445inter8, gate445inter9, gate445inter10, gate445inter11, gate445inter12, gate250inter0, gate250inter1, gate250inter2, gate250inter3, gate250inter4, gate250inter5, gate250inter6, gate250inter7, gate250inter8, gate250inter9, gate250inter10, gate250inter11, gate250inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate456inter0, gate456inter1, gate456inter2, gate456inter3, gate456inter4, gate456inter5, gate456inter6, gate456inter7, gate456inter8, gate456inter9, gate456inter10, gate456inter11, gate456inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate49inter0, gate49inter1, gate49inter2, gate49inter3, gate49inter4, gate49inter5, gate49inter6, gate49inter7, gate49inter8, gate49inter9, gate49inter10, gate49inter11, gate49inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate226inter0, gate226inter1, gate226inter2, gate226inter3, gate226inter4, gate226inter5, gate226inter6, gate226inter7, gate226inter8, gate226inter9, gate226inter10, gate226inter11, gate226inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate470inter0, gate470inter1, gate470inter2, gate470inter3, gate470inter4, gate470inter5, gate470inter6, gate470inter7, gate470inter8, gate470inter9, gate470inter10, gate470inter11, gate470inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate389inter0, gate389inter1, gate389inter2, gate389inter3, gate389inter4, gate389inter5, gate389inter6, gate389inter7, gate389inter8, gate389inter9, gate389inter10, gate389inter11, gate389inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate109inter0, gate109inter1, gate109inter2, gate109inter3, gate109inter4, gate109inter5, gate109inter6, gate109inter7, gate109inter8, gate109inter9, gate109inter10, gate109inter11, gate109inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate503inter0, gate503inter1, gate503inter2, gate503inter3, gate503inter4, gate503inter5, gate503inter6, gate503inter7, gate503inter8, gate503inter9, gate503inter10, gate503inter11, gate503inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate507inter0, gate507inter1, gate507inter2, gate507inter3, gate507inter4, gate507inter5, gate507inter6, gate507inter7, gate507inter8, gate507inter9, gate507inter10, gate507inter11, gate507inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate414inter0, gate414inter1, gate414inter2, gate414inter3, gate414inter4, gate414inter5, gate414inter6, gate414inter7, gate414inter8, gate414inter9, gate414inter10, gate414inter11, gate414inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate93inter0, gate93inter1, gate93inter2, gate93inter3, gate93inter4, gate93inter5, gate93inter6, gate93inter7, gate93inter8, gate93inter9, gate93inter10, gate93inter11, gate93inter12, gate436inter0, gate436inter1, gate436inter2, gate436inter3, gate436inter4, gate436inter5, gate436inter6, gate436inter7, gate436inter8, gate436inter9, gate436inter10, gate436inter11, gate436inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12, gate45inter0, gate45inter1, gate45inter2, gate45inter3, gate45inter4, gate45inter5, gate45inter6, gate45inter7, gate45inter8, gate45inter9, gate45inter10, gate45inter11, gate45inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate434inter0, gate434inter1, gate434inter2, gate434inter3, gate434inter4, gate434inter5, gate434inter6, gate434inter7, gate434inter8, gate434inter9, gate434inter10, gate434inter11, gate434inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate2507(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate2508(.a(gate12inter0), .b(s_280), .O(gate12inter1));
  and2  gate2509(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate2510(.a(s_280), .O(gate12inter3));
  inv1  gate2511(.a(s_281), .O(gate12inter4));
  nand2 gate2512(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate2513(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate2514(.a(G7), .O(gate12inter7));
  inv1  gate2515(.a(G8), .O(gate12inter8));
  nand2 gate2516(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate2517(.a(s_281), .b(gate12inter3), .O(gate12inter10));
  nor2  gate2518(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate2519(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate2520(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );

  xor2  gate1919(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate1920(.a(gate14inter0), .b(s_196), .O(gate14inter1));
  and2  gate1921(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate1922(.a(s_196), .O(gate14inter3));
  inv1  gate1923(.a(s_197), .O(gate14inter4));
  nand2 gate1924(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate1925(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate1926(.a(G11), .O(gate14inter7));
  inv1  gate1927(.a(G12), .O(gate14inter8));
  nand2 gate1928(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate1929(.a(s_197), .b(gate14inter3), .O(gate14inter10));
  nor2  gate1930(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate1931(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate1932(.a(gate14inter12), .b(gate14inter1), .O(G281));
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate2423(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate2424(.a(gate16inter0), .b(s_268), .O(gate16inter1));
  and2  gate2425(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate2426(.a(s_268), .O(gate16inter3));
  inv1  gate2427(.a(s_269), .O(gate16inter4));
  nand2 gate2428(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate2429(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate2430(.a(G15), .O(gate16inter7));
  inv1  gate2431(.a(G16), .O(gate16inter8));
  nand2 gate2432(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate2433(.a(s_269), .b(gate16inter3), .O(gate16inter10));
  nor2  gate2434(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate2435(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate2436(.a(gate16inter12), .b(gate16inter1), .O(G287));

  xor2  gate2283(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate2284(.a(gate17inter0), .b(s_248), .O(gate17inter1));
  and2  gate2285(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate2286(.a(s_248), .O(gate17inter3));
  inv1  gate2287(.a(s_249), .O(gate17inter4));
  nand2 gate2288(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate2289(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate2290(.a(G17), .O(gate17inter7));
  inv1  gate2291(.a(G18), .O(gate17inter8));
  nand2 gate2292(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate2293(.a(s_249), .b(gate17inter3), .O(gate17inter10));
  nor2  gate2294(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate2295(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate2296(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate2045(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate2046(.a(gate22inter0), .b(s_214), .O(gate22inter1));
  and2  gate2047(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate2048(.a(s_214), .O(gate22inter3));
  inv1  gate2049(.a(s_215), .O(gate22inter4));
  nand2 gate2050(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate2051(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate2052(.a(G27), .O(gate22inter7));
  inv1  gate2053(.a(G28), .O(gate22inter8));
  nand2 gate2054(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate2055(.a(s_215), .b(gate22inter3), .O(gate22inter10));
  nor2  gate2056(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate2057(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate2058(.a(gate22inter12), .b(gate22inter1), .O(G305));

  xor2  gate2171(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate2172(.a(gate23inter0), .b(s_232), .O(gate23inter1));
  and2  gate2173(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate2174(.a(s_232), .O(gate23inter3));
  inv1  gate2175(.a(s_233), .O(gate23inter4));
  nand2 gate2176(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate2177(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate2178(.a(G29), .O(gate23inter7));
  inv1  gate2179(.a(G30), .O(gate23inter8));
  nand2 gate2180(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate2181(.a(s_233), .b(gate23inter3), .O(gate23inter10));
  nor2  gate2182(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate2183(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate2184(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate1989(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate1990(.a(gate25inter0), .b(s_206), .O(gate25inter1));
  and2  gate1991(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate1992(.a(s_206), .O(gate25inter3));
  inv1  gate1993(.a(s_207), .O(gate25inter4));
  nand2 gate1994(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate1995(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate1996(.a(G1), .O(gate25inter7));
  inv1  gate1997(.a(G5), .O(gate25inter8));
  nand2 gate1998(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate1999(.a(s_207), .b(gate25inter3), .O(gate25inter10));
  nor2  gate2000(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate2001(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate2002(.a(gate25inter12), .b(gate25inter1), .O(G314));

  xor2  gate659(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate660(.a(gate26inter0), .b(s_16), .O(gate26inter1));
  and2  gate661(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate662(.a(s_16), .O(gate26inter3));
  inv1  gate663(.a(s_17), .O(gate26inter4));
  nand2 gate664(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate665(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate666(.a(G9), .O(gate26inter7));
  inv1  gate667(.a(G13), .O(gate26inter8));
  nand2 gate668(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate669(.a(s_17), .b(gate26inter3), .O(gate26inter10));
  nor2  gate670(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate671(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate672(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );

  xor2  gate1611(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate1612(.a(gate32inter0), .b(s_152), .O(gate32inter1));
  and2  gate1613(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate1614(.a(s_152), .O(gate32inter3));
  inv1  gate1615(.a(s_153), .O(gate32inter4));
  nand2 gate1616(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate1617(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate1618(.a(G12), .O(gate32inter7));
  inv1  gate1619(.a(G16), .O(gate32inter8));
  nand2 gate1620(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate1621(.a(s_153), .b(gate32inter3), .O(gate32inter10));
  nor2  gate1622(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate1623(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate1624(.a(gate32inter12), .b(gate32inter1), .O(G335));

  xor2  gate1443(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate1444(.a(gate33inter0), .b(s_128), .O(gate33inter1));
  and2  gate1445(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate1446(.a(s_128), .O(gate33inter3));
  inv1  gate1447(.a(s_129), .O(gate33inter4));
  nand2 gate1448(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate1449(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate1450(.a(G17), .O(gate33inter7));
  inv1  gate1451(.a(G21), .O(gate33inter8));
  nand2 gate1452(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate1453(.a(s_129), .b(gate33inter3), .O(gate33inter10));
  nor2  gate1454(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate1455(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate1456(.a(gate33inter12), .b(gate33inter1), .O(G338));
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );

  xor2  gate855(.a(G30), .b(G26), .O(gate36inter0));
  nand2 gate856(.a(gate36inter0), .b(s_44), .O(gate36inter1));
  and2  gate857(.a(G30), .b(G26), .O(gate36inter2));
  inv1  gate858(.a(s_44), .O(gate36inter3));
  inv1  gate859(.a(s_45), .O(gate36inter4));
  nand2 gate860(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate861(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate862(.a(G26), .O(gate36inter7));
  inv1  gate863(.a(G30), .O(gate36inter8));
  nand2 gate864(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate865(.a(s_45), .b(gate36inter3), .O(gate36inter10));
  nor2  gate866(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate867(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate868(.a(gate36inter12), .b(gate36inter1), .O(G347));
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate2185(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate2186(.a(gate39inter0), .b(s_234), .O(gate39inter1));
  and2  gate2187(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate2188(.a(s_234), .O(gate39inter3));
  inv1  gate2189(.a(s_235), .O(gate39inter4));
  nand2 gate2190(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate2191(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate2192(.a(G20), .O(gate39inter7));
  inv1  gate2193(.a(G24), .O(gate39inter8));
  nand2 gate2194(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate2195(.a(s_235), .b(gate39inter3), .O(gate39inter10));
  nor2  gate2196(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate2197(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate2198(.a(gate39inter12), .b(gate39inter1), .O(G356));
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate2521(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate2522(.a(gate43inter0), .b(s_282), .O(gate43inter1));
  and2  gate2523(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate2524(.a(s_282), .O(gate43inter3));
  inv1  gate2525(.a(s_283), .O(gate43inter4));
  nand2 gate2526(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate2527(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate2528(.a(G3), .O(gate43inter7));
  inv1  gate2529(.a(G269), .O(gate43inter8));
  nand2 gate2530(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate2531(.a(s_283), .b(gate43inter3), .O(gate43inter10));
  nor2  gate2532(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate2533(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate2534(.a(gate43inter12), .b(gate43inter1), .O(G364));

  xor2  gate2773(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate2774(.a(gate44inter0), .b(s_318), .O(gate44inter1));
  and2  gate2775(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate2776(.a(s_318), .O(gate44inter3));
  inv1  gate2777(.a(s_319), .O(gate44inter4));
  nand2 gate2778(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate2779(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate2780(.a(G4), .O(gate44inter7));
  inv1  gate2781(.a(G269), .O(gate44inter8));
  nand2 gate2782(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate2783(.a(s_319), .b(gate44inter3), .O(gate44inter10));
  nor2  gate2784(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate2785(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate2786(.a(gate44inter12), .b(gate44inter1), .O(G365));

  xor2  gate2465(.a(G272), .b(G5), .O(gate45inter0));
  nand2 gate2466(.a(gate45inter0), .b(s_274), .O(gate45inter1));
  and2  gate2467(.a(G272), .b(G5), .O(gate45inter2));
  inv1  gate2468(.a(s_274), .O(gate45inter3));
  inv1  gate2469(.a(s_275), .O(gate45inter4));
  nand2 gate2470(.a(gate45inter4), .b(gate45inter3), .O(gate45inter5));
  nor2  gate2471(.a(gate45inter5), .b(gate45inter2), .O(gate45inter6));
  inv1  gate2472(.a(G5), .O(gate45inter7));
  inv1  gate2473(.a(G272), .O(gate45inter8));
  nand2 gate2474(.a(gate45inter8), .b(gate45inter7), .O(gate45inter9));
  nand2 gate2475(.a(s_275), .b(gate45inter3), .O(gate45inter10));
  nor2  gate2476(.a(gate45inter10), .b(gate45inter9), .O(gate45inter11));
  nor2  gate2477(.a(gate45inter11), .b(gate45inter6), .O(gate45inter12));
  nand2 gate2478(.a(gate45inter12), .b(gate45inter1), .O(G366));
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );

  xor2  gate1219(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate1220(.a(gate48inter0), .b(s_96), .O(gate48inter1));
  and2  gate1221(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate1222(.a(s_96), .O(gate48inter3));
  inv1  gate1223(.a(s_97), .O(gate48inter4));
  nand2 gate1224(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate1225(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate1226(.a(G8), .O(gate48inter7));
  inv1  gate1227(.a(G275), .O(gate48inter8));
  nand2 gate1228(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate1229(.a(s_97), .b(gate48inter3), .O(gate48inter10));
  nor2  gate1230(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate1231(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate1232(.a(gate48inter12), .b(gate48inter1), .O(G369));

  xor2  gate1541(.a(G278), .b(G9), .O(gate49inter0));
  nand2 gate1542(.a(gate49inter0), .b(s_142), .O(gate49inter1));
  and2  gate1543(.a(G278), .b(G9), .O(gate49inter2));
  inv1  gate1544(.a(s_142), .O(gate49inter3));
  inv1  gate1545(.a(s_143), .O(gate49inter4));
  nand2 gate1546(.a(gate49inter4), .b(gate49inter3), .O(gate49inter5));
  nor2  gate1547(.a(gate49inter5), .b(gate49inter2), .O(gate49inter6));
  inv1  gate1548(.a(G9), .O(gate49inter7));
  inv1  gate1549(.a(G278), .O(gate49inter8));
  nand2 gate1550(.a(gate49inter8), .b(gate49inter7), .O(gate49inter9));
  nand2 gate1551(.a(s_143), .b(gate49inter3), .O(gate49inter10));
  nor2  gate1552(.a(gate49inter10), .b(gate49inter9), .O(gate49inter11));
  nor2  gate1553(.a(gate49inter11), .b(gate49inter6), .O(gate49inter12));
  nand2 gate1554(.a(gate49inter12), .b(gate49inter1), .O(G370));
nand2 gate50( .a(G10), .b(G278), .O(G371) );

  xor2  gate2255(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate2256(.a(gate51inter0), .b(s_244), .O(gate51inter1));
  and2  gate2257(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate2258(.a(s_244), .O(gate51inter3));
  inv1  gate2259(.a(s_245), .O(gate51inter4));
  nand2 gate2260(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate2261(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate2262(.a(G11), .O(gate51inter7));
  inv1  gate2263(.a(G281), .O(gate51inter8));
  nand2 gate2264(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate2265(.a(s_245), .b(gate51inter3), .O(gate51inter10));
  nor2  gate2266(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate2267(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate2268(.a(gate51inter12), .b(gate51inter1), .O(G372));

  xor2  gate2619(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate2620(.a(gate52inter0), .b(s_296), .O(gate52inter1));
  and2  gate2621(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate2622(.a(s_296), .O(gate52inter3));
  inv1  gate2623(.a(s_297), .O(gate52inter4));
  nand2 gate2624(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate2625(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate2626(.a(G12), .O(gate52inter7));
  inv1  gate2627(.a(G281), .O(gate52inter8));
  nand2 gate2628(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate2629(.a(s_297), .b(gate52inter3), .O(gate52inter10));
  nor2  gate2630(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate2631(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate2632(.a(gate52inter12), .b(gate52inter1), .O(G373));

  xor2  gate2661(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate2662(.a(gate53inter0), .b(s_302), .O(gate53inter1));
  and2  gate2663(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate2664(.a(s_302), .O(gate53inter3));
  inv1  gate2665(.a(s_303), .O(gate53inter4));
  nand2 gate2666(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate2667(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate2668(.a(G13), .O(gate53inter7));
  inv1  gate2669(.a(G284), .O(gate53inter8));
  nand2 gate2670(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate2671(.a(s_303), .b(gate53inter3), .O(gate53inter10));
  nor2  gate2672(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate2673(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate2674(.a(gate53inter12), .b(gate53inter1), .O(G374));
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate939(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate940(.a(gate59inter0), .b(s_56), .O(gate59inter1));
  and2  gate941(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate942(.a(s_56), .O(gate59inter3));
  inv1  gate943(.a(s_57), .O(gate59inter4));
  nand2 gate944(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate945(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate946(.a(G19), .O(gate59inter7));
  inv1  gate947(.a(G293), .O(gate59inter8));
  nand2 gate948(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate949(.a(s_57), .b(gate59inter3), .O(gate59inter10));
  nor2  gate950(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate951(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate952(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate1289(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate1290(.a(gate67inter0), .b(s_106), .O(gate67inter1));
  and2  gate1291(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate1292(.a(s_106), .O(gate67inter3));
  inv1  gate1293(.a(s_107), .O(gate67inter4));
  nand2 gate1294(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate1295(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate1296(.a(G27), .O(gate67inter7));
  inv1  gate1297(.a(G305), .O(gate67inter8));
  nand2 gate1298(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate1299(.a(s_107), .b(gate67inter3), .O(gate67inter10));
  nor2  gate1300(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate1301(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate1302(.a(gate67inter12), .b(gate67inter1), .O(G388));

  xor2  gate2395(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate2396(.a(gate68inter0), .b(s_264), .O(gate68inter1));
  and2  gate2397(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate2398(.a(s_264), .O(gate68inter3));
  inv1  gate2399(.a(s_265), .O(gate68inter4));
  nand2 gate2400(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate2401(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate2402(.a(G28), .O(gate68inter7));
  inv1  gate2403(.a(G305), .O(gate68inter8));
  nand2 gate2404(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate2405(.a(s_265), .b(gate68inter3), .O(gate68inter10));
  nor2  gate2406(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate2407(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate2408(.a(gate68inter12), .b(gate68inter1), .O(G389));

  xor2  gate603(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate604(.a(gate69inter0), .b(s_8), .O(gate69inter1));
  and2  gate605(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate606(.a(s_8), .O(gate69inter3));
  inv1  gate607(.a(s_9), .O(gate69inter4));
  nand2 gate608(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate609(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate610(.a(G29), .O(gate69inter7));
  inv1  gate611(.a(G308), .O(gate69inter8));
  nand2 gate612(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate613(.a(s_9), .b(gate69inter3), .O(gate69inter10));
  nor2  gate614(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate615(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate616(.a(gate69inter12), .b(gate69inter1), .O(G390));

  xor2  gate1625(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate1626(.a(gate70inter0), .b(s_154), .O(gate70inter1));
  and2  gate1627(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate1628(.a(s_154), .O(gate70inter3));
  inv1  gate1629(.a(s_155), .O(gate70inter4));
  nand2 gate1630(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate1631(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate1632(.a(G30), .O(gate70inter7));
  inv1  gate1633(.a(G308), .O(gate70inter8));
  nand2 gate1634(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate1635(.a(s_155), .b(gate70inter3), .O(gate70inter10));
  nor2  gate1636(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate1637(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate1638(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );

  xor2  gate1569(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate1570(.a(gate72inter0), .b(s_146), .O(gate72inter1));
  and2  gate1571(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate1572(.a(s_146), .O(gate72inter3));
  inv1  gate1573(.a(s_147), .O(gate72inter4));
  nand2 gate1574(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate1575(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate1576(.a(G32), .O(gate72inter7));
  inv1  gate1577(.a(G311), .O(gate72inter8));
  nand2 gate1578(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate1579(.a(s_147), .b(gate72inter3), .O(gate72inter10));
  nor2  gate1580(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate1581(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate1582(.a(gate72inter12), .b(gate72inter1), .O(G393));

  xor2  gate1135(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate1136(.a(gate73inter0), .b(s_84), .O(gate73inter1));
  and2  gate1137(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate1138(.a(s_84), .O(gate73inter3));
  inv1  gate1139(.a(s_85), .O(gate73inter4));
  nand2 gate1140(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate1141(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate1142(.a(G1), .O(gate73inter7));
  inv1  gate1143(.a(G314), .O(gate73inter8));
  nand2 gate1144(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate1145(.a(s_85), .b(gate73inter3), .O(gate73inter10));
  nor2  gate1146(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate1147(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate1148(.a(gate73inter12), .b(gate73inter1), .O(G394));
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate911(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate912(.a(gate75inter0), .b(s_52), .O(gate75inter1));
  and2  gate913(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate914(.a(s_52), .O(gate75inter3));
  inv1  gate915(.a(s_53), .O(gate75inter4));
  nand2 gate916(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate917(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate918(.a(G9), .O(gate75inter7));
  inv1  gate919(.a(G317), .O(gate75inter8));
  nand2 gate920(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate921(.a(s_53), .b(gate75inter3), .O(gate75inter10));
  nor2  gate922(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate923(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate924(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate1387(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate1388(.a(gate77inter0), .b(s_120), .O(gate77inter1));
  and2  gate1389(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate1390(.a(s_120), .O(gate77inter3));
  inv1  gate1391(.a(s_121), .O(gate77inter4));
  nand2 gate1392(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate1393(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate1394(.a(G2), .O(gate77inter7));
  inv1  gate1395(.a(G320), .O(gate77inter8));
  nand2 gate1396(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate1397(.a(s_121), .b(gate77inter3), .O(gate77inter10));
  nor2  gate1398(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate1399(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate1400(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );

  xor2  gate2143(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate2144(.a(gate83inter0), .b(s_228), .O(gate83inter1));
  and2  gate2145(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate2146(.a(s_228), .O(gate83inter3));
  inv1  gate2147(.a(s_229), .O(gate83inter4));
  nand2 gate2148(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate2149(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate2150(.a(G11), .O(gate83inter7));
  inv1  gate2151(.a(G329), .O(gate83inter8));
  nand2 gate2152(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate2153(.a(s_229), .b(gate83inter3), .O(gate83inter10));
  nor2  gate2154(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate2155(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate2156(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate1401(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate1402(.a(gate86inter0), .b(s_122), .O(gate86inter1));
  and2  gate1403(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate1404(.a(s_122), .O(gate86inter3));
  inv1  gate1405(.a(s_123), .O(gate86inter4));
  nand2 gate1406(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate1407(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate1408(.a(G8), .O(gate86inter7));
  inv1  gate1409(.a(G332), .O(gate86inter8));
  nand2 gate1410(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate1411(.a(s_123), .b(gate86inter3), .O(gate86inter10));
  nor2  gate1412(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate1413(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate1414(.a(gate86inter12), .b(gate86inter1), .O(G407));

  xor2  gate2339(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate2340(.a(gate87inter0), .b(s_256), .O(gate87inter1));
  and2  gate2341(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate2342(.a(s_256), .O(gate87inter3));
  inv1  gate2343(.a(s_257), .O(gate87inter4));
  nand2 gate2344(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate2345(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate2346(.a(G12), .O(gate87inter7));
  inv1  gate2347(.a(G335), .O(gate87inter8));
  nand2 gate2348(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate2349(.a(s_257), .b(gate87inter3), .O(gate87inter10));
  nor2  gate2350(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate2351(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate2352(.a(gate87inter12), .b(gate87inter1), .O(G408));

  xor2  gate981(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate982(.a(gate88inter0), .b(s_62), .O(gate88inter1));
  and2  gate983(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate984(.a(s_62), .O(gate88inter3));
  inv1  gate985(.a(s_63), .O(gate88inter4));
  nand2 gate986(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate987(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate988(.a(G16), .O(gate88inter7));
  inv1  gate989(.a(G335), .O(gate88inter8));
  nand2 gate990(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate991(.a(s_63), .b(gate88inter3), .O(gate88inter10));
  nor2  gate992(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate993(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate994(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );

  xor2  gate1653(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate1654(.a(gate92inter0), .b(s_158), .O(gate92inter1));
  and2  gate1655(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate1656(.a(s_158), .O(gate92inter3));
  inv1  gate1657(.a(s_159), .O(gate92inter4));
  nand2 gate1658(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate1659(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate1660(.a(G29), .O(gate92inter7));
  inv1  gate1661(.a(G341), .O(gate92inter8));
  nand2 gate1662(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate1663(.a(s_159), .b(gate92inter3), .O(gate92inter10));
  nor2  gate1664(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate1665(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate1666(.a(gate92inter12), .b(gate92inter1), .O(G413));

  xor2  gate2297(.a(G344), .b(G18), .O(gate93inter0));
  nand2 gate2298(.a(gate93inter0), .b(s_250), .O(gate93inter1));
  and2  gate2299(.a(G344), .b(G18), .O(gate93inter2));
  inv1  gate2300(.a(s_250), .O(gate93inter3));
  inv1  gate2301(.a(s_251), .O(gate93inter4));
  nand2 gate2302(.a(gate93inter4), .b(gate93inter3), .O(gate93inter5));
  nor2  gate2303(.a(gate93inter5), .b(gate93inter2), .O(gate93inter6));
  inv1  gate2304(.a(G18), .O(gate93inter7));
  inv1  gate2305(.a(G344), .O(gate93inter8));
  nand2 gate2306(.a(gate93inter8), .b(gate93inter7), .O(gate93inter9));
  nand2 gate2307(.a(s_251), .b(gate93inter3), .O(gate93inter10));
  nor2  gate2308(.a(gate93inter10), .b(gate93inter9), .O(gate93inter11));
  nor2  gate2309(.a(gate93inter11), .b(gate93inter6), .O(gate93inter12));
  nand2 gate2310(.a(gate93inter12), .b(gate93inter1), .O(G414));
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate1723(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate1724(.a(gate95inter0), .b(s_168), .O(gate95inter1));
  and2  gate1725(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate1726(.a(s_168), .O(gate95inter3));
  inv1  gate1727(.a(s_169), .O(gate95inter4));
  nand2 gate1728(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate1729(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate1730(.a(G26), .O(gate95inter7));
  inv1  gate1731(.a(G347), .O(gate95inter8));
  nand2 gate1732(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate1733(.a(s_169), .b(gate95inter3), .O(gate95inter10));
  nor2  gate1734(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate1735(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate1736(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate1639(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate1640(.a(gate104inter0), .b(s_156), .O(gate104inter1));
  and2  gate1641(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate1642(.a(s_156), .O(gate104inter3));
  inv1  gate1643(.a(s_157), .O(gate104inter4));
  nand2 gate1644(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate1645(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate1646(.a(G32), .O(gate104inter7));
  inv1  gate1647(.a(G359), .O(gate104inter8));
  nand2 gate1648(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate1649(.a(s_157), .b(gate104inter3), .O(gate104inter10));
  nor2  gate1650(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate1651(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate1652(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );

  xor2  gate813(.a(G369), .b(G368), .O(gate108inter0));
  nand2 gate814(.a(gate108inter0), .b(s_38), .O(gate108inter1));
  and2  gate815(.a(G369), .b(G368), .O(gate108inter2));
  inv1  gate816(.a(s_38), .O(gate108inter3));
  inv1  gate817(.a(s_39), .O(gate108inter4));
  nand2 gate818(.a(gate108inter4), .b(gate108inter3), .O(gate108inter5));
  nor2  gate819(.a(gate108inter5), .b(gate108inter2), .O(gate108inter6));
  inv1  gate820(.a(G368), .O(gate108inter7));
  inv1  gate821(.a(G369), .O(gate108inter8));
  nand2 gate822(.a(gate108inter8), .b(gate108inter7), .O(gate108inter9));
  nand2 gate823(.a(s_39), .b(gate108inter3), .O(gate108inter10));
  nor2  gate824(.a(gate108inter10), .b(gate108inter9), .O(gate108inter11));
  nor2  gate825(.a(gate108inter11), .b(gate108inter6), .O(gate108inter12));
  nand2 gate826(.a(gate108inter12), .b(gate108inter1), .O(G435));

  xor2  gate2003(.a(G371), .b(G370), .O(gate109inter0));
  nand2 gate2004(.a(gate109inter0), .b(s_208), .O(gate109inter1));
  and2  gate2005(.a(G371), .b(G370), .O(gate109inter2));
  inv1  gate2006(.a(s_208), .O(gate109inter3));
  inv1  gate2007(.a(s_209), .O(gate109inter4));
  nand2 gate2008(.a(gate109inter4), .b(gate109inter3), .O(gate109inter5));
  nor2  gate2009(.a(gate109inter5), .b(gate109inter2), .O(gate109inter6));
  inv1  gate2010(.a(G370), .O(gate109inter7));
  inv1  gate2011(.a(G371), .O(gate109inter8));
  nand2 gate2012(.a(gate109inter8), .b(gate109inter7), .O(gate109inter9));
  nand2 gate2013(.a(s_209), .b(gate109inter3), .O(gate109inter10));
  nor2  gate2014(.a(gate109inter10), .b(gate109inter9), .O(gate109inter11));
  nor2  gate2015(.a(gate109inter11), .b(gate109inter6), .O(gate109inter12));
  nand2 gate2016(.a(gate109inter12), .b(gate109inter1), .O(G438));
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate2269(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate2270(.a(gate124inter0), .b(s_246), .O(gate124inter1));
  and2  gate2271(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate2272(.a(s_246), .O(gate124inter3));
  inv1  gate2273(.a(s_247), .O(gate124inter4));
  nand2 gate2274(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate2275(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate2276(.a(G400), .O(gate124inter7));
  inv1  gate2277(.a(G401), .O(gate124inter8));
  nand2 gate2278(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate2279(.a(s_247), .b(gate124inter3), .O(gate124inter10));
  nor2  gate2280(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate2281(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate2282(.a(gate124inter12), .b(gate124inter1), .O(G483));
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate1331(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate1332(.a(gate132inter0), .b(s_112), .O(gate132inter1));
  and2  gate1333(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate1334(.a(s_112), .O(gate132inter3));
  inv1  gate1335(.a(s_113), .O(gate132inter4));
  nand2 gate1336(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate1337(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate1338(.a(G416), .O(gate132inter7));
  inv1  gate1339(.a(G417), .O(gate132inter8));
  nand2 gate1340(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate1341(.a(s_113), .b(gate132inter3), .O(gate132inter10));
  nor2  gate1342(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate1343(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate1344(.a(gate132inter12), .b(gate132inter1), .O(G507));

  xor2  gate2199(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate2200(.a(gate133inter0), .b(s_236), .O(gate133inter1));
  and2  gate2201(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate2202(.a(s_236), .O(gate133inter3));
  inv1  gate2203(.a(s_237), .O(gate133inter4));
  nand2 gate2204(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate2205(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate2206(.a(G418), .O(gate133inter7));
  inv1  gate2207(.a(G419), .O(gate133inter8));
  nand2 gate2208(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate2209(.a(s_237), .b(gate133inter3), .O(gate133inter10));
  nor2  gate2210(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate2211(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate2212(.a(gate133inter12), .b(gate133inter1), .O(G510));
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate2437(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate2438(.a(gate135inter0), .b(s_270), .O(gate135inter1));
  and2  gate2439(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate2440(.a(s_270), .O(gate135inter3));
  inv1  gate2441(.a(s_271), .O(gate135inter4));
  nand2 gate2442(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate2443(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate2444(.a(G422), .O(gate135inter7));
  inv1  gate2445(.a(G423), .O(gate135inter8));
  nand2 gate2446(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate2447(.a(s_271), .b(gate135inter3), .O(gate135inter10));
  nor2  gate2448(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate2449(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate2450(.a(gate135inter12), .b(gate135inter1), .O(G516));

  xor2  gate1947(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate1948(.a(gate136inter0), .b(s_200), .O(gate136inter1));
  and2  gate1949(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate1950(.a(s_200), .O(gate136inter3));
  inv1  gate1951(.a(s_201), .O(gate136inter4));
  nand2 gate1952(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate1953(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate1954(.a(G424), .O(gate136inter7));
  inv1  gate1955(.a(G425), .O(gate136inter8));
  nand2 gate1956(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate1957(.a(s_201), .b(gate136inter3), .O(gate136inter10));
  nor2  gate1958(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate1959(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate1960(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );

  xor2  gate1681(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate1682(.a(gate138inter0), .b(s_162), .O(gate138inter1));
  and2  gate1683(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate1684(.a(s_162), .O(gate138inter3));
  inv1  gate1685(.a(s_163), .O(gate138inter4));
  nand2 gate1686(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate1687(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate1688(.a(G432), .O(gate138inter7));
  inv1  gate1689(.a(G435), .O(gate138inter8));
  nand2 gate1690(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate1691(.a(s_163), .b(gate138inter3), .O(gate138inter10));
  nor2  gate1692(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate1693(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate1694(.a(gate138inter12), .b(gate138inter1), .O(G525));

  xor2  gate2325(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate2326(.a(gate139inter0), .b(s_254), .O(gate139inter1));
  and2  gate2327(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate2328(.a(s_254), .O(gate139inter3));
  inv1  gate2329(.a(s_255), .O(gate139inter4));
  nand2 gate2330(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate2331(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate2332(.a(G438), .O(gate139inter7));
  inv1  gate2333(.a(G441), .O(gate139inter8));
  nand2 gate2334(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate2335(.a(s_255), .b(gate139inter3), .O(gate139inter10));
  nor2  gate2336(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate2337(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate2338(.a(gate139inter12), .b(gate139inter1), .O(G528));
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate645(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate646(.a(gate143inter0), .b(s_14), .O(gate143inter1));
  and2  gate647(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate648(.a(s_14), .O(gate143inter3));
  inv1  gate649(.a(s_15), .O(gate143inter4));
  nand2 gate650(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate651(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate652(.a(G462), .O(gate143inter7));
  inv1  gate653(.a(G465), .O(gate143inter8));
  nand2 gate654(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate655(.a(s_15), .b(gate143inter3), .O(gate143inter10));
  nor2  gate656(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate657(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate658(.a(gate143inter12), .b(gate143inter1), .O(G540));
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );

  xor2  gate715(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate716(.a(gate146inter0), .b(s_24), .O(gate146inter1));
  and2  gate717(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate718(.a(s_24), .O(gate146inter3));
  inv1  gate719(.a(s_25), .O(gate146inter4));
  nand2 gate720(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate721(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate722(.a(G480), .O(gate146inter7));
  inv1  gate723(.a(G483), .O(gate146inter8));
  nand2 gate724(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate725(.a(s_25), .b(gate146inter3), .O(gate146inter10));
  nor2  gate726(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate727(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate728(.a(gate146inter12), .b(gate146inter1), .O(G549));

  xor2  gate1247(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate1248(.a(gate147inter0), .b(s_100), .O(gate147inter1));
  and2  gate1249(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate1250(.a(s_100), .O(gate147inter3));
  inv1  gate1251(.a(s_101), .O(gate147inter4));
  nand2 gate1252(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate1253(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate1254(.a(G486), .O(gate147inter7));
  inv1  gate1255(.a(G489), .O(gate147inter8));
  nand2 gate1256(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate1257(.a(s_101), .b(gate147inter3), .O(gate147inter10));
  nor2  gate1258(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate1259(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate1260(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate687(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate688(.a(gate149inter0), .b(s_20), .O(gate149inter1));
  and2  gate689(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate690(.a(s_20), .O(gate149inter3));
  inv1  gate691(.a(s_21), .O(gate149inter4));
  nand2 gate692(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate693(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate694(.a(G498), .O(gate149inter7));
  inv1  gate695(.a(G501), .O(gate149inter8));
  nand2 gate696(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate697(.a(s_21), .b(gate149inter3), .O(gate149inter10));
  nor2  gate698(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate699(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate700(.a(gate149inter12), .b(gate149inter1), .O(G558));

  xor2  gate771(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate772(.a(gate150inter0), .b(s_32), .O(gate150inter1));
  and2  gate773(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate774(.a(s_32), .O(gate150inter3));
  inv1  gate775(.a(s_33), .O(gate150inter4));
  nand2 gate776(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate777(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate778(.a(G504), .O(gate150inter7));
  inv1  gate779(.a(G507), .O(gate150inter8));
  nand2 gate780(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate781(.a(s_33), .b(gate150inter3), .O(gate150inter10));
  nor2  gate782(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate783(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate784(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );

  xor2  gate1205(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate1206(.a(gate154inter0), .b(s_94), .O(gate154inter1));
  and2  gate1207(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate1208(.a(s_94), .O(gate154inter3));
  inv1  gate1209(.a(s_95), .O(gate154inter4));
  nand2 gate1210(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate1211(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate1212(.a(G429), .O(gate154inter7));
  inv1  gate1213(.a(G522), .O(gate154inter8));
  nand2 gate1214(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate1215(.a(s_95), .b(gate154inter3), .O(gate154inter10));
  nor2  gate1216(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate1217(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate1218(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate2675(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate2676(.a(gate157inter0), .b(s_304), .O(gate157inter1));
  and2  gate2677(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate2678(.a(s_304), .O(gate157inter3));
  inv1  gate2679(.a(s_305), .O(gate157inter4));
  nand2 gate2680(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate2681(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate2682(.a(G438), .O(gate157inter7));
  inv1  gate2683(.a(G528), .O(gate157inter8));
  nand2 gate2684(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate2685(.a(s_305), .b(gate157inter3), .O(gate157inter10));
  nor2  gate2686(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate2687(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate2688(.a(gate157inter12), .b(gate157inter1), .O(G574));

  xor2  gate1695(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate1696(.a(gate158inter0), .b(s_164), .O(gate158inter1));
  and2  gate1697(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate1698(.a(s_164), .O(gate158inter3));
  inv1  gate1699(.a(s_165), .O(gate158inter4));
  nand2 gate1700(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate1701(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate1702(.a(G441), .O(gate158inter7));
  inv1  gate1703(.a(G528), .O(gate158inter8));
  nand2 gate1704(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate1705(.a(s_165), .b(gate158inter3), .O(gate158inter10));
  nor2  gate1706(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate1707(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate1708(.a(gate158inter12), .b(gate158inter1), .O(G575));
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );

  xor2  gate673(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate674(.a(gate163inter0), .b(s_18), .O(gate163inter1));
  and2  gate675(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate676(.a(s_18), .O(gate163inter3));
  inv1  gate677(.a(s_19), .O(gate163inter4));
  nand2 gate678(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate679(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate680(.a(G456), .O(gate163inter7));
  inv1  gate681(.a(G537), .O(gate163inter8));
  nand2 gate682(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate683(.a(s_19), .b(gate163inter3), .O(gate163inter10));
  nor2  gate684(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate685(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate686(.a(gate163inter12), .b(gate163inter1), .O(G580));

  xor2  gate729(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate730(.a(gate164inter0), .b(s_26), .O(gate164inter1));
  and2  gate731(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate732(.a(s_26), .O(gate164inter3));
  inv1  gate733(.a(s_27), .O(gate164inter4));
  nand2 gate734(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate735(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate736(.a(G459), .O(gate164inter7));
  inv1  gate737(.a(G537), .O(gate164inter8));
  nand2 gate738(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate739(.a(s_27), .b(gate164inter3), .O(gate164inter10));
  nor2  gate740(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate741(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate742(.a(gate164inter12), .b(gate164inter1), .O(G581));

  xor2  gate1751(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate1752(.a(gate165inter0), .b(s_172), .O(gate165inter1));
  and2  gate1753(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate1754(.a(s_172), .O(gate165inter3));
  inv1  gate1755(.a(s_173), .O(gate165inter4));
  nand2 gate1756(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate1757(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate1758(.a(G462), .O(gate165inter7));
  inv1  gate1759(.a(G540), .O(gate165inter8));
  nand2 gate1760(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate1761(.a(s_173), .b(gate165inter3), .O(gate165inter10));
  nor2  gate1762(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate1763(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate1764(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate2591(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate2592(.a(gate170inter0), .b(s_292), .O(gate170inter1));
  and2  gate2593(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate2594(.a(s_292), .O(gate170inter3));
  inv1  gate2595(.a(s_293), .O(gate170inter4));
  nand2 gate2596(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate2597(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate2598(.a(G477), .O(gate170inter7));
  inv1  gate2599(.a(G546), .O(gate170inter8));
  nand2 gate2600(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate2601(.a(s_293), .b(gate170inter3), .O(gate170inter10));
  nor2  gate2602(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate2603(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate2604(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate1905(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate1906(.a(gate172inter0), .b(s_194), .O(gate172inter1));
  and2  gate1907(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate1908(.a(s_194), .O(gate172inter3));
  inv1  gate1909(.a(s_195), .O(gate172inter4));
  nand2 gate1910(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate1911(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate1912(.a(G483), .O(gate172inter7));
  inv1  gate1913(.a(G549), .O(gate172inter8));
  nand2 gate1914(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate1915(.a(s_195), .b(gate172inter3), .O(gate172inter10));
  nor2  gate1916(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate1917(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate1918(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );

  xor2  gate561(.a(G555), .b(G495), .O(gate176inter0));
  nand2 gate562(.a(gate176inter0), .b(s_2), .O(gate176inter1));
  and2  gate563(.a(G555), .b(G495), .O(gate176inter2));
  inv1  gate564(.a(s_2), .O(gate176inter3));
  inv1  gate565(.a(s_3), .O(gate176inter4));
  nand2 gate566(.a(gate176inter4), .b(gate176inter3), .O(gate176inter5));
  nor2  gate567(.a(gate176inter5), .b(gate176inter2), .O(gate176inter6));
  inv1  gate568(.a(G495), .O(gate176inter7));
  inv1  gate569(.a(G555), .O(gate176inter8));
  nand2 gate570(.a(gate176inter8), .b(gate176inter7), .O(gate176inter9));
  nand2 gate571(.a(s_3), .b(gate176inter3), .O(gate176inter10));
  nor2  gate572(.a(gate176inter10), .b(gate176inter9), .O(gate176inter11));
  nor2  gate573(.a(gate176inter11), .b(gate176inter6), .O(gate176inter12));
  nand2 gate574(.a(gate176inter12), .b(gate176inter1), .O(G593));
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate897(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate898(.a(gate178inter0), .b(s_50), .O(gate178inter1));
  and2  gate899(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate900(.a(s_50), .O(gate178inter3));
  inv1  gate901(.a(s_51), .O(gate178inter4));
  nand2 gate902(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate903(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate904(.a(G501), .O(gate178inter7));
  inv1  gate905(.a(G558), .O(gate178inter8));
  nand2 gate906(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate907(.a(s_51), .b(gate178inter3), .O(gate178inter10));
  nor2  gate908(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate909(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate910(.a(gate178inter12), .b(gate178inter1), .O(G595));
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate1583(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate1584(.a(gate180inter0), .b(s_148), .O(gate180inter1));
  and2  gate1585(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate1586(.a(s_148), .O(gate180inter3));
  inv1  gate1587(.a(s_149), .O(gate180inter4));
  nand2 gate1588(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate1589(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate1590(.a(G507), .O(gate180inter7));
  inv1  gate1591(.a(G561), .O(gate180inter8));
  nand2 gate1592(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate1593(.a(s_149), .b(gate180inter3), .O(gate180inter10));
  nor2  gate1594(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate1595(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate1596(.a(gate180inter12), .b(gate180inter1), .O(G597));
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate2745(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate2746(.a(gate183inter0), .b(s_314), .O(gate183inter1));
  and2  gate2747(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate2748(.a(s_314), .O(gate183inter3));
  inv1  gate2749(.a(s_315), .O(gate183inter4));
  nand2 gate2750(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate2751(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate2752(.a(G516), .O(gate183inter7));
  inv1  gate2753(.a(G567), .O(gate183inter8));
  nand2 gate2754(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate2755(.a(s_315), .b(gate183inter3), .O(gate183inter10));
  nor2  gate2756(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate2757(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate2758(.a(gate183inter12), .b(gate183inter1), .O(G600));

  xor2  gate1429(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate1430(.a(gate184inter0), .b(s_126), .O(gate184inter1));
  and2  gate1431(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate1432(.a(s_126), .O(gate184inter3));
  inv1  gate1433(.a(s_127), .O(gate184inter4));
  nand2 gate1434(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate1435(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate1436(.a(G519), .O(gate184inter7));
  inv1  gate1437(.a(G567), .O(gate184inter8));
  nand2 gate1438(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate1439(.a(s_127), .b(gate184inter3), .O(gate184inter10));
  nor2  gate1440(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate1441(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate1442(.a(gate184inter12), .b(gate184inter1), .O(G601));
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate1275(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate1276(.a(gate186inter0), .b(s_104), .O(gate186inter1));
  and2  gate1277(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate1278(.a(s_104), .O(gate186inter3));
  inv1  gate1279(.a(s_105), .O(gate186inter4));
  nand2 gate1280(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate1281(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate1282(.a(G572), .O(gate186inter7));
  inv1  gate1283(.a(G573), .O(gate186inter8));
  nand2 gate1284(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate1285(.a(s_105), .b(gate186inter3), .O(gate186inter10));
  nor2  gate1286(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate1287(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate1288(.a(gate186inter12), .b(gate186inter1), .O(G607));

  xor2  gate1933(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate1934(.a(gate187inter0), .b(s_198), .O(gate187inter1));
  and2  gate1935(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate1936(.a(s_198), .O(gate187inter3));
  inv1  gate1937(.a(s_199), .O(gate187inter4));
  nand2 gate1938(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate1939(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate1940(.a(G574), .O(gate187inter7));
  inv1  gate1941(.a(G575), .O(gate187inter8));
  nand2 gate1942(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate1943(.a(s_199), .b(gate187inter3), .O(gate187inter10));
  nor2  gate1944(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate1945(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate1946(.a(gate187inter12), .b(gate187inter1), .O(G612));
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );

  xor2  gate2815(.a(G581), .b(G580), .O(gate190inter0));
  nand2 gate2816(.a(gate190inter0), .b(s_324), .O(gate190inter1));
  and2  gate2817(.a(G581), .b(G580), .O(gate190inter2));
  inv1  gate2818(.a(s_324), .O(gate190inter3));
  inv1  gate2819(.a(s_325), .O(gate190inter4));
  nand2 gate2820(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate2821(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate2822(.a(G580), .O(gate190inter7));
  inv1  gate2823(.a(G581), .O(gate190inter8));
  nand2 gate2824(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate2825(.a(s_325), .b(gate190inter3), .O(gate190inter10));
  nor2  gate2826(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate2827(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate2828(.a(gate190inter12), .b(gate190inter1), .O(G627));

  xor2  gate827(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate828(.a(gate191inter0), .b(s_40), .O(gate191inter1));
  and2  gate829(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate830(.a(s_40), .O(gate191inter3));
  inv1  gate831(.a(s_41), .O(gate191inter4));
  nand2 gate832(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate833(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate834(.a(G582), .O(gate191inter7));
  inv1  gate835(.a(G583), .O(gate191inter8));
  nand2 gate836(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate837(.a(s_41), .b(gate191inter3), .O(gate191inter10));
  nor2  gate838(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate839(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate840(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );

  xor2  gate1709(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate1710(.a(gate199inter0), .b(s_166), .O(gate199inter1));
  and2  gate1711(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate1712(.a(s_166), .O(gate199inter3));
  inv1  gate1713(.a(s_167), .O(gate199inter4));
  nand2 gate1714(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate1715(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate1716(.a(G598), .O(gate199inter7));
  inv1  gate1717(.a(G599), .O(gate199inter8));
  nand2 gate1718(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate1719(.a(s_167), .b(gate199inter3), .O(gate199inter10));
  nor2  gate1720(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate1721(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate1722(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate785(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate786(.a(gate201inter0), .b(s_34), .O(gate201inter1));
  and2  gate787(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate788(.a(s_34), .O(gate201inter3));
  inv1  gate789(.a(s_35), .O(gate201inter4));
  nand2 gate790(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate791(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate792(.a(G602), .O(gate201inter7));
  inv1  gate793(.a(G607), .O(gate201inter8));
  nand2 gate794(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate795(.a(s_35), .b(gate201inter3), .O(gate201inter10));
  nor2  gate796(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate797(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate798(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate869(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate870(.a(gate203inter0), .b(s_46), .O(gate203inter1));
  and2  gate871(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate872(.a(s_46), .O(gate203inter3));
  inv1  gate873(.a(s_47), .O(gate203inter4));
  nand2 gate874(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate875(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate876(.a(G602), .O(gate203inter7));
  inv1  gate877(.a(G612), .O(gate203inter8));
  nand2 gate878(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate879(.a(s_47), .b(gate203inter3), .O(gate203inter10));
  nor2  gate880(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate881(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate882(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate2451(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate2452(.a(gate205inter0), .b(s_272), .O(gate205inter1));
  and2  gate2453(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate2454(.a(s_272), .O(gate205inter3));
  inv1  gate2455(.a(s_273), .O(gate205inter4));
  nand2 gate2456(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate2457(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate2458(.a(G622), .O(gate205inter7));
  inv1  gate2459(.a(G627), .O(gate205inter8));
  nand2 gate2460(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate2461(.a(s_273), .b(gate205inter3), .O(gate205inter10));
  nor2  gate2462(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate2463(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate2464(.a(gate205inter12), .b(gate205inter1), .O(G678));
nand2 gate206( .a(G632), .b(G637), .O(G681) );

  xor2  gate2857(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate2858(.a(gate207inter0), .b(s_330), .O(gate207inter1));
  and2  gate2859(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate2860(.a(s_330), .O(gate207inter3));
  inv1  gate2861(.a(s_331), .O(gate207inter4));
  nand2 gate2862(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate2863(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate2864(.a(G622), .O(gate207inter7));
  inv1  gate2865(.a(G632), .O(gate207inter8));
  nand2 gate2866(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate2867(.a(s_331), .b(gate207inter3), .O(gate207inter10));
  nor2  gate2868(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate2869(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate2870(.a(gate207inter12), .b(gate207inter1), .O(G684));
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate2717(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate2718(.a(gate211inter0), .b(s_310), .O(gate211inter1));
  and2  gate2719(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate2720(.a(s_310), .O(gate211inter3));
  inv1  gate2721(.a(s_311), .O(gate211inter4));
  nand2 gate2722(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate2723(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate2724(.a(G612), .O(gate211inter7));
  inv1  gate2725(.a(G669), .O(gate211inter8));
  nand2 gate2726(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate2727(.a(s_311), .b(gate211inter3), .O(gate211inter10));
  nor2  gate2728(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate2729(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate2730(.a(gate211inter12), .b(gate211inter1), .O(G692));

  xor2  gate1149(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate1150(.a(gate212inter0), .b(s_86), .O(gate212inter1));
  and2  gate1151(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate1152(.a(s_86), .O(gate212inter3));
  inv1  gate1153(.a(s_87), .O(gate212inter4));
  nand2 gate1154(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate1155(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate1156(.a(G617), .O(gate212inter7));
  inv1  gate1157(.a(G669), .O(gate212inter8));
  nand2 gate1158(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate1159(.a(s_87), .b(gate212inter3), .O(gate212inter10));
  nor2  gate1160(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate1161(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate1162(.a(gate212inter12), .b(gate212inter1), .O(G693));
nand2 gate213( .a(G602), .b(G672), .O(G694) );

  xor2  gate2535(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate2536(.a(gate214inter0), .b(s_284), .O(gate214inter1));
  and2  gate2537(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate2538(.a(s_284), .O(gate214inter3));
  inv1  gate2539(.a(s_285), .O(gate214inter4));
  nand2 gate2540(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate2541(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate2542(.a(G612), .O(gate214inter7));
  inv1  gate2543(.a(G672), .O(gate214inter8));
  nand2 gate2544(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate2545(.a(s_285), .b(gate214inter3), .O(gate214inter10));
  nor2  gate2546(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate2547(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate2548(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );

  xor2  gate1821(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate1822(.a(gate221inter0), .b(s_182), .O(gate221inter1));
  and2  gate1823(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate1824(.a(s_182), .O(gate221inter3));
  inv1  gate1825(.a(s_183), .O(gate221inter4));
  nand2 gate1826(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate1827(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate1828(.a(G622), .O(gate221inter7));
  inv1  gate1829(.a(G684), .O(gate221inter8));
  nand2 gate1830(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate1831(.a(s_183), .b(gate221inter3), .O(gate221inter10));
  nor2  gate1832(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate1833(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate1834(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate1499(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate1500(.a(gate223inter0), .b(s_136), .O(gate223inter1));
  and2  gate1501(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate1502(.a(s_136), .O(gate223inter3));
  inv1  gate1503(.a(s_137), .O(gate223inter4));
  nand2 gate1504(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate1505(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate1506(.a(G627), .O(gate223inter7));
  inv1  gate1507(.a(G687), .O(gate223inter8));
  nand2 gate1508(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate1509(.a(s_137), .b(gate223inter3), .O(gate223inter10));
  nor2  gate1510(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate1511(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate1512(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );

  xor2  gate1121(.a(G691), .b(G690), .O(gate225inter0));
  nand2 gate1122(.a(gate225inter0), .b(s_82), .O(gate225inter1));
  and2  gate1123(.a(G691), .b(G690), .O(gate225inter2));
  inv1  gate1124(.a(s_82), .O(gate225inter3));
  inv1  gate1125(.a(s_83), .O(gate225inter4));
  nand2 gate1126(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate1127(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate1128(.a(G690), .O(gate225inter7));
  inv1  gate1129(.a(G691), .O(gate225inter8));
  nand2 gate1130(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate1131(.a(s_83), .b(gate225inter3), .O(gate225inter10));
  nor2  gate1132(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate1133(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate1134(.a(gate225inter12), .b(gate225inter1), .O(G706));

  xor2  gate1667(.a(G693), .b(G692), .O(gate226inter0));
  nand2 gate1668(.a(gate226inter0), .b(s_160), .O(gate226inter1));
  and2  gate1669(.a(G693), .b(G692), .O(gate226inter2));
  inv1  gate1670(.a(s_160), .O(gate226inter3));
  inv1  gate1671(.a(s_161), .O(gate226inter4));
  nand2 gate1672(.a(gate226inter4), .b(gate226inter3), .O(gate226inter5));
  nor2  gate1673(.a(gate226inter5), .b(gate226inter2), .O(gate226inter6));
  inv1  gate1674(.a(G692), .O(gate226inter7));
  inv1  gate1675(.a(G693), .O(gate226inter8));
  nand2 gate1676(.a(gate226inter8), .b(gate226inter7), .O(gate226inter9));
  nand2 gate1677(.a(s_161), .b(gate226inter3), .O(gate226inter10));
  nor2  gate1678(.a(gate226inter10), .b(gate226inter9), .O(gate226inter11));
  nor2  gate1679(.a(gate226inter11), .b(gate226inter6), .O(gate226inter12));
  nand2 gate1680(.a(gate226inter12), .b(gate226inter1), .O(G709));
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate1527(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate1528(.a(gate228inter0), .b(s_140), .O(gate228inter1));
  and2  gate1529(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate1530(.a(s_140), .O(gate228inter3));
  inv1  gate1531(.a(s_141), .O(gate228inter4));
  nand2 gate1532(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate1533(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate1534(.a(G696), .O(gate228inter7));
  inv1  gate1535(.a(G697), .O(gate228inter8));
  nand2 gate1536(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate1537(.a(s_141), .b(gate228inter3), .O(gate228inter10));
  nor2  gate1538(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate1539(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate1540(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate2031(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate2032(.a(gate231inter0), .b(s_212), .O(gate231inter1));
  and2  gate2033(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate2034(.a(s_212), .O(gate231inter3));
  inv1  gate2035(.a(s_213), .O(gate231inter4));
  nand2 gate2036(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate2037(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate2038(.a(G702), .O(gate231inter7));
  inv1  gate2039(.a(G703), .O(gate231inter8));
  nand2 gate2040(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate2041(.a(s_213), .b(gate231inter3), .O(gate231inter10));
  nor2  gate2042(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate2043(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate2044(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );

  xor2  gate1597(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate1598(.a(gate235inter0), .b(s_150), .O(gate235inter1));
  and2  gate1599(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate1600(.a(s_150), .O(gate235inter3));
  inv1  gate1601(.a(s_151), .O(gate235inter4));
  nand2 gate1602(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate1603(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate1604(.a(G248), .O(gate235inter7));
  inv1  gate1605(.a(G724), .O(gate235inter8));
  nand2 gate1606(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate1607(.a(s_151), .b(gate235inter3), .O(gate235inter10));
  nor2  gate1608(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate1609(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate1610(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate2703(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate2704(.a(gate240inter0), .b(s_308), .O(gate240inter1));
  and2  gate2705(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate2706(.a(s_308), .O(gate240inter3));
  inv1  gate2707(.a(s_309), .O(gate240inter4));
  nand2 gate2708(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate2709(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate2710(.a(G263), .O(gate240inter7));
  inv1  gate2711(.a(G715), .O(gate240inter8));
  nand2 gate2712(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate2713(.a(s_309), .b(gate240inter3), .O(gate240inter10));
  nor2  gate2714(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate2715(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate2716(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate2731(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate2732(.a(gate243inter0), .b(s_312), .O(gate243inter1));
  and2  gate2733(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate2734(.a(s_312), .O(gate243inter3));
  inv1  gate2735(.a(s_313), .O(gate243inter4));
  nand2 gate2736(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate2737(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate2738(.a(G245), .O(gate243inter7));
  inv1  gate2739(.a(G733), .O(gate243inter8));
  nand2 gate2740(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate2741(.a(s_313), .b(gate243inter3), .O(gate243inter10));
  nor2  gate2742(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate2743(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate2744(.a(gate243inter12), .b(gate243inter1), .O(G756));

  xor2  gate617(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate618(.a(gate244inter0), .b(s_10), .O(gate244inter1));
  and2  gate619(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate620(.a(s_10), .O(gate244inter3));
  inv1  gate621(.a(s_11), .O(gate244inter4));
  nand2 gate622(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate623(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate624(.a(G721), .O(gate244inter7));
  inv1  gate625(.a(G733), .O(gate244inter8));
  nand2 gate626(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate627(.a(s_11), .b(gate244inter3), .O(gate244inter10));
  nor2  gate628(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate629(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate630(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate1261(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate1262(.a(gate249inter0), .b(s_102), .O(gate249inter1));
  and2  gate1263(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate1264(.a(s_102), .O(gate249inter3));
  inv1  gate1265(.a(s_103), .O(gate249inter4));
  nand2 gate1266(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate1267(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate1268(.a(G254), .O(gate249inter7));
  inv1  gate1269(.a(G742), .O(gate249inter8));
  nand2 gate1270(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate1271(.a(s_103), .b(gate249inter3), .O(gate249inter10));
  nor2  gate1272(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate1273(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate1274(.a(gate249inter12), .b(gate249inter1), .O(G762));

  xor2  gate1065(.a(G742), .b(G706), .O(gate250inter0));
  nand2 gate1066(.a(gate250inter0), .b(s_74), .O(gate250inter1));
  and2  gate1067(.a(G742), .b(G706), .O(gate250inter2));
  inv1  gate1068(.a(s_74), .O(gate250inter3));
  inv1  gate1069(.a(s_75), .O(gate250inter4));
  nand2 gate1070(.a(gate250inter4), .b(gate250inter3), .O(gate250inter5));
  nor2  gate1071(.a(gate250inter5), .b(gate250inter2), .O(gate250inter6));
  inv1  gate1072(.a(G706), .O(gate250inter7));
  inv1  gate1073(.a(G742), .O(gate250inter8));
  nand2 gate1074(.a(gate250inter8), .b(gate250inter7), .O(gate250inter9));
  nand2 gate1075(.a(s_75), .b(gate250inter3), .O(gate250inter10));
  nor2  gate1076(.a(gate250inter10), .b(gate250inter9), .O(gate250inter11));
  nor2  gate1077(.a(gate250inter11), .b(gate250inter6), .O(gate250inter12));
  nand2 gate1078(.a(gate250inter12), .b(gate250inter1), .O(G763));
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate2563(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate2564(.a(gate252inter0), .b(s_288), .O(gate252inter1));
  and2  gate2565(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate2566(.a(s_288), .O(gate252inter3));
  inv1  gate2567(.a(s_289), .O(gate252inter4));
  nand2 gate2568(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate2569(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate2570(.a(G709), .O(gate252inter7));
  inv1  gate2571(.a(G745), .O(gate252inter8));
  nand2 gate2572(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate2573(.a(s_289), .b(gate252inter3), .O(gate252inter10));
  nor2  gate2574(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate2575(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate2576(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );

  xor2  gate1849(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate1850(.a(gate254inter0), .b(s_186), .O(gate254inter1));
  and2  gate1851(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate1852(.a(s_186), .O(gate254inter3));
  inv1  gate1853(.a(s_187), .O(gate254inter4));
  nand2 gate1854(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate1855(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate1856(.a(G712), .O(gate254inter7));
  inv1  gate1857(.a(G748), .O(gate254inter8));
  nand2 gate1858(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate1859(.a(s_187), .b(gate254inter3), .O(gate254inter10));
  nor2  gate1860(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate1861(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate1862(.a(gate254inter12), .b(gate254inter1), .O(G767));

  xor2  gate2605(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate2606(.a(gate255inter0), .b(s_294), .O(gate255inter1));
  and2  gate2607(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate2608(.a(s_294), .O(gate255inter3));
  inv1  gate2609(.a(s_295), .O(gate255inter4));
  nand2 gate2610(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate2611(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate2612(.a(G263), .O(gate255inter7));
  inv1  gate2613(.a(G751), .O(gate255inter8));
  nand2 gate2614(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate2615(.a(s_295), .b(gate255inter3), .O(gate255inter10));
  nor2  gate2616(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate2617(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate2618(.a(gate255inter12), .b(gate255inter1), .O(G768));

  xor2  gate1345(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate1346(.a(gate256inter0), .b(s_114), .O(gate256inter1));
  and2  gate1347(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate1348(.a(s_114), .O(gate256inter3));
  inv1  gate1349(.a(s_115), .O(gate256inter4));
  nand2 gate1350(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate1351(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate1352(.a(G715), .O(gate256inter7));
  inv1  gate1353(.a(G751), .O(gate256inter8));
  nand2 gate1354(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate1355(.a(s_115), .b(gate256inter3), .O(gate256inter10));
  nor2  gate1356(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate1357(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate1358(.a(gate256inter12), .b(gate256inter1), .O(G769));
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate757(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate758(.a(gate261inter0), .b(s_30), .O(gate261inter1));
  and2  gate759(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate760(.a(s_30), .O(gate261inter3));
  inv1  gate761(.a(s_31), .O(gate261inter4));
  nand2 gate762(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate763(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate764(.a(G762), .O(gate261inter7));
  inv1  gate765(.a(G763), .O(gate261inter8));
  nand2 gate766(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate767(.a(s_31), .b(gate261inter3), .O(gate261inter10));
  nor2  gate768(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate769(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate770(.a(gate261inter12), .b(gate261inter1), .O(G782));
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate1163(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate1164(.a(gate263inter0), .b(s_88), .O(gate263inter1));
  and2  gate1165(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate1166(.a(s_88), .O(gate263inter3));
  inv1  gate1167(.a(s_89), .O(gate263inter4));
  nand2 gate1168(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate1169(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate1170(.a(G766), .O(gate263inter7));
  inv1  gate1171(.a(G767), .O(gate263inter8));
  nand2 gate1172(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate1173(.a(s_89), .b(gate263inter3), .O(gate263inter10));
  nor2  gate1174(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate1175(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate1176(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate1961(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate1962(.a(gate265inter0), .b(s_202), .O(gate265inter1));
  and2  gate1963(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate1964(.a(s_202), .O(gate265inter3));
  inv1  gate1965(.a(s_203), .O(gate265inter4));
  nand2 gate1966(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate1967(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate1968(.a(G642), .O(gate265inter7));
  inv1  gate1969(.a(G770), .O(gate265inter8));
  nand2 gate1970(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate1971(.a(s_203), .b(gate265inter3), .O(gate265inter10));
  nor2  gate1972(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate1973(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate1974(.a(gate265inter12), .b(gate265inter1), .O(G794));
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate2017(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate2018(.a(gate267inter0), .b(s_210), .O(gate267inter1));
  and2  gate2019(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate2020(.a(s_210), .O(gate267inter3));
  inv1  gate2021(.a(s_211), .O(gate267inter4));
  nand2 gate2022(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate2023(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate2024(.a(G648), .O(gate267inter7));
  inv1  gate2025(.a(G776), .O(gate267inter8));
  nand2 gate2026(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate2027(.a(s_211), .b(gate267inter3), .O(gate267inter10));
  nor2  gate2028(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate2029(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate2030(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate575(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate576(.a(gate271inter0), .b(s_4), .O(gate271inter1));
  and2  gate577(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate578(.a(s_4), .O(gate271inter3));
  inv1  gate579(.a(s_5), .O(gate271inter4));
  nand2 gate580(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate581(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate582(.a(G660), .O(gate271inter7));
  inv1  gate583(.a(G788), .O(gate271inter8));
  nand2 gate584(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate585(.a(s_5), .b(gate271inter3), .O(gate271inter10));
  nor2  gate586(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate587(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate588(.a(gate271inter12), .b(gate271inter1), .O(G812));

  xor2  gate2549(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate2550(.a(gate272inter0), .b(s_286), .O(gate272inter1));
  and2  gate2551(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate2552(.a(s_286), .O(gate272inter3));
  inv1  gate2553(.a(s_287), .O(gate272inter4));
  nand2 gate2554(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate2555(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate2556(.a(G663), .O(gate272inter7));
  inv1  gate2557(.a(G791), .O(gate272inter8));
  nand2 gate2558(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate2559(.a(s_287), .b(gate272inter3), .O(gate272inter10));
  nor2  gate2560(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate2561(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate2562(.a(gate272inter12), .b(gate272inter1), .O(G815));

  xor2  gate1107(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate1108(.a(gate273inter0), .b(s_80), .O(gate273inter1));
  and2  gate1109(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate1110(.a(s_80), .O(gate273inter3));
  inv1  gate1111(.a(s_81), .O(gate273inter4));
  nand2 gate1112(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate1113(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate1114(.a(G642), .O(gate273inter7));
  inv1  gate1115(.a(G794), .O(gate273inter8));
  nand2 gate1116(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate1117(.a(s_81), .b(gate273inter3), .O(gate273inter10));
  nor2  gate1118(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate1119(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate1120(.a(gate273inter12), .b(gate273inter1), .O(G818));
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate1891(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate1892(.a(gate280inter0), .b(s_192), .O(gate280inter1));
  and2  gate1893(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate1894(.a(s_192), .O(gate280inter3));
  inv1  gate1895(.a(s_193), .O(gate280inter4));
  nand2 gate1896(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate1897(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate1898(.a(G779), .O(gate280inter7));
  inv1  gate1899(.a(G803), .O(gate280inter8));
  nand2 gate1900(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate1901(.a(s_193), .b(gate280inter3), .O(gate280inter10));
  nor2  gate1902(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate1903(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate1904(.a(gate280inter12), .b(gate280inter1), .O(G825));
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate2241(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate2242(.a(gate282inter0), .b(s_242), .O(gate282inter1));
  and2  gate2243(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate2244(.a(s_242), .O(gate282inter3));
  inv1  gate2245(.a(s_243), .O(gate282inter4));
  nand2 gate2246(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate2247(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate2248(.a(G782), .O(gate282inter7));
  inv1  gate2249(.a(G806), .O(gate282inter8));
  nand2 gate2250(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate2251(.a(s_243), .b(gate282inter3), .O(gate282inter10));
  nor2  gate2252(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate2253(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate2254(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );

  xor2  gate2577(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate2578(.a(gate284inter0), .b(s_290), .O(gate284inter1));
  and2  gate2579(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate2580(.a(s_290), .O(gate284inter3));
  inv1  gate2581(.a(s_291), .O(gate284inter4));
  nand2 gate2582(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate2583(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate2584(.a(G785), .O(gate284inter7));
  inv1  gate2585(.a(G809), .O(gate284inter8));
  nand2 gate2586(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate2587(.a(s_291), .b(gate284inter3), .O(gate284inter10));
  nor2  gate2588(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate2589(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate2590(.a(gate284inter12), .b(gate284inter1), .O(G829));

  xor2  gate2115(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate2116(.a(gate285inter0), .b(s_224), .O(gate285inter1));
  and2  gate2117(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate2118(.a(s_224), .O(gate285inter3));
  inv1  gate2119(.a(s_225), .O(gate285inter4));
  nand2 gate2120(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate2121(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate2122(.a(G660), .O(gate285inter7));
  inv1  gate2123(.a(G812), .O(gate285inter8));
  nand2 gate2124(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate2125(.a(s_225), .b(gate285inter3), .O(gate285inter10));
  nor2  gate2126(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate2127(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate2128(.a(gate285inter12), .b(gate285inter1), .O(G830));

  xor2  gate2493(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate2494(.a(gate286inter0), .b(s_278), .O(gate286inter1));
  and2  gate2495(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate2496(.a(s_278), .O(gate286inter3));
  inv1  gate2497(.a(s_279), .O(gate286inter4));
  nand2 gate2498(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate2499(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate2500(.a(G788), .O(gate286inter7));
  inv1  gate2501(.a(G812), .O(gate286inter8));
  nand2 gate2502(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate2503(.a(s_279), .b(gate286inter3), .O(gate286inter10));
  nor2  gate2504(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate2505(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate2506(.a(gate286inter12), .b(gate286inter1), .O(G831));

  xor2  gate1471(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate1472(.a(gate287inter0), .b(s_132), .O(gate287inter1));
  and2  gate1473(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate1474(.a(s_132), .O(gate287inter3));
  inv1  gate1475(.a(s_133), .O(gate287inter4));
  nand2 gate1476(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate1477(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate1478(.a(G663), .O(gate287inter7));
  inv1  gate1479(.a(G815), .O(gate287inter8));
  nand2 gate1480(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate1481(.a(s_133), .b(gate287inter3), .O(gate287inter10));
  nor2  gate1482(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate1483(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate1484(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate2101(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate2102(.a(gate292inter0), .b(s_222), .O(gate292inter1));
  and2  gate2103(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate2104(.a(s_222), .O(gate292inter3));
  inv1  gate2105(.a(s_223), .O(gate292inter4));
  nand2 gate2106(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate2107(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate2108(.a(G824), .O(gate292inter7));
  inv1  gate2109(.a(G825), .O(gate292inter8));
  nand2 gate2110(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate2111(.a(s_223), .b(gate292inter3), .O(gate292inter10));
  nor2  gate2112(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate2113(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate2114(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate2829(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate2830(.a(gate295inter0), .b(s_326), .O(gate295inter1));
  and2  gate2831(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate2832(.a(s_326), .O(gate295inter3));
  inv1  gate2833(.a(s_327), .O(gate295inter4));
  nand2 gate2834(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate2835(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate2836(.a(G830), .O(gate295inter7));
  inv1  gate2837(.a(G831), .O(gate295inter8));
  nand2 gate2838(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate2839(.a(s_327), .b(gate295inter3), .O(gate295inter10));
  nor2  gate2840(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate2841(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate2842(.a(gate295inter12), .b(gate295inter1), .O(G912));
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate1317(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate1318(.a(gate387inter0), .b(s_110), .O(gate387inter1));
  and2  gate1319(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate1320(.a(s_110), .O(gate387inter3));
  inv1  gate1321(.a(s_111), .O(gate387inter4));
  nand2 gate1322(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate1323(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate1324(.a(G1), .O(gate387inter7));
  inv1  gate1325(.a(G1036), .O(gate387inter8));
  nand2 gate1326(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate1327(.a(s_111), .b(gate387inter3), .O(gate387inter10));
  nor2  gate1328(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate1329(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate1330(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );

  xor2  gate1807(.a(G1042), .b(G3), .O(gate389inter0));
  nand2 gate1808(.a(gate389inter0), .b(s_180), .O(gate389inter1));
  and2  gate1809(.a(G1042), .b(G3), .O(gate389inter2));
  inv1  gate1810(.a(s_180), .O(gate389inter3));
  inv1  gate1811(.a(s_181), .O(gate389inter4));
  nand2 gate1812(.a(gate389inter4), .b(gate389inter3), .O(gate389inter5));
  nor2  gate1813(.a(gate389inter5), .b(gate389inter2), .O(gate389inter6));
  inv1  gate1814(.a(G3), .O(gate389inter7));
  inv1  gate1815(.a(G1042), .O(gate389inter8));
  nand2 gate1816(.a(gate389inter8), .b(gate389inter7), .O(gate389inter9));
  nand2 gate1817(.a(s_181), .b(gate389inter3), .O(gate389inter10));
  nor2  gate1818(.a(gate389inter10), .b(gate389inter9), .O(gate389inter11));
  nor2  gate1819(.a(gate389inter11), .b(gate389inter6), .O(gate389inter12));
  nand2 gate1820(.a(gate389inter12), .b(gate389inter1), .O(G1138));
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate1191(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate1192(.a(gate391inter0), .b(s_92), .O(gate391inter1));
  and2  gate1193(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate1194(.a(s_92), .O(gate391inter3));
  inv1  gate1195(.a(s_93), .O(gate391inter4));
  nand2 gate1196(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate1197(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate1198(.a(G5), .O(gate391inter7));
  inv1  gate1199(.a(G1048), .O(gate391inter8));
  nand2 gate1200(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate1201(.a(s_93), .b(gate391inter3), .O(gate391inter10));
  nor2  gate1202(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate1203(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate1204(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );

  xor2  gate1975(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate1976(.a(gate399inter0), .b(s_204), .O(gate399inter1));
  and2  gate1977(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate1978(.a(s_204), .O(gate399inter3));
  inv1  gate1979(.a(s_205), .O(gate399inter4));
  nand2 gate1980(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate1981(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate1982(.a(G13), .O(gate399inter7));
  inv1  gate1983(.a(G1072), .O(gate399inter8));
  nand2 gate1984(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate1985(.a(s_205), .b(gate399inter3), .O(gate399inter10));
  nor2  gate1986(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate1987(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate1988(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );

  xor2  gate2381(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate2382(.a(gate404inter0), .b(s_262), .O(gate404inter1));
  and2  gate2383(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate2384(.a(s_262), .O(gate404inter3));
  inv1  gate2385(.a(s_263), .O(gate404inter4));
  nand2 gate2386(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate2387(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate2388(.a(G18), .O(gate404inter7));
  inv1  gate2389(.a(G1087), .O(gate404inter8));
  nand2 gate2390(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate2391(.a(s_263), .b(gate404inter3), .O(gate404inter10));
  nor2  gate2392(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate2393(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate2394(.a(gate404inter12), .b(gate404inter1), .O(G1183));

  xor2  gate883(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate884(.a(gate405inter0), .b(s_48), .O(gate405inter1));
  and2  gate885(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate886(.a(s_48), .O(gate405inter3));
  inv1  gate887(.a(s_49), .O(gate405inter4));
  nand2 gate888(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate889(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate890(.a(G19), .O(gate405inter7));
  inv1  gate891(.a(G1090), .O(gate405inter8));
  nand2 gate892(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate893(.a(s_49), .b(gate405inter3), .O(gate405inter10));
  nor2  gate894(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate895(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate896(.a(gate405inter12), .b(gate405inter1), .O(G1186));
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate1555(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate1556(.a(gate407inter0), .b(s_144), .O(gate407inter1));
  and2  gate1557(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate1558(.a(s_144), .O(gate407inter3));
  inv1  gate1559(.a(s_145), .O(gate407inter4));
  nand2 gate1560(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate1561(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate1562(.a(G21), .O(gate407inter7));
  inv1  gate1563(.a(G1096), .O(gate407inter8));
  nand2 gate1564(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate1565(.a(s_145), .b(gate407inter3), .O(gate407inter10));
  nor2  gate1566(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate1567(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate1568(.a(gate407inter12), .b(gate407inter1), .O(G1192));
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate1513(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate1514(.a(gate413inter0), .b(s_138), .O(gate413inter1));
  and2  gate1515(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate1516(.a(s_138), .O(gate413inter3));
  inv1  gate1517(.a(s_139), .O(gate413inter4));
  nand2 gate1518(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate1519(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate1520(.a(G27), .O(gate413inter7));
  inv1  gate1521(.a(G1114), .O(gate413inter8));
  nand2 gate1522(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate1523(.a(s_139), .b(gate413inter3), .O(gate413inter10));
  nor2  gate1524(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate1525(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate1526(.a(gate413inter12), .b(gate413inter1), .O(G1210));

  xor2  gate2213(.a(G1117), .b(G28), .O(gate414inter0));
  nand2 gate2214(.a(gate414inter0), .b(s_238), .O(gate414inter1));
  and2  gate2215(.a(G1117), .b(G28), .O(gate414inter2));
  inv1  gate2216(.a(s_238), .O(gate414inter3));
  inv1  gate2217(.a(s_239), .O(gate414inter4));
  nand2 gate2218(.a(gate414inter4), .b(gate414inter3), .O(gate414inter5));
  nor2  gate2219(.a(gate414inter5), .b(gate414inter2), .O(gate414inter6));
  inv1  gate2220(.a(G28), .O(gate414inter7));
  inv1  gate2221(.a(G1117), .O(gate414inter8));
  nand2 gate2222(.a(gate414inter8), .b(gate414inter7), .O(gate414inter9));
  nand2 gate2223(.a(s_239), .b(gate414inter3), .O(gate414inter10));
  nor2  gate2224(.a(gate414inter10), .b(gate414inter9), .O(gate414inter11));
  nor2  gate2225(.a(gate414inter11), .b(gate414inter6), .O(gate414inter12));
  nand2 gate2226(.a(gate414inter12), .b(gate414inter1), .O(G1213));

  xor2  gate1079(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate1080(.a(gate415inter0), .b(s_76), .O(gate415inter1));
  and2  gate1081(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate1082(.a(s_76), .O(gate415inter3));
  inv1  gate1083(.a(s_77), .O(gate415inter4));
  nand2 gate1084(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate1085(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate1086(.a(G29), .O(gate415inter7));
  inv1  gate1087(.a(G1120), .O(gate415inter8));
  nand2 gate1088(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate1089(.a(s_77), .b(gate415inter3), .O(gate415inter10));
  nor2  gate1090(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate1091(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate1092(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );

  xor2  gate2689(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate2690(.a(gate421inter0), .b(s_306), .O(gate421inter1));
  and2  gate2691(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate2692(.a(s_306), .O(gate421inter3));
  inv1  gate2693(.a(s_307), .O(gate421inter4));
  nand2 gate2694(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate2695(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate2696(.a(G2), .O(gate421inter7));
  inv1  gate2697(.a(G1135), .O(gate421inter8));
  nand2 gate2698(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate2699(.a(s_307), .b(gate421inter3), .O(gate421inter10));
  nor2  gate2700(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate2701(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate2702(.a(gate421inter12), .b(gate421inter1), .O(G1230));

  xor2  gate2843(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate2844(.a(gate422inter0), .b(s_328), .O(gate422inter1));
  and2  gate2845(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate2846(.a(s_328), .O(gate422inter3));
  inv1  gate2847(.a(s_329), .O(gate422inter4));
  nand2 gate2848(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate2849(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate2850(.a(G1039), .O(gate422inter7));
  inv1  gate2851(.a(G1135), .O(gate422inter8));
  nand2 gate2852(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate2853(.a(s_329), .b(gate422inter3), .O(gate422inter10));
  nor2  gate2854(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate2855(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate2856(.a(gate422inter12), .b(gate422inter1), .O(G1231));

  xor2  gate2073(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate2074(.a(gate423inter0), .b(s_218), .O(gate423inter1));
  and2  gate2075(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate2076(.a(s_218), .O(gate423inter3));
  inv1  gate2077(.a(s_219), .O(gate423inter4));
  nand2 gate2078(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate2079(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate2080(.a(G3), .O(gate423inter7));
  inv1  gate2081(.a(G1138), .O(gate423inter8));
  nand2 gate2082(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate2083(.a(s_219), .b(gate423inter3), .O(gate423inter10));
  nor2  gate2084(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate2085(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate2086(.a(gate423inter12), .b(gate423inter1), .O(G1232));
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate1177(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate1178(.a(gate425inter0), .b(s_90), .O(gate425inter1));
  and2  gate1179(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate1180(.a(s_90), .O(gate425inter3));
  inv1  gate1181(.a(s_91), .O(gate425inter4));
  nand2 gate1182(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1183(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1184(.a(G4), .O(gate425inter7));
  inv1  gate1185(.a(G1141), .O(gate425inter8));
  nand2 gate1186(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1187(.a(s_91), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1188(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1189(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1190(.a(gate425inter12), .b(gate425inter1), .O(G1234));

  xor2  gate925(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate926(.a(gate426inter0), .b(s_54), .O(gate426inter1));
  and2  gate927(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate928(.a(s_54), .O(gate426inter3));
  inv1  gate929(.a(s_55), .O(gate426inter4));
  nand2 gate930(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate931(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate932(.a(G1045), .O(gate426inter7));
  inv1  gate933(.a(G1141), .O(gate426inter8));
  nand2 gate934(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate935(.a(s_55), .b(gate426inter3), .O(gate426inter10));
  nor2  gate936(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate937(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate938(.a(gate426inter12), .b(gate426inter1), .O(G1235));

  xor2  gate1779(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate1780(.a(gate427inter0), .b(s_176), .O(gate427inter1));
  and2  gate1781(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate1782(.a(s_176), .O(gate427inter3));
  inv1  gate1783(.a(s_177), .O(gate427inter4));
  nand2 gate1784(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate1785(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate1786(.a(G5), .O(gate427inter7));
  inv1  gate1787(.a(G1144), .O(gate427inter8));
  nand2 gate1788(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate1789(.a(s_177), .b(gate427inter3), .O(gate427inter10));
  nor2  gate1790(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate1791(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate1792(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );

  xor2  gate2633(.a(G1153), .b(G1057), .O(gate434inter0));
  nand2 gate2634(.a(gate434inter0), .b(s_298), .O(gate434inter1));
  and2  gate2635(.a(G1153), .b(G1057), .O(gate434inter2));
  inv1  gate2636(.a(s_298), .O(gate434inter3));
  inv1  gate2637(.a(s_299), .O(gate434inter4));
  nand2 gate2638(.a(gate434inter4), .b(gate434inter3), .O(gate434inter5));
  nor2  gate2639(.a(gate434inter5), .b(gate434inter2), .O(gate434inter6));
  inv1  gate2640(.a(G1057), .O(gate434inter7));
  inv1  gate2641(.a(G1153), .O(gate434inter8));
  nand2 gate2642(.a(gate434inter8), .b(gate434inter7), .O(gate434inter9));
  nand2 gate2643(.a(s_299), .b(gate434inter3), .O(gate434inter10));
  nor2  gate2644(.a(gate434inter10), .b(gate434inter9), .O(gate434inter11));
  nor2  gate2645(.a(gate434inter11), .b(gate434inter6), .O(gate434inter12));
  nand2 gate2646(.a(gate434inter12), .b(gate434inter1), .O(G1243));

  xor2  gate1093(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate1094(.a(gate435inter0), .b(s_78), .O(gate435inter1));
  and2  gate1095(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate1096(.a(s_78), .O(gate435inter3));
  inv1  gate1097(.a(s_79), .O(gate435inter4));
  nand2 gate1098(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate1099(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate1100(.a(G9), .O(gate435inter7));
  inv1  gate1101(.a(G1156), .O(gate435inter8));
  nand2 gate1102(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate1103(.a(s_79), .b(gate435inter3), .O(gate435inter10));
  nor2  gate1104(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate1105(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate1106(.a(gate435inter12), .b(gate435inter1), .O(G1244));

  xor2  gate2311(.a(G1156), .b(G1060), .O(gate436inter0));
  nand2 gate2312(.a(gate436inter0), .b(s_252), .O(gate436inter1));
  and2  gate2313(.a(G1156), .b(G1060), .O(gate436inter2));
  inv1  gate2314(.a(s_252), .O(gate436inter3));
  inv1  gate2315(.a(s_253), .O(gate436inter4));
  nand2 gate2316(.a(gate436inter4), .b(gate436inter3), .O(gate436inter5));
  nor2  gate2317(.a(gate436inter5), .b(gate436inter2), .O(gate436inter6));
  inv1  gate2318(.a(G1060), .O(gate436inter7));
  inv1  gate2319(.a(G1156), .O(gate436inter8));
  nand2 gate2320(.a(gate436inter8), .b(gate436inter7), .O(gate436inter9));
  nand2 gate2321(.a(s_253), .b(gate436inter3), .O(gate436inter10));
  nor2  gate2322(.a(gate436inter10), .b(gate436inter9), .O(gate436inter11));
  nor2  gate2323(.a(gate436inter11), .b(gate436inter6), .O(gate436inter12));
  nand2 gate2324(.a(gate436inter12), .b(gate436inter1), .O(G1245));

  xor2  gate2479(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate2480(.a(gate437inter0), .b(s_276), .O(gate437inter1));
  and2  gate2481(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate2482(.a(s_276), .O(gate437inter3));
  inv1  gate2483(.a(s_277), .O(gate437inter4));
  nand2 gate2484(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate2485(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate2486(.a(G10), .O(gate437inter7));
  inv1  gate2487(.a(G1159), .O(gate437inter8));
  nand2 gate2488(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate2489(.a(s_277), .b(gate437inter3), .O(gate437inter10));
  nor2  gate2490(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate2491(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate2492(.a(gate437inter12), .b(gate437inter1), .O(G1246));

  xor2  gate2409(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate2410(.a(gate438inter0), .b(s_266), .O(gate438inter1));
  and2  gate2411(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate2412(.a(s_266), .O(gate438inter3));
  inv1  gate2413(.a(s_267), .O(gate438inter4));
  nand2 gate2414(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate2415(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate2416(.a(G1063), .O(gate438inter7));
  inv1  gate2417(.a(G1159), .O(gate438inter8));
  nand2 gate2418(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate2419(.a(s_267), .b(gate438inter3), .O(gate438inter10));
  nor2  gate2420(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate2421(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate2422(.a(gate438inter12), .b(gate438inter1), .O(G1247));
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate2353(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate2354(.a(gate441inter0), .b(s_258), .O(gate441inter1));
  and2  gate2355(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate2356(.a(s_258), .O(gate441inter3));
  inv1  gate2357(.a(s_259), .O(gate441inter4));
  nand2 gate2358(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate2359(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate2360(.a(G12), .O(gate441inter7));
  inv1  gate2361(.a(G1165), .O(gate441inter8));
  nand2 gate2362(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate2363(.a(s_259), .b(gate441inter3), .O(gate441inter10));
  nor2  gate2364(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate2365(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate2366(.a(gate441inter12), .b(gate441inter1), .O(G1250));
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );

  xor2  gate953(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate954(.a(gate443inter0), .b(s_58), .O(gate443inter1));
  and2  gate955(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate956(.a(s_58), .O(gate443inter3));
  inv1  gate957(.a(s_59), .O(gate443inter4));
  nand2 gate958(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate959(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate960(.a(G13), .O(gate443inter7));
  inv1  gate961(.a(G1168), .O(gate443inter8));
  nand2 gate962(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate963(.a(s_59), .b(gate443inter3), .O(gate443inter10));
  nor2  gate964(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate965(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate966(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );

  xor2  gate1051(.a(G1171), .b(G14), .O(gate445inter0));
  nand2 gate1052(.a(gate445inter0), .b(s_72), .O(gate445inter1));
  and2  gate1053(.a(G1171), .b(G14), .O(gate445inter2));
  inv1  gate1054(.a(s_72), .O(gate445inter3));
  inv1  gate1055(.a(s_73), .O(gate445inter4));
  nand2 gate1056(.a(gate445inter4), .b(gate445inter3), .O(gate445inter5));
  nor2  gate1057(.a(gate445inter5), .b(gate445inter2), .O(gate445inter6));
  inv1  gate1058(.a(G14), .O(gate445inter7));
  inv1  gate1059(.a(G1171), .O(gate445inter8));
  nand2 gate1060(.a(gate445inter8), .b(gate445inter7), .O(gate445inter9));
  nand2 gate1061(.a(s_73), .b(gate445inter3), .O(gate445inter10));
  nor2  gate1062(.a(gate445inter10), .b(gate445inter9), .O(gate445inter11));
  nor2  gate1063(.a(gate445inter11), .b(gate445inter6), .O(gate445inter12));
  nand2 gate1064(.a(gate445inter12), .b(gate445inter1), .O(G1254));

  xor2  gate1877(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate1878(.a(gate446inter0), .b(s_190), .O(gate446inter1));
  and2  gate1879(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate1880(.a(s_190), .O(gate446inter3));
  inv1  gate1881(.a(s_191), .O(gate446inter4));
  nand2 gate1882(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate1883(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate1884(.a(G1075), .O(gate446inter7));
  inv1  gate1885(.a(G1171), .O(gate446inter8));
  nand2 gate1886(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate1887(.a(s_191), .b(gate446inter3), .O(gate446inter10));
  nor2  gate1888(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate1889(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate1890(.a(gate446inter12), .b(gate446inter1), .O(G1255));
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate2367(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate2368(.a(gate448inter0), .b(s_260), .O(gate448inter1));
  and2  gate2369(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate2370(.a(s_260), .O(gate448inter3));
  inv1  gate2371(.a(s_261), .O(gate448inter4));
  nand2 gate2372(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate2373(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate2374(.a(G1078), .O(gate448inter7));
  inv1  gate2375(.a(G1174), .O(gate448inter8));
  nand2 gate2376(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate2377(.a(s_261), .b(gate448inter3), .O(gate448inter10));
  nor2  gate2378(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate2379(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate2380(.a(gate448inter12), .b(gate448inter1), .O(G1257));

  xor2  gate2647(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate2648(.a(gate449inter0), .b(s_300), .O(gate449inter1));
  and2  gate2649(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate2650(.a(s_300), .O(gate449inter3));
  inv1  gate2651(.a(s_301), .O(gate449inter4));
  nand2 gate2652(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate2653(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate2654(.a(G16), .O(gate449inter7));
  inv1  gate2655(.a(G1177), .O(gate449inter8));
  nand2 gate2656(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate2657(.a(s_301), .b(gate449inter3), .O(gate449inter10));
  nor2  gate2658(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate2659(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate2660(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );

  xor2  gate631(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate632(.a(gate451inter0), .b(s_12), .O(gate451inter1));
  and2  gate633(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate634(.a(s_12), .O(gate451inter3));
  inv1  gate635(.a(s_13), .O(gate451inter4));
  nand2 gate636(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate637(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate638(.a(G17), .O(gate451inter7));
  inv1  gate639(.a(G1180), .O(gate451inter8));
  nand2 gate640(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate641(.a(s_13), .b(gate451inter3), .O(gate451inter10));
  nor2  gate642(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate643(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate644(.a(gate451inter12), .b(gate451inter1), .O(G1260));
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate589(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate590(.a(gate453inter0), .b(s_6), .O(gate453inter1));
  and2  gate591(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate592(.a(s_6), .O(gate453inter3));
  inv1  gate593(.a(s_7), .O(gate453inter4));
  nand2 gate594(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate595(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate596(.a(G18), .O(gate453inter7));
  inv1  gate597(.a(G1183), .O(gate453inter8));
  nand2 gate598(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate599(.a(s_7), .b(gate453inter3), .O(gate453inter10));
  nor2  gate600(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate601(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate602(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );

  xor2  gate1233(.a(G1186), .b(G1090), .O(gate456inter0));
  nand2 gate1234(.a(gate456inter0), .b(s_98), .O(gate456inter1));
  and2  gate1235(.a(G1186), .b(G1090), .O(gate456inter2));
  inv1  gate1236(.a(s_98), .O(gate456inter3));
  inv1  gate1237(.a(s_99), .O(gate456inter4));
  nand2 gate1238(.a(gate456inter4), .b(gate456inter3), .O(gate456inter5));
  nor2  gate1239(.a(gate456inter5), .b(gate456inter2), .O(gate456inter6));
  inv1  gate1240(.a(G1090), .O(gate456inter7));
  inv1  gate1241(.a(G1186), .O(gate456inter8));
  nand2 gate1242(.a(gate456inter8), .b(gate456inter7), .O(gate456inter9));
  nand2 gate1243(.a(s_99), .b(gate456inter3), .O(gate456inter10));
  nor2  gate1244(.a(gate456inter10), .b(gate456inter9), .O(gate456inter11));
  nor2  gate1245(.a(gate456inter11), .b(gate456inter6), .O(gate456inter12));
  nand2 gate1246(.a(gate456inter12), .b(gate456inter1), .O(G1265));

  xor2  gate1765(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate1766(.a(gate457inter0), .b(s_174), .O(gate457inter1));
  and2  gate1767(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate1768(.a(s_174), .O(gate457inter3));
  inv1  gate1769(.a(s_175), .O(gate457inter4));
  nand2 gate1770(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate1771(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate1772(.a(G20), .O(gate457inter7));
  inv1  gate1773(.a(G1189), .O(gate457inter8));
  nand2 gate1774(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate1775(.a(s_175), .b(gate457inter3), .O(gate457inter10));
  nor2  gate1776(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate1777(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate1778(.a(gate457inter12), .b(gate457inter1), .O(G1266));

  xor2  gate1863(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate1864(.a(gate458inter0), .b(s_188), .O(gate458inter1));
  and2  gate1865(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate1866(.a(s_188), .O(gate458inter3));
  inv1  gate1867(.a(s_189), .O(gate458inter4));
  nand2 gate1868(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate1869(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate1870(.a(G1093), .O(gate458inter7));
  inv1  gate1871(.a(G1189), .O(gate458inter8));
  nand2 gate1872(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate1873(.a(s_189), .b(gate458inter3), .O(gate458inter10));
  nor2  gate1874(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate1875(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate1876(.a(gate458inter12), .b(gate458inter1), .O(G1267));

  xor2  gate547(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate548(.a(gate459inter0), .b(s_0), .O(gate459inter1));
  and2  gate549(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate550(.a(s_0), .O(gate459inter3));
  inv1  gate551(.a(s_1), .O(gate459inter4));
  nand2 gate552(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate553(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate554(.a(G21), .O(gate459inter7));
  inv1  gate555(.a(G1192), .O(gate459inter8));
  nand2 gate556(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate557(.a(s_1), .b(gate459inter3), .O(gate459inter10));
  nor2  gate558(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate559(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate560(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate1835(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate1836(.a(gate461inter0), .b(s_184), .O(gate461inter1));
  and2  gate1837(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate1838(.a(s_184), .O(gate461inter3));
  inv1  gate1839(.a(s_185), .O(gate461inter4));
  nand2 gate1840(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate1841(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate1842(.a(G22), .O(gate461inter7));
  inv1  gate1843(.a(G1195), .O(gate461inter8));
  nand2 gate1844(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate1845(.a(s_185), .b(gate461inter3), .O(gate461inter10));
  nor2  gate1846(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate1847(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate1848(.a(gate461inter12), .b(gate461inter1), .O(G1270));

  xor2  gate2087(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate2088(.a(gate462inter0), .b(s_220), .O(gate462inter1));
  and2  gate2089(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate2090(.a(s_220), .O(gate462inter3));
  inv1  gate2091(.a(s_221), .O(gate462inter4));
  nand2 gate2092(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate2093(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate2094(.a(G1099), .O(gate462inter7));
  inv1  gate2095(.a(G1195), .O(gate462inter8));
  nand2 gate2096(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate2097(.a(s_221), .b(gate462inter3), .O(gate462inter10));
  nor2  gate2098(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate2099(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate2100(.a(gate462inter12), .b(gate462inter1), .O(G1271));

  xor2  gate743(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate744(.a(gate463inter0), .b(s_28), .O(gate463inter1));
  and2  gate745(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate746(.a(s_28), .O(gate463inter3));
  inv1  gate747(.a(s_29), .O(gate463inter4));
  nand2 gate748(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate749(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate750(.a(G23), .O(gate463inter7));
  inv1  gate751(.a(G1198), .O(gate463inter8));
  nand2 gate752(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate753(.a(s_29), .b(gate463inter3), .O(gate463inter10));
  nor2  gate754(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate755(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate756(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate1037(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate1038(.a(gate465inter0), .b(s_70), .O(gate465inter1));
  and2  gate1039(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate1040(.a(s_70), .O(gate465inter3));
  inv1  gate1041(.a(s_71), .O(gate465inter4));
  nand2 gate1042(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate1043(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate1044(.a(G24), .O(gate465inter7));
  inv1  gate1045(.a(G1201), .O(gate465inter8));
  nand2 gate1046(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate1047(.a(s_71), .b(gate465inter3), .O(gate465inter10));
  nor2  gate1048(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate1049(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate1050(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );

  xor2  gate1485(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate1486(.a(gate468inter0), .b(s_134), .O(gate468inter1));
  and2  gate1487(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate1488(.a(s_134), .O(gate468inter3));
  inv1  gate1489(.a(s_135), .O(gate468inter4));
  nand2 gate1490(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate1491(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate1492(.a(G1108), .O(gate468inter7));
  inv1  gate1493(.a(G1204), .O(gate468inter8));
  nand2 gate1494(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate1495(.a(s_135), .b(gate468inter3), .O(gate468inter10));
  nor2  gate1496(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate1497(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate1498(.a(gate468inter12), .b(gate468inter1), .O(G1277));

  xor2  gate2801(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate2802(.a(gate469inter0), .b(s_322), .O(gate469inter1));
  and2  gate2803(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate2804(.a(s_322), .O(gate469inter3));
  inv1  gate2805(.a(s_323), .O(gate469inter4));
  nand2 gate2806(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate2807(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate2808(.a(G26), .O(gate469inter7));
  inv1  gate2809(.a(G1207), .O(gate469inter8));
  nand2 gate2810(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate2811(.a(s_323), .b(gate469inter3), .O(gate469inter10));
  nor2  gate2812(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate2813(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate2814(.a(gate469inter12), .b(gate469inter1), .O(G1278));

  xor2  gate1737(.a(G1207), .b(G1111), .O(gate470inter0));
  nand2 gate1738(.a(gate470inter0), .b(s_170), .O(gate470inter1));
  and2  gate1739(.a(G1207), .b(G1111), .O(gate470inter2));
  inv1  gate1740(.a(s_170), .O(gate470inter3));
  inv1  gate1741(.a(s_171), .O(gate470inter4));
  nand2 gate1742(.a(gate470inter4), .b(gate470inter3), .O(gate470inter5));
  nor2  gate1743(.a(gate470inter5), .b(gate470inter2), .O(gate470inter6));
  inv1  gate1744(.a(G1111), .O(gate470inter7));
  inv1  gate1745(.a(G1207), .O(gate470inter8));
  nand2 gate1746(.a(gate470inter8), .b(gate470inter7), .O(gate470inter9));
  nand2 gate1747(.a(s_171), .b(gate470inter3), .O(gate470inter10));
  nor2  gate1748(.a(gate470inter10), .b(gate470inter9), .O(gate470inter11));
  nor2  gate1749(.a(gate470inter11), .b(gate470inter6), .O(gate470inter12));
  nand2 gate1750(.a(gate470inter12), .b(gate470inter1), .O(G1279));

  xor2  gate2787(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate2788(.a(gate471inter0), .b(s_320), .O(gate471inter1));
  and2  gate2789(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate2790(.a(s_320), .O(gate471inter3));
  inv1  gate2791(.a(s_321), .O(gate471inter4));
  nand2 gate2792(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate2793(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate2794(.a(G27), .O(gate471inter7));
  inv1  gate2795(.a(G1210), .O(gate471inter8));
  nand2 gate2796(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate2797(.a(s_321), .b(gate471inter3), .O(gate471inter10));
  nor2  gate2798(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate2799(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate2800(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate1457(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate1458(.a(gate475inter0), .b(s_130), .O(gate475inter1));
  and2  gate1459(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate1460(.a(s_130), .O(gate475inter3));
  inv1  gate1461(.a(s_131), .O(gate475inter4));
  nand2 gate1462(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate1463(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate1464(.a(G29), .O(gate475inter7));
  inv1  gate1465(.a(G1216), .O(gate475inter8));
  nand2 gate1466(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate1467(.a(s_131), .b(gate475inter3), .O(gate475inter10));
  nor2  gate1468(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate1469(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate1470(.a(gate475inter12), .b(gate475inter1), .O(G1284));

  xor2  gate701(.a(G1216), .b(G1120), .O(gate476inter0));
  nand2 gate702(.a(gate476inter0), .b(s_22), .O(gate476inter1));
  and2  gate703(.a(G1216), .b(G1120), .O(gate476inter2));
  inv1  gate704(.a(s_22), .O(gate476inter3));
  inv1  gate705(.a(s_23), .O(gate476inter4));
  nand2 gate706(.a(gate476inter4), .b(gate476inter3), .O(gate476inter5));
  nor2  gate707(.a(gate476inter5), .b(gate476inter2), .O(gate476inter6));
  inv1  gate708(.a(G1120), .O(gate476inter7));
  inv1  gate709(.a(G1216), .O(gate476inter8));
  nand2 gate710(.a(gate476inter8), .b(gate476inter7), .O(gate476inter9));
  nand2 gate711(.a(s_23), .b(gate476inter3), .O(gate476inter10));
  nor2  gate712(.a(gate476inter10), .b(gate476inter9), .O(gate476inter11));
  nor2  gate713(.a(gate476inter11), .b(gate476inter6), .O(gate476inter12));
  nand2 gate714(.a(gate476inter12), .b(gate476inter1), .O(G1285));

  xor2  gate1373(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate1374(.a(gate477inter0), .b(s_118), .O(gate477inter1));
  and2  gate1375(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate1376(.a(s_118), .O(gate477inter3));
  inv1  gate1377(.a(s_119), .O(gate477inter4));
  nand2 gate1378(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate1379(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate1380(.a(G30), .O(gate477inter7));
  inv1  gate1381(.a(G1219), .O(gate477inter8));
  nand2 gate1382(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate1383(.a(s_119), .b(gate477inter3), .O(gate477inter10));
  nor2  gate1384(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate1385(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate1386(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );

  xor2  gate841(.a(G1225), .b(G32), .O(gate481inter0));
  nand2 gate842(.a(gate481inter0), .b(s_42), .O(gate481inter1));
  and2  gate843(.a(G1225), .b(G32), .O(gate481inter2));
  inv1  gate844(.a(s_42), .O(gate481inter3));
  inv1  gate845(.a(s_43), .O(gate481inter4));
  nand2 gate846(.a(gate481inter4), .b(gate481inter3), .O(gate481inter5));
  nor2  gate847(.a(gate481inter5), .b(gate481inter2), .O(gate481inter6));
  inv1  gate848(.a(G32), .O(gate481inter7));
  inv1  gate849(.a(G1225), .O(gate481inter8));
  nand2 gate850(.a(gate481inter8), .b(gate481inter7), .O(gate481inter9));
  nand2 gate851(.a(s_43), .b(gate481inter3), .O(gate481inter10));
  nor2  gate852(.a(gate481inter10), .b(gate481inter9), .O(gate481inter11));
  nor2  gate853(.a(gate481inter11), .b(gate481inter6), .O(gate481inter12));
  nand2 gate854(.a(gate481inter12), .b(gate481inter1), .O(G1290));
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate2129(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate2130(.a(gate485inter0), .b(s_226), .O(gate485inter1));
  and2  gate2131(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate2132(.a(s_226), .O(gate485inter3));
  inv1  gate2133(.a(s_227), .O(gate485inter4));
  nand2 gate2134(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate2135(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate2136(.a(G1232), .O(gate485inter7));
  inv1  gate2137(.a(G1233), .O(gate485inter8));
  nand2 gate2138(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate2139(.a(s_227), .b(gate485inter3), .O(gate485inter10));
  nor2  gate2140(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate2141(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate2142(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate799(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate800(.a(gate487inter0), .b(s_36), .O(gate487inter1));
  and2  gate801(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate802(.a(s_36), .O(gate487inter3));
  inv1  gate803(.a(s_37), .O(gate487inter4));
  nand2 gate804(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate805(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate806(.a(G1236), .O(gate487inter7));
  inv1  gate807(.a(G1237), .O(gate487inter8));
  nand2 gate808(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate809(.a(s_37), .b(gate487inter3), .O(gate487inter10));
  nor2  gate810(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate811(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate812(.a(gate487inter12), .b(gate487inter1), .O(G1296));

  xor2  gate1359(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate1360(.a(gate488inter0), .b(s_116), .O(gate488inter1));
  and2  gate1361(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate1362(.a(s_116), .O(gate488inter3));
  inv1  gate1363(.a(s_117), .O(gate488inter4));
  nand2 gate1364(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate1365(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate1366(.a(G1238), .O(gate488inter7));
  inv1  gate1367(.a(G1239), .O(gate488inter8));
  nand2 gate1368(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate1369(.a(s_117), .b(gate488inter3), .O(gate488inter10));
  nor2  gate1370(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate1371(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate1372(.a(gate488inter12), .b(gate488inter1), .O(G1297));

  xor2  gate1793(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate1794(.a(gate489inter0), .b(s_178), .O(gate489inter1));
  and2  gate1795(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate1796(.a(s_178), .O(gate489inter3));
  inv1  gate1797(.a(s_179), .O(gate489inter4));
  nand2 gate1798(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate1799(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate1800(.a(G1240), .O(gate489inter7));
  inv1  gate1801(.a(G1241), .O(gate489inter8));
  nand2 gate1802(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate1803(.a(s_179), .b(gate489inter3), .O(gate489inter10));
  nor2  gate1804(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate1805(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate1806(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate967(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate968(.a(gate491inter0), .b(s_60), .O(gate491inter1));
  and2  gate969(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate970(.a(s_60), .O(gate491inter3));
  inv1  gate971(.a(s_61), .O(gate491inter4));
  nand2 gate972(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate973(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate974(.a(G1244), .O(gate491inter7));
  inv1  gate975(.a(G1245), .O(gate491inter8));
  nand2 gate976(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate977(.a(s_61), .b(gate491inter3), .O(gate491inter10));
  nor2  gate978(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate979(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate980(.a(gate491inter12), .b(gate491inter1), .O(G1300));

  xor2  gate1303(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate1304(.a(gate492inter0), .b(s_108), .O(gate492inter1));
  and2  gate1305(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate1306(.a(s_108), .O(gate492inter3));
  inv1  gate1307(.a(s_109), .O(gate492inter4));
  nand2 gate1308(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate1309(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate1310(.a(G1246), .O(gate492inter7));
  inv1  gate1311(.a(G1247), .O(gate492inter8));
  nand2 gate1312(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate1313(.a(s_109), .b(gate492inter3), .O(gate492inter10));
  nor2  gate1314(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate1315(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate1316(.a(gate492inter12), .b(gate492inter1), .O(G1301));
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate2227(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate2228(.a(gate496inter0), .b(s_240), .O(gate496inter1));
  and2  gate2229(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate2230(.a(s_240), .O(gate496inter3));
  inv1  gate2231(.a(s_241), .O(gate496inter4));
  nand2 gate2232(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate2233(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate2234(.a(G1254), .O(gate496inter7));
  inv1  gate2235(.a(G1255), .O(gate496inter8));
  nand2 gate2236(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate2237(.a(s_241), .b(gate496inter3), .O(gate496inter10));
  nor2  gate2238(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate2239(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate2240(.a(gate496inter12), .b(gate496inter1), .O(G1305));
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );

  xor2  gate2059(.a(G1269), .b(G1268), .O(gate503inter0));
  nand2 gate2060(.a(gate503inter0), .b(s_216), .O(gate503inter1));
  and2  gate2061(.a(G1269), .b(G1268), .O(gate503inter2));
  inv1  gate2062(.a(s_216), .O(gate503inter3));
  inv1  gate2063(.a(s_217), .O(gate503inter4));
  nand2 gate2064(.a(gate503inter4), .b(gate503inter3), .O(gate503inter5));
  nor2  gate2065(.a(gate503inter5), .b(gate503inter2), .O(gate503inter6));
  inv1  gate2066(.a(G1268), .O(gate503inter7));
  inv1  gate2067(.a(G1269), .O(gate503inter8));
  nand2 gate2068(.a(gate503inter8), .b(gate503inter7), .O(gate503inter9));
  nand2 gate2069(.a(s_217), .b(gate503inter3), .O(gate503inter10));
  nor2  gate2070(.a(gate503inter10), .b(gate503inter9), .O(gate503inter11));
  nor2  gate2071(.a(gate503inter11), .b(gate503inter6), .O(gate503inter12));
  nand2 gate2072(.a(gate503inter12), .b(gate503inter1), .O(G1312));

  xor2  gate995(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate996(.a(gate504inter0), .b(s_64), .O(gate504inter1));
  and2  gate997(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate998(.a(s_64), .O(gate504inter3));
  inv1  gate999(.a(s_65), .O(gate504inter4));
  nand2 gate1000(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate1001(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate1002(.a(G1270), .O(gate504inter7));
  inv1  gate1003(.a(G1271), .O(gate504inter8));
  nand2 gate1004(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate1005(.a(s_65), .b(gate504inter3), .O(gate504inter10));
  nor2  gate1006(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate1007(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate1008(.a(gate504inter12), .b(gate504inter1), .O(G1313));

  xor2  gate1023(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate1024(.a(gate505inter0), .b(s_68), .O(gate505inter1));
  and2  gate1025(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate1026(.a(s_68), .O(gate505inter3));
  inv1  gate1027(.a(s_69), .O(gate505inter4));
  nand2 gate1028(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate1029(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate1030(.a(G1272), .O(gate505inter7));
  inv1  gate1031(.a(G1273), .O(gate505inter8));
  nand2 gate1032(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate1033(.a(s_69), .b(gate505inter3), .O(gate505inter10));
  nor2  gate1034(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate1035(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate1036(.a(gate505inter12), .b(gate505inter1), .O(G1314));
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );

  xor2  gate2157(.a(G1277), .b(G1276), .O(gate507inter0));
  nand2 gate2158(.a(gate507inter0), .b(s_230), .O(gate507inter1));
  and2  gate2159(.a(G1277), .b(G1276), .O(gate507inter2));
  inv1  gate2160(.a(s_230), .O(gate507inter3));
  inv1  gate2161(.a(s_231), .O(gate507inter4));
  nand2 gate2162(.a(gate507inter4), .b(gate507inter3), .O(gate507inter5));
  nor2  gate2163(.a(gate507inter5), .b(gate507inter2), .O(gate507inter6));
  inv1  gate2164(.a(G1276), .O(gate507inter7));
  inv1  gate2165(.a(G1277), .O(gate507inter8));
  nand2 gate2166(.a(gate507inter8), .b(gate507inter7), .O(gate507inter9));
  nand2 gate2167(.a(s_231), .b(gate507inter3), .O(gate507inter10));
  nor2  gate2168(.a(gate507inter10), .b(gate507inter9), .O(gate507inter11));
  nor2  gate2169(.a(gate507inter11), .b(gate507inter6), .O(gate507inter12));
  nand2 gate2170(.a(gate507inter12), .b(gate507inter1), .O(G1316));

  xor2  gate1415(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate1416(.a(gate508inter0), .b(s_124), .O(gate508inter1));
  and2  gate1417(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate1418(.a(s_124), .O(gate508inter3));
  inv1  gate1419(.a(s_125), .O(gate508inter4));
  nand2 gate1420(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate1421(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate1422(.a(G1278), .O(gate508inter7));
  inv1  gate1423(.a(G1279), .O(gate508inter8));
  nand2 gate1424(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate1425(.a(s_125), .b(gate508inter3), .O(gate508inter10));
  nor2  gate1426(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate1427(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate1428(.a(gate508inter12), .b(gate508inter1), .O(G1317));

  xor2  gate2759(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate2760(.a(gate509inter0), .b(s_316), .O(gate509inter1));
  and2  gate2761(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate2762(.a(s_316), .O(gate509inter3));
  inv1  gate2763(.a(s_317), .O(gate509inter4));
  nand2 gate2764(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate2765(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate2766(.a(G1280), .O(gate509inter7));
  inv1  gate2767(.a(G1281), .O(gate509inter8));
  nand2 gate2768(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate2769(.a(s_317), .b(gate509inter3), .O(gate509inter10));
  nor2  gate2770(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate2771(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate2772(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );

  xor2  gate1009(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate1010(.a(gate512inter0), .b(s_66), .O(gate512inter1));
  and2  gate1011(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate1012(.a(s_66), .O(gate512inter3));
  inv1  gate1013(.a(s_67), .O(gate512inter4));
  nand2 gate1014(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate1015(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate1016(.a(G1286), .O(gate512inter7));
  inv1  gate1017(.a(G1287), .O(gate512inter8));
  nand2 gate1018(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate1019(.a(s_67), .b(gate512inter3), .O(gate512inter10));
  nor2  gate1020(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate1021(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate1022(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule