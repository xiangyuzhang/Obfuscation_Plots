module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281, s_282, s_283, s_284, s_285, s_286, s_287, s_288, s_289, s_290, s_291, s_292, s_293, s_294, s_295, s_296, s_297, s_298, s_299, s_300, s_301, s_302, s_303, s_304, s_305, s_306, s_307, s_308, s_309, s_310, s_311, s_312, s_313, s_314, s_315, s_316, s_317, s_318, s_319, s_320, s_321, s_322, s_323, s_324, s_325, s_326, s_327, s_328, s_329, s_330, s_331, s_332, s_333, s_334, s_335, s_336, s_337, s_338, s_339, s_340, s_341, s_342, s_343, s_344, s_345, s_346, s_347, s_348, s_349, s_350, s_351;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate119inter0, gate119inter1, gate119inter2, gate119inter3, gate119inter4, gate119inter5, gate119inter6, gate119inter7, gate119inter8, gate119inter9, gate119inter10, gate119inter11, gate119inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate78inter0, gate78inter1, gate78inter2, gate78inter3, gate78inter4, gate78inter5, gate78inter6, gate78inter7, gate78inter8, gate78inter9, gate78inter10, gate78inter11, gate78inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate416inter0, gate416inter1, gate416inter2, gate416inter3, gate416inter4, gate416inter5, gate416inter6, gate416inter7, gate416inter8, gate416inter9, gate416inter10, gate416inter11, gate416inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate267inter0, gate267inter1, gate267inter2, gate267inter3, gate267inter4, gate267inter5, gate267inter6, gate267inter7, gate267inter8, gate267inter9, gate267inter10, gate267inter11, gate267inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate44inter0, gate44inter1, gate44inter2, gate44inter3, gate44inter4, gate44inter5, gate44inter6, gate44inter7, gate44inter8, gate44inter9, gate44inter10, gate44inter11, gate44inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate132inter0, gate132inter1, gate132inter2, gate132inter3, gate132inter4, gate132inter5, gate132inter6, gate132inter7, gate132inter8, gate132inter9, gate132inter10, gate132inter11, gate132inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate234inter0, gate234inter1, gate234inter2, gate234inter3, gate234inter4, gate234inter5, gate234inter6, gate234inter7, gate234inter8, gate234inter9, gate234inter10, gate234inter11, gate234inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate450inter0, gate450inter1, gate450inter2, gate450inter3, gate450inter4, gate450inter5, gate450inter6, gate450inter7, gate450inter8, gate450inter9, gate450inter10, gate450inter11, gate450inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate469inter0, gate469inter1, gate469inter2, gate469inter3, gate469inter4, gate469inter5, gate469inter6, gate469inter7, gate469inter8, gate469inter9, gate469inter10, gate469inter11, gate469inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate398inter0, gate398inter1, gate398inter2, gate398inter3, gate398inter4, gate398inter5, gate398inter6, gate398inter7, gate398inter8, gate398inter9, gate398inter10, gate398inter11, gate398inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate448inter0, gate448inter1, gate448inter2, gate448inter3, gate448inter4, gate448inter5, gate448inter6, gate448inter7, gate448inter8, gate448inter9, gate448inter10, gate448inter11, gate448inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate239inter0, gate239inter1, gate239inter2, gate239inter3, gate239inter4, gate239inter5, gate239inter6, gate239inter7, gate239inter8, gate239inter9, gate239inter10, gate239inter11, gate239inter12, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate245inter0, gate245inter1, gate245inter2, gate245inter3, gate245inter4, gate245inter5, gate245inter6, gate245inter7, gate245inter8, gate245inter9, gate245inter10, gate245inter11, gate245inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate451inter0, gate451inter1, gate451inter2, gate451inter3, gate451inter4, gate451inter5, gate451inter6, gate451inter7, gate451inter8, gate451inter9, gate451inter10, gate451inter11, gate451inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate96inter0, gate96inter1, gate96inter2, gate96inter3, gate96inter4, gate96inter5, gate96inter6, gate96inter7, gate96inter8, gate96inter9, gate96inter10, gate96inter11, gate96inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate399inter0, gate399inter1, gate399inter2, gate399inter3, gate399inter4, gate399inter5, gate399inter6, gate399inter7, gate399inter8, gate399inter9, gate399inter10, gate399inter11, gate399inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate169inter0, gate169inter1, gate169inter2, gate169inter3, gate169inter4, gate169inter5, gate169inter6, gate169inter7, gate169inter8, gate169inter9, gate169inter10, gate169inter11, gate169inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate112inter0, gate112inter1, gate112inter2, gate112inter3, gate112inter4, gate112inter5, gate112inter6, gate112inter7, gate112inter8, gate112inter9, gate112inter10, gate112inter11, gate112inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate64inter0, gate64inter1, gate64inter2, gate64inter3, gate64inter4, gate64inter5, gate64inter6, gate64inter7, gate64inter8, gate64inter9, gate64inter10, gate64inter11, gate64inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate813(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate814(.a(gate9inter0), .b(s_38), .O(gate9inter1));
  and2  gate815(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate816(.a(s_38), .O(gate9inter3));
  inv1  gate817(.a(s_39), .O(gate9inter4));
  nand2 gate818(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate819(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate820(.a(G1), .O(gate9inter7));
  inv1  gate821(.a(G2), .O(gate9inter8));
  nand2 gate822(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate823(.a(s_39), .b(gate9inter3), .O(gate9inter10));
  nor2  gate824(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate825(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate826(.a(gate9inter12), .b(gate9inter1), .O(G266));

  xor2  gate687(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate688(.a(gate10inter0), .b(s_20), .O(gate10inter1));
  and2  gate689(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate690(.a(s_20), .O(gate10inter3));
  inv1  gate691(.a(s_21), .O(gate10inter4));
  nand2 gate692(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate693(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate694(.a(G3), .O(gate10inter7));
  inv1  gate695(.a(G4), .O(gate10inter8));
  nand2 gate696(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate697(.a(s_21), .b(gate10inter3), .O(gate10inter10));
  nor2  gate698(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate699(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate700(.a(gate10inter12), .b(gate10inter1), .O(G269));

  xor2  gate2395(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate2396(.a(gate11inter0), .b(s_264), .O(gate11inter1));
  and2  gate2397(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate2398(.a(s_264), .O(gate11inter3));
  inv1  gate2399(.a(s_265), .O(gate11inter4));
  nand2 gate2400(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate2401(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate2402(.a(G5), .O(gate11inter7));
  inv1  gate2403(.a(G6), .O(gate11inter8));
  nand2 gate2404(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate2405(.a(s_265), .b(gate11inter3), .O(gate11inter10));
  nor2  gate2406(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate2407(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate2408(.a(gate11inter12), .b(gate11inter1), .O(G272));

  xor2  gate2269(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate2270(.a(gate12inter0), .b(s_246), .O(gate12inter1));
  and2  gate2271(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate2272(.a(s_246), .O(gate12inter3));
  inv1  gate2273(.a(s_247), .O(gate12inter4));
  nand2 gate2274(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate2275(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate2276(.a(G7), .O(gate12inter7));
  inv1  gate2277(.a(G8), .O(gate12inter8));
  nand2 gate2278(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate2279(.a(s_247), .b(gate12inter3), .O(gate12inter10));
  nor2  gate2280(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate2281(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate2282(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );

  xor2  gate1821(.a(G12), .b(G11), .O(gate14inter0));
  nand2 gate1822(.a(gate14inter0), .b(s_182), .O(gate14inter1));
  and2  gate1823(.a(G12), .b(G11), .O(gate14inter2));
  inv1  gate1824(.a(s_182), .O(gate14inter3));
  inv1  gate1825(.a(s_183), .O(gate14inter4));
  nand2 gate1826(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate1827(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate1828(.a(G11), .O(gate14inter7));
  inv1  gate1829(.a(G12), .O(gate14inter8));
  nand2 gate1830(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate1831(.a(s_183), .b(gate14inter3), .O(gate14inter10));
  nor2  gate1832(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate1833(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate1834(.a(gate14inter12), .b(gate14inter1), .O(G281));

  xor2  gate2409(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate2410(.a(gate15inter0), .b(s_266), .O(gate15inter1));
  and2  gate2411(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate2412(.a(s_266), .O(gate15inter3));
  inv1  gate2413(.a(s_267), .O(gate15inter4));
  nand2 gate2414(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate2415(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate2416(.a(G13), .O(gate15inter7));
  inv1  gate2417(.a(G14), .O(gate15inter8));
  nand2 gate2418(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate2419(.a(s_267), .b(gate15inter3), .O(gate15inter10));
  nor2  gate2420(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate2421(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate2422(.a(gate15inter12), .b(gate15inter1), .O(G284));

  xor2  gate1009(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate1010(.a(gate16inter0), .b(s_66), .O(gate16inter1));
  and2  gate1011(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate1012(.a(s_66), .O(gate16inter3));
  inv1  gate1013(.a(s_67), .O(gate16inter4));
  nand2 gate1014(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate1015(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate1016(.a(G15), .O(gate16inter7));
  inv1  gate1017(.a(G16), .O(gate16inter8));
  nand2 gate1018(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate1019(.a(s_67), .b(gate16inter3), .O(gate16inter10));
  nor2  gate1020(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate1021(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate1022(.a(gate16inter12), .b(gate16inter1), .O(G287));

  xor2  gate1863(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate1864(.a(gate17inter0), .b(s_188), .O(gate17inter1));
  and2  gate1865(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate1866(.a(s_188), .O(gate17inter3));
  inv1  gate1867(.a(s_189), .O(gate17inter4));
  nand2 gate1868(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate1869(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate1870(.a(G17), .O(gate17inter7));
  inv1  gate1871(.a(G18), .O(gate17inter8));
  nand2 gate1872(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate1873(.a(s_189), .b(gate17inter3), .O(gate17inter10));
  nor2  gate1874(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate1875(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate1876(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate1765(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate1766(.a(gate19inter0), .b(s_174), .O(gate19inter1));
  and2  gate1767(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate1768(.a(s_174), .O(gate19inter3));
  inv1  gate1769(.a(s_175), .O(gate19inter4));
  nand2 gate1770(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate1771(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate1772(.a(G21), .O(gate19inter7));
  inv1  gate1773(.a(G22), .O(gate19inter8));
  nand2 gate1774(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate1775(.a(s_175), .b(gate19inter3), .O(gate19inter10));
  nor2  gate1776(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate1777(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate1778(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate883(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate884(.a(gate21inter0), .b(s_48), .O(gate21inter1));
  and2  gate885(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate886(.a(s_48), .O(gate21inter3));
  inv1  gate887(.a(s_49), .O(gate21inter4));
  nand2 gate888(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate889(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate890(.a(G25), .O(gate21inter7));
  inv1  gate891(.a(G26), .O(gate21inter8));
  nand2 gate892(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate893(.a(s_49), .b(gate21inter3), .O(gate21inter10));
  nor2  gate894(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate895(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate896(.a(gate21inter12), .b(gate21inter1), .O(G302));
nand2 gate22( .a(G27), .b(G28), .O(G305) );

  xor2  gate1205(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate1206(.a(gate23inter0), .b(s_94), .O(gate23inter1));
  and2  gate1207(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate1208(.a(s_94), .O(gate23inter3));
  inv1  gate1209(.a(s_95), .O(gate23inter4));
  nand2 gate1210(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate1211(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate1212(.a(G29), .O(gate23inter7));
  inv1  gate1213(.a(G30), .O(gate23inter8));
  nand2 gate1214(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate1215(.a(s_95), .b(gate23inter3), .O(gate23inter10));
  nor2  gate1216(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate1217(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate1218(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate1877(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate1878(.a(gate25inter0), .b(s_190), .O(gate25inter1));
  and2  gate1879(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate1880(.a(s_190), .O(gate25inter3));
  inv1  gate1881(.a(s_191), .O(gate25inter4));
  nand2 gate1882(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate1883(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate1884(.a(G1), .O(gate25inter7));
  inv1  gate1885(.a(G5), .O(gate25inter8));
  nand2 gate1886(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate1887(.a(s_191), .b(gate25inter3), .O(gate25inter10));
  nor2  gate1888(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate1889(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate1890(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate2717(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate2718(.a(gate27inter0), .b(s_310), .O(gate27inter1));
  and2  gate2719(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate2720(.a(s_310), .O(gate27inter3));
  inv1  gate2721(.a(s_311), .O(gate27inter4));
  nand2 gate2722(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate2723(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate2724(.a(G2), .O(gate27inter7));
  inv1  gate2725(.a(G6), .O(gate27inter8));
  nand2 gate2726(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate2727(.a(s_311), .b(gate27inter3), .O(gate27inter10));
  nor2  gate2728(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate2729(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate2730(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );

  xor2  gate2619(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate2620(.a(gate33inter0), .b(s_296), .O(gate33inter1));
  and2  gate2621(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate2622(.a(s_296), .O(gate33inter3));
  inv1  gate2623(.a(s_297), .O(gate33inter4));
  nand2 gate2624(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate2625(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate2626(.a(G17), .O(gate33inter7));
  inv1  gate2627(.a(G21), .O(gate33inter8));
  nand2 gate2628(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate2629(.a(s_297), .b(gate33inter3), .O(gate33inter10));
  nor2  gate2630(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate2631(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate2632(.a(gate33inter12), .b(gate33inter1), .O(G338));
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate1555(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate1556(.a(gate37inter0), .b(s_144), .O(gate37inter1));
  and2  gate1557(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate1558(.a(s_144), .O(gate37inter3));
  inv1  gate1559(.a(s_145), .O(gate37inter4));
  nand2 gate1560(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate1561(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate1562(.a(G19), .O(gate37inter7));
  inv1  gate1563(.a(G23), .O(gate37inter8));
  nand2 gate1564(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate1565(.a(s_145), .b(gate37inter3), .O(gate37inter10));
  nor2  gate1566(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate1567(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate1568(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );

  xor2  gate967(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate968(.a(gate40inter0), .b(s_60), .O(gate40inter1));
  and2  gate969(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate970(.a(s_60), .O(gate40inter3));
  inv1  gate971(.a(s_61), .O(gate40inter4));
  nand2 gate972(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate973(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate974(.a(G28), .O(gate40inter7));
  inv1  gate975(.a(G32), .O(gate40inter8));
  nand2 gate976(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate977(.a(s_61), .b(gate40inter3), .O(gate40inter10));
  nor2  gate978(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate979(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate980(.a(gate40inter12), .b(gate40inter1), .O(G359));
nand2 gate41( .a(G1), .b(G266), .O(G362) );

  xor2  gate1933(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate1934(.a(gate42inter0), .b(s_198), .O(gate42inter1));
  and2  gate1935(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate1936(.a(s_198), .O(gate42inter3));
  inv1  gate1937(.a(s_199), .O(gate42inter4));
  nand2 gate1938(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate1939(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate1940(.a(G2), .O(gate42inter7));
  inv1  gate1941(.a(G266), .O(gate42inter8));
  nand2 gate1942(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate1943(.a(s_199), .b(gate42inter3), .O(gate42inter10));
  nor2  gate1944(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate1945(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate1946(.a(gate42inter12), .b(gate42inter1), .O(G363));

  xor2  gate911(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate912(.a(gate43inter0), .b(s_52), .O(gate43inter1));
  and2  gate913(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate914(.a(s_52), .O(gate43inter3));
  inv1  gate915(.a(s_53), .O(gate43inter4));
  nand2 gate916(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate917(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate918(.a(G3), .O(gate43inter7));
  inv1  gate919(.a(G269), .O(gate43inter8));
  nand2 gate920(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate921(.a(s_53), .b(gate43inter3), .O(gate43inter10));
  nor2  gate922(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate923(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate924(.a(gate43inter12), .b(gate43inter1), .O(G364));

  xor2  gate1415(.a(G269), .b(G4), .O(gate44inter0));
  nand2 gate1416(.a(gate44inter0), .b(s_124), .O(gate44inter1));
  and2  gate1417(.a(G269), .b(G4), .O(gate44inter2));
  inv1  gate1418(.a(s_124), .O(gate44inter3));
  inv1  gate1419(.a(s_125), .O(gate44inter4));
  nand2 gate1420(.a(gate44inter4), .b(gate44inter3), .O(gate44inter5));
  nor2  gate1421(.a(gate44inter5), .b(gate44inter2), .O(gate44inter6));
  inv1  gate1422(.a(G4), .O(gate44inter7));
  inv1  gate1423(.a(G269), .O(gate44inter8));
  nand2 gate1424(.a(gate44inter8), .b(gate44inter7), .O(gate44inter9));
  nand2 gate1425(.a(s_125), .b(gate44inter3), .O(gate44inter10));
  nor2  gate1426(.a(gate44inter10), .b(gate44inter9), .O(gate44inter11));
  nor2  gate1427(.a(gate44inter11), .b(gate44inter6), .O(gate44inter12));
  nand2 gate1428(.a(gate44inter12), .b(gate44inter1), .O(G365));
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate1387(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate1388(.a(gate46inter0), .b(s_120), .O(gate46inter1));
  and2  gate1389(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate1390(.a(s_120), .O(gate46inter3));
  inv1  gate1391(.a(s_121), .O(gate46inter4));
  nand2 gate1392(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate1393(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate1394(.a(G6), .O(gate46inter7));
  inv1  gate1395(.a(G272), .O(gate46inter8));
  nand2 gate1396(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate1397(.a(s_121), .b(gate46inter3), .O(gate46inter10));
  nor2  gate1398(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate1399(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate1400(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );

  xor2  gate1247(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate1248(.a(gate50inter0), .b(s_100), .O(gate50inter1));
  and2  gate1249(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate1250(.a(s_100), .O(gate50inter3));
  inv1  gate1251(.a(s_101), .O(gate50inter4));
  nand2 gate1252(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate1253(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate1254(.a(G10), .O(gate50inter7));
  inv1  gate1255(.a(G278), .O(gate50inter8));
  nand2 gate1256(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate1257(.a(s_101), .b(gate50inter3), .O(gate50inter10));
  nor2  gate1258(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate1259(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate1260(.a(gate50inter12), .b(gate50inter1), .O(G371));
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate869(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate870(.a(gate54inter0), .b(s_46), .O(gate54inter1));
  and2  gate871(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate872(.a(s_46), .O(gate54inter3));
  inv1  gate873(.a(s_47), .O(gate54inter4));
  nand2 gate874(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate875(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate876(.a(G14), .O(gate54inter7));
  inv1  gate877(.a(G284), .O(gate54inter8));
  nand2 gate878(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate879(.a(s_47), .b(gate54inter3), .O(gate54inter10));
  nor2  gate880(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate881(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate882(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );

  xor2  gate2521(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate2522(.a(gate56inter0), .b(s_282), .O(gate56inter1));
  and2  gate2523(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate2524(.a(s_282), .O(gate56inter3));
  inv1  gate2525(.a(s_283), .O(gate56inter4));
  nand2 gate2526(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate2527(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate2528(.a(G16), .O(gate56inter7));
  inv1  gate2529(.a(G287), .O(gate56inter8));
  nand2 gate2530(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate2531(.a(s_283), .b(gate56inter3), .O(gate56inter10));
  nor2  gate2532(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate2533(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate2534(.a(gate56inter12), .b(gate56inter1), .O(G377));

  xor2  gate2451(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate2452(.a(gate57inter0), .b(s_272), .O(gate57inter1));
  and2  gate2453(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate2454(.a(s_272), .O(gate57inter3));
  inv1  gate2455(.a(s_273), .O(gate57inter4));
  nand2 gate2456(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate2457(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate2458(.a(G17), .O(gate57inter7));
  inv1  gate2459(.a(G290), .O(gate57inter8));
  nand2 gate2460(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate2461(.a(s_273), .b(gate57inter3), .O(gate57inter10));
  nor2  gate2462(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate2463(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate2464(.a(gate57inter12), .b(gate57inter1), .O(G378));

  xor2  gate925(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate926(.a(gate58inter0), .b(s_54), .O(gate58inter1));
  and2  gate927(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate928(.a(s_54), .O(gate58inter3));
  inv1  gate929(.a(s_55), .O(gate58inter4));
  nand2 gate930(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate931(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate932(.a(G18), .O(gate58inter7));
  inv1  gate933(.a(G290), .O(gate58inter8));
  nand2 gate934(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate935(.a(s_55), .b(gate58inter3), .O(gate58inter10));
  nor2  gate936(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate937(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate938(.a(gate58inter12), .b(gate58inter1), .O(G379));
nand2 gate59( .a(G19), .b(G293), .O(G380) );

  xor2  gate1163(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate1164(.a(gate60inter0), .b(s_88), .O(gate60inter1));
  and2  gate1165(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate1166(.a(s_88), .O(gate60inter3));
  inv1  gate1167(.a(s_89), .O(gate60inter4));
  nand2 gate1168(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate1169(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate1170(.a(G20), .O(gate60inter7));
  inv1  gate1171(.a(G293), .O(gate60inter8));
  nand2 gate1172(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate1173(.a(s_89), .b(gate60inter3), .O(gate60inter10));
  nor2  gate1174(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate1175(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate1176(.a(gate60inter12), .b(gate60inter1), .O(G381));

  xor2  gate1989(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate1990(.a(gate61inter0), .b(s_206), .O(gate61inter1));
  and2  gate1991(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate1992(.a(s_206), .O(gate61inter3));
  inv1  gate1993(.a(s_207), .O(gate61inter4));
  nand2 gate1994(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate1995(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate1996(.a(G21), .O(gate61inter7));
  inv1  gate1997(.a(G296), .O(gate61inter8));
  nand2 gate1998(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate1999(.a(s_207), .b(gate61inter3), .O(gate61inter10));
  nor2  gate2000(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate2001(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate2002(.a(gate61inter12), .b(gate61inter1), .O(G382));
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate1191(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate1192(.a(gate63inter0), .b(s_92), .O(gate63inter1));
  and2  gate1193(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate1194(.a(s_92), .O(gate63inter3));
  inv1  gate1195(.a(s_93), .O(gate63inter4));
  nand2 gate1196(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate1197(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate1198(.a(G23), .O(gate63inter7));
  inv1  gate1199(.a(G299), .O(gate63inter8));
  nand2 gate1200(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate1201(.a(s_93), .b(gate63inter3), .O(gate63inter10));
  nor2  gate1202(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate1203(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate1204(.a(gate63inter12), .b(gate63inter1), .O(G384));

  xor2  gate2983(.a(G299), .b(G24), .O(gate64inter0));
  nand2 gate2984(.a(gate64inter0), .b(s_348), .O(gate64inter1));
  and2  gate2985(.a(G299), .b(G24), .O(gate64inter2));
  inv1  gate2986(.a(s_348), .O(gate64inter3));
  inv1  gate2987(.a(s_349), .O(gate64inter4));
  nand2 gate2988(.a(gate64inter4), .b(gate64inter3), .O(gate64inter5));
  nor2  gate2989(.a(gate64inter5), .b(gate64inter2), .O(gate64inter6));
  inv1  gate2990(.a(G24), .O(gate64inter7));
  inv1  gate2991(.a(G299), .O(gate64inter8));
  nand2 gate2992(.a(gate64inter8), .b(gate64inter7), .O(gate64inter9));
  nand2 gate2993(.a(s_349), .b(gate64inter3), .O(gate64inter10));
  nor2  gate2994(.a(gate64inter10), .b(gate64inter9), .O(gate64inter11));
  nor2  gate2995(.a(gate64inter11), .b(gate64inter6), .O(gate64inter12));
  nand2 gate2996(.a(gate64inter12), .b(gate64inter1), .O(G385));

  xor2  gate2325(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate2326(.a(gate65inter0), .b(s_254), .O(gate65inter1));
  and2  gate2327(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate2328(.a(s_254), .O(gate65inter3));
  inv1  gate2329(.a(s_255), .O(gate65inter4));
  nand2 gate2330(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate2331(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate2332(.a(G25), .O(gate65inter7));
  inv1  gate2333(.a(G302), .O(gate65inter8));
  nand2 gate2334(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate2335(.a(s_255), .b(gate65inter3), .O(gate65inter10));
  nor2  gate2336(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate2337(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate2338(.a(gate65inter12), .b(gate65inter1), .O(G386));
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );

  xor2  gate2199(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate2200(.a(gate72inter0), .b(s_236), .O(gate72inter1));
  and2  gate2201(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate2202(.a(s_236), .O(gate72inter3));
  inv1  gate2203(.a(s_237), .O(gate72inter4));
  nand2 gate2204(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate2205(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate2206(.a(G32), .O(gate72inter7));
  inv1  gate2207(.a(G311), .O(gate72inter8));
  nand2 gate2208(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate2209(.a(s_237), .b(gate72inter3), .O(gate72inter10));
  nor2  gate2210(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate2211(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate2212(.a(gate72inter12), .b(gate72inter1), .O(G393));
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate645(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate646(.a(gate77inter0), .b(s_14), .O(gate77inter1));
  and2  gate647(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate648(.a(s_14), .O(gate77inter3));
  inv1  gate649(.a(s_15), .O(gate77inter4));
  nand2 gate650(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate651(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate652(.a(G2), .O(gate77inter7));
  inv1  gate653(.a(G320), .O(gate77inter8));
  nand2 gate654(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate655(.a(s_15), .b(gate77inter3), .O(gate77inter10));
  nor2  gate656(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate657(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate658(.a(gate77inter12), .b(gate77inter1), .O(G398));

  xor2  gate701(.a(G320), .b(G6), .O(gate78inter0));
  nand2 gate702(.a(gate78inter0), .b(s_22), .O(gate78inter1));
  and2  gate703(.a(G320), .b(G6), .O(gate78inter2));
  inv1  gate704(.a(s_22), .O(gate78inter3));
  inv1  gate705(.a(s_23), .O(gate78inter4));
  nand2 gate706(.a(gate78inter4), .b(gate78inter3), .O(gate78inter5));
  nor2  gate707(.a(gate78inter5), .b(gate78inter2), .O(gate78inter6));
  inv1  gate708(.a(G6), .O(gate78inter7));
  inv1  gate709(.a(G320), .O(gate78inter8));
  nand2 gate710(.a(gate78inter8), .b(gate78inter7), .O(gate78inter9));
  nand2 gate711(.a(s_23), .b(gate78inter3), .O(gate78inter10));
  nor2  gate712(.a(gate78inter10), .b(gate78inter9), .O(gate78inter11));
  nor2  gate713(.a(gate78inter11), .b(gate78inter6), .O(gate78inter12));
  nand2 gate714(.a(gate78inter12), .b(gate78inter1), .O(G399));
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate617(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate618(.a(gate81inter0), .b(s_10), .O(gate81inter1));
  and2  gate619(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate620(.a(s_10), .O(gate81inter3));
  inv1  gate621(.a(s_11), .O(gate81inter4));
  nand2 gate622(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate623(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate624(.a(G3), .O(gate81inter7));
  inv1  gate625(.a(G326), .O(gate81inter8));
  nand2 gate626(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate627(.a(s_11), .b(gate81inter3), .O(gate81inter10));
  nor2  gate628(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate629(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate630(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );

  xor2  gate1429(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate1430(.a(gate83inter0), .b(s_126), .O(gate83inter1));
  and2  gate1431(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate1432(.a(s_126), .O(gate83inter3));
  inv1  gate1433(.a(s_127), .O(gate83inter4));
  nand2 gate1434(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate1435(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate1436(.a(G11), .O(gate83inter7));
  inv1  gate1437(.a(G329), .O(gate83inter8));
  nand2 gate1438(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate1439(.a(s_127), .b(gate83inter3), .O(gate83inter10));
  nor2  gate1440(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate1441(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate1442(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );

  xor2  gate729(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate730(.a(gate86inter0), .b(s_26), .O(gate86inter1));
  and2  gate731(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate732(.a(s_26), .O(gate86inter3));
  inv1  gate733(.a(s_27), .O(gate86inter4));
  nand2 gate734(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate735(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate736(.a(G8), .O(gate86inter7));
  inv1  gate737(.a(G332), .O(gate86inter8));
  nand2 gate738(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate739(.a(s_27), .b(gate86inter3), .O(gate86inter10));
  nor2  gate740(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate741(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate742(.a(gate86inter12), .b(gate86inter1), .O(G407));

  xor2  gate1177(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate1178(.a(gate87inter0), .b(s_90), .O(gate87inter1));
  and2  gate1179(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate1180(.a(s_90), .O(gate87inter3));
  inv1  gate1181(.a(s_91), .O(gate87inter4));
  nand2 gate1182(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate1183(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate1184(.a(G12), .O(gate87inter7));
  inv1  gate1185(.a(G335), .O(gate87inter8));
  nand2 gate1186(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate1187(.a(s_91), .b(gate87inter3), .O(gate87inter10));
  nor2  gate1188(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate1189(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate1190(.a(gate87inter12), .b(gate87inter1), .O(G408));

  xor2  gate1457(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate1458(.a(gate88inter0), .b(s_130), .O(gate88inter1));
  and2  gate1459(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate1460(.a(s_130), .O(gate88inter3));
  inv1  gate1461(.a(s_131), .O(gate88inter4));
  nand2 gate1462(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate1463(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate1464(.a(G16), .O(gate88inter7));
  inv1  gate1465(.a(G335), .O(gate88inter8));
  nand2 gate1466(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate1467(.a(s_131), .b(gate88inter3), .O(gate88inter10));
  nor2  gate1468(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate1469(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate1470(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate2465(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate2466(.a(gate90inter0), .b(s_274), .O(gate90inter1));
  and2  gate2467(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate2468(.a(s_274), .O(gate90inter3));
  inv1  gate2469(.a(s_275), .O(gate90inter4));
  nand2 gate2470(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate2471(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate2472(.a(G21), .O(gate90inter7));
  inv1  gate2473(.a(G338), .O(gate90inter8));
  nand2 gate2474(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate2475(.a(s_275), .b(gate90inter3), .O(gate90inter10));
  nor2  gate2476(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate2477(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate2478(.a(gate90inter12), .b(gate90inter1), .O(G411));
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate1121(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate1122(.a(gate95inter0), .b(s_82), .O(gate95inter1));
  and2  gate1123(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate1124(.a(s_82), .O(gate95inter3));
  inv1  gate1125(.a(s_83), .O(gate95inter4));
  nand2 gate1126(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate1127(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate1128(.a(G26), .O(gate95inter7));
  inv1  gate1129(.a(G347), .O(gate95inter8));
  nand2 gate1130(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate1131(.a(s_83), .b(gate95inter3), .O(gate95inter10));
  nor2  gate1132(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate1133(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate1134(.a(gate95inter12), .b(gate95inter1), .O(G416));

  xor2  gate2381(.a(G347), .b(G30), .O(gate96inter0));
  nand2 gate2382(.a(gate96inter0), .b(s_262), .O(gate96inter1));
  and2  gate2383(.a(G347), .b(G30), .O(gate96inter2));
  inv1  gate2384(.a(s_262), .O(gate96inter3));
  inv1  gate2385(.a(s_263), .O(gate96inter4));
  nand2 gate2386(.a(gate96inter4), .b(gate96inter3), .O(gate96inter5));
  nor2  gate2387(.a(gate96inter5), .b(gate96inter2), .O(gate96inter6));
  inv1  gate2388(.a(G30), .O(gate96inter7));
  inv1  gate2389(.a(G347), .O(gate96inter8));
  nand2 gate2390(.a(gate96inter8), .b(gate96inter7), .O(gate96inter9));
  nand2 gate2391(.a(s_263), .b(gate96inter3), .O(gate96inter10));
  nor2  gate2392(.a(gate96inter10), .b(gate96inter9), .O(gate96inter11));
  nor2  gate2393(.a(gate96inter11), .b(gate96inter6), .O(gate96inter12));
  nand2 gate2394(.a(gate96inter12), .b(gate96inter1), .O(G417));
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate1905(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate1906(.a(gate100inter0), .b(s_194), .O(gate100inter1));
  and2  gate1907(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate1908(.a(s_194), .O(gate100inter3));
  inv1  gate1909(.a(s_195), .O(gate100inter4));
  nand2 gate1910(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate1911(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate1912(.a(G31), .O(gate100inter7));
  inv1  gate1913(.a(G353), .O(gate100inter8));
  nand2 gate1914(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate1915(.a(s_195), .b(gate100inter3), .O(gate100inter10));
  nor2  gate1916(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate1917(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate1918(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate2787(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate2788(.a(gate102inter0), .b(s_320), .O(gate102inter1));
  and2  gate2789(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate2790(.a(s_320), .O(gate102inter3));
  inv1  gate2791(.a(s_321), .O(gate102inter4));
  nand2 gate2792(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate2793(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate2794(.a(G24), .O(gate102inter7));
  inv1  gate2795(.a(G356), .O(gate102inter8));
  nand2 gate2796(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate2797(.a(s_321), .b(gate102inter3), .O(gate102inter10));
  nor2  gate2798(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate2799(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate2800(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate2115(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate2116(.a(gate104inter0), .b(s_224), .O(gate104inter1));
  and2  gate2117(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate2118(.a(s_224), .O(gate104inter3));
  inv1  gate2119(.a(s_225), .O(gate104inter4));
  nand2 gate2120(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate2121(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate2122(.a(G32), .O(gate104inter7));
  inv1  gate2123(.a(G359), .O(gate104inter8));
  nand2 gate2124(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate2125(.a(s_225), .b(gate104inter3), .O(gate104inter10));
  nor2  gate2126(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate2127(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate2128(.a(gate104inter12), .b(gate104inter1), .O(G425));
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );

  xor2  gate1611(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate1612(.a(gate111inter0), .b(s_152), .O(gate111inter1));
  and2  gate1613(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate1614(.a(s_152), .O(gate111inter3));
  inv1  gate1615(.a(s_153), .O(gate111inter4));
  nand2 gate1616(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate1617(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate1618(.a(G374), .O(gate111inter7));
  inv1  gate1619(.a(G375), .O(gate111inter8));
  nand2 gate1620(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate1621(.a(s_153), .b(gate111inter3), .O(gate111inter10));
  nor2  gate1622(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate1623(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate1624(.a(gate111inter12), .b(gate111inter1), .O(G444));

  xor2  gate2955(.a(G377), .b(G376), .O(gate112inter0));
  nand2 gate2956(.a(gate112inter0), .b(s_344), .O(gate112inter1));
  and2  gate2957(.a(G377), .b(G376), .O(gate112inter2));
  inv1  gate2958(.a(s_344), .O(gate112inter3));
  inv1  gate2959(.a(s_345), .O(gate112inter4));
  nand2 gate2960(.a(gate112inter4), .b(gate112inter3), .O(gate112inter5));
  nor2  gate2961(.a(gate112inter5), .b(gate112inter2), .O(gate112inter6));
  inv1  gate2962(.a(G376), .O(gate112inter7));
  inv1  gate2963(.a(G377), .O(gate112inter8));
  nand2 gate2964(.a(gate112inter8), .b(gate112inter7), .O(gate112inter9));
  nand2 gate2965(.a(s_345), .b(gate112inter3), .O(gate112inter10));
  nor2  gate2966(.a(gate112inter10), .b(gate112inter9), .O(gate112inter11));
  nor2  gate2967(.a(gate112inter11), .b(gate112inter6), .O(gate112inter12));
  nand2 gate2968(.a(gate112inter12), .b(gate112inter1), .O(G447));

  xor2  gate757(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate758(.a(gate113inter0), .b(s_30), .O(gate113inter1));
  and2  gate759(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate760(.a(s_30), .O(gate113inter3));
  inv1  gate761(.a(s_31), .O(gate113inter4));
  nand2 gate762(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate763(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate764(.a(G378), .O(gate113inter7));
  inv1  gate765(.a(G379), .O(gate113inter8));
  nand2 gate766(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate767(.a(s_31), .b(gate113inter3), .O(gate113inter10));
  nor2  gate768(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate769(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate770(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate2577(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate2578(.a(gate117inter0), .b(s_290), .O(gate117inter1));
  and2  gate2579(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate2580(.a(s_290), .O(gate117inter3));
  inv1  gate2581(.a(s_291), .O(gate117inter4));
  nand2 gate2582(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate2583(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate2584(.a(G386), .O(gate117inter7));
  inv1  gate2585(.a(G387), .O(gate117inter8));
  nand2 gate2586(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate2587(.a(s_291), .b(gate117inter3), .O(gate117inter10));
  nor2  gate2588(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate2589(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate2590(.a(gate117inter12), .b(gate117inter1), .O(G462));

  xor2  gate2647(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate2648(.a(gate118inter0), .b(s_300), .O(gate118inter1));
  and2  gate2649(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate2650(.a(s_300), .O(gate118inter3));
  inv1  gate2651(.a(s_301), .O(gate118inter4));
  nand2 gate2652(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate2653(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate2654(.a(G388), .O(gate118inter7));
  inv1  gate2655(.a(G389), .O(gate118inter8));
  nand2 gate2656(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate2657(.a(s_301), .b(gate118inter3), .O(gate118inter10));
  nor2  gate2658(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate2659(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate2660(.a(gate118inter12), .b(gate118inter1), .O(G465));

  xor2  gate603(.a(G391), .b(G390), .O(gate119inter0));
  nand2 gate604(.a(gate119inter0), .b(s_8), .O(gate119inter1));
  and2  gate605(.a(G391), .b(G390), .O(gate119inter2));
  inv1  gate606(.a(s_8), .O(gate119inter3));
  inv1  gate607(.a(s_9), .O(gate119inter4));
  nand2 gate608(.a(gate119inter4), .b(gate119inter3), .O(gate119inter5));
  nor2  gate609(.a(gate119inter5), .b(gate119inter2), .O(gate119inter6));
  inv1  gate610(.a(G390), .O(gate119inter7));
  inv1  gate611(.a(G391), .O(gate119inter8));
  nand2 gate612(.a(gate119inter8), .b(gate119inter7), .O(gate119inter9));
  nand2 gate613(.a(s_9), .b(gate119inter3), .O(gate119inter10));
  nor2  gate614(.a(gate119inter10), .b(gate119inter9), .O(gate119inter11));
  nor2  gate615(.a(gate119inter11), .b(gate119inter6), .O(gate119inter12));
  nand2 gate616(.a(gate119inter12), .b(gate119inter1), .O(G468));
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate2773(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate2774(.a(gate125inter0), .b(s_318), .O(gate125inter1));
  and2  gate2775(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate2776(.a(s_318), .O(gate125inter3));
  inv1  gate2777(.a(s_319), .O(gate125inter4));
  nand2 gate2778(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate2779(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate2780(.a(G402), .O(gate125inter7));
  inv1  gate2781(.a(G403), .O(gate125inter8));
  nand2 gate2782(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate2783(.a(s_319), .b(gate125inter3), .O(gate125inter10));
  nor2  gate2784(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate2785(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate2786(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );

  xor2  gate1485(.a(G417), .b(G416), .O(gate132inter0));
  nand2 gate1486(.a(gate132inter0), .b(s_134), .O(gate132inter1));
  and2  gate1487(.a(G417), .b(G416), .O(gate132inter2));
  inv1  gate1488(.a(s_134), .O(gate132inter3));
  inv1  gate1489(.a(s_135), .O(gate132inter4));
  nand2 gate1490(.a(gate132inter4), .b(gate132inter3), .O(gate132inter5));
  nor2  gate1491(.a(gate132inter5), .b(gate132inter2), .O(gate132inter6));
  inv1  gate1492(.a(G416), .O(gate132inter7));
  inv1  gate1493(.a(G417), .O(gate132inter8));
  nand2 gate1494(.a(gate132inter8), .b(gate132inter7), .O(gate132inter9));
  nand2 gate1495(.a(s_135), .b(gate132inter3), .O(gate132inter10));
  nor2  gate1496(.a(gate132inter10), .b(gate132inter9), .O(gate132inter11));
  nor2  gate1497(.a(gate132inter11), .b(gate132inter6), .O(gate132inter12));
  nand2 gate1498(.a(gate132inter12), .b(gate132inter1), .O(G507));
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate1051(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate1052(.a(gate136inter0), .b(s_72), .O(gate136inter1));
  and2  gate1053(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate1054(.a(s_72), .O(gate136inter3));
  inv1  gate1055(.a(s_73), .O(gate136inter4));
  nand2 gate1056(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate1057(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate1058(.a(G424), .O(gate136inter7));
  inv1  gate1059(.a(G425), .O(gate136inter8));
  nand2 gate1060(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate1061(.a(s_73), .b(gate136inter3), .O(gate136inter10));
  nor2  gate1062(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate1063(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate1064(.a(gate136inter12), .b(gate136inter1), .O(G519));

  xor2  gate1709(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate1710(.a(gate137inter0), .b(s_166), .O(gate137inter1));
  and2  gate1711(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate1712(.a(s_166), .O(gate137inter3));
  inv1  gate1713(.a(s_167), .O(gate137inter4));
  nand2 gate1714(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate1715(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate1716(.a(G426), .O(gate137inter7));
  inv1  gate1717(.a(G429), .O(gate137inter8));
  nand2 gate1718(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate1719(.a(s_167), .b(gate137inter3), .O(gate137inter10));
  nor2  gate1720(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate1721(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate1722(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );

  xor2  gate1807(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate1808(.a(gate141inter0), .b(s_180), .O(gate141inter1));
  and2  gate1809(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate1810(.a(s_180), .O(gate141inter3));
  inv1  gate1811(.a(s_181), .O(gate141inter4));
  nand2 gate1812(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate1813(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate1814(.a(G450), .O(gate141inter7));
  inv1  gate1815(.a(G453), .O(gate141inter8));
  nand2 gate1816(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate1817(.a(s_181), .b(gate141inter3), .O(gate141inter10));
  nor2  gate1818(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate1819(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate1820(.a(gate141inter12), .b(gate141inter1), .O(G534));
nand2 gate142( .a(G456), .b(G459), .O(G537) );

  xor2  gate1345(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate1346(.a(gate143inter0), .b(s_114), .O(gate143inter1));
  and2  gate1347(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate1348(.a(s_114), .O(gate143inter3));
  inv1  gate1349(.a(s_115), .O(gate143inter4));
  nand2 gate1350(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate1351(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate1352(.a(G462), .O(gate143inter7));
  inv1  gate1353(.a(G465), .O(gate143inter8));
  nand2 gate1354(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate1355(.a(s_115), .b(gate143inter3), .O(gate143inter10));
  nor2  gate1356(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate1357(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate1358(.a(gate143inter12), .b(gate143inter1), .O(G540));

  xor2  gate2017(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate2018(.a(gate144inter0), .b(s_210), .O(gate144inter1));
  and2  gate2019(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate2020(.a(s_210), .O(gate144inter3));
  inv1  gate2021(.a(s_211), .O(gate144inter4));
  nand2 gate2022(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate2023(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate2024(.a(G468), .O(gate144inter7));
  inv1  gate2025(.a(G471), .O(gate144inter8));
  nand2 gate2026(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate2027(.a(s_211), .b(gate144inter3), .O(gate144inter10));
  nor2  gate2028(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate2029(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate2030(.a(gate144inter12), .b(gate144inter1), .O(G543));

  xor2  gate2675(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate2676(.a(gate145inter0), .b(s_304), .O(gate145inter1));
  and2  gate2677(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate2678(.a(s_304), .O(gate145inter3));
  inv1  gate2679(.a(s_305), .O(gate145inter4));
  nand2 gate2680(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate2681(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate2682(.a(G474), .O(gate145inter7));
  inv1  gate2683(.a(G477), .O(gate145inter8));
  nand2 gate2684(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate2685(.a(s_305), .b(gate145inter3), .O(gate145inter10));
  nor2  gate2686(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate2687(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate2688(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );

  xor2  gate2045(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate2046(.a(gate147inter0), .b(s_214), .O(gate147inter1));
  and2  gate2047(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate2048(.a(s_214), .O(gate147inter3));
  inv1  gate2049(.a(s_215), .O(gate147inter4));
  nand2 gate2050(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate2051(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate2052(.a(G486), .O(gate147inter7));
  inv1  gate2053(.a(G489), .O(gate147inter8));
  nand2 gate2054(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate2055(.a(s_215), .b(gate147inter3), .O(gate147inter10));
  nor2  gate2056(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate2057(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate2058(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate1443(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate1444(.a(gate149inter0), .b(s_128), .O(gate149inter1));
  and2  gate1445(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate1446(.a(s_128), .O(gate149inter3));
  inv1  gate1447(.a(s_129), .O(gate149inter4));
  nand2 gate1448(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate1449(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate1450(.a(G498), .O(gate149inter7));
  inv1  gate1451(.a(G501), .O(gate149inter8));
  nand2 gate1452(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate1453(.a(s_129), .b(gate149inter3), .O(gate149inter10));
  nor2  gate1454(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate1455(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate1456(.a(gate149inter12), .b(gate149inter1), .O(G558));

  xor2  gate2703(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate2704(.a(gate150inter0), .b(s_308), .O(gate150inter1));
  and2  gate2705(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate2706(.a(s_308), .O(gate150inter3));
  inv1  gate2707(.a(s_309), .O(gate150inter4));
  nand2 gate2708(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate2709(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate2710(.a(G504), .O(gate150inter7));
  inv1  gate2711(.a(G507), .O(gate150inter8));
  nand2 gate2712(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate2713(.a(s_309), .b(gate150inter3), .O(gate150inter10));
  nor2  gate2714(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate2715(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate2716(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate1079(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate1080(.a(gate153inter0), .b(s_76), .O(gate153inter1));
  and2  gate1081(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate1082(.a(s_76), .O(gate153inter3));
  inv1  gate1083(.a(s_77), .O(gate153inter4));
  nand2 gate1084(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate1085(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate1086(.a(G426), .O(gate153inter7));
  inv1  gate1087(.a(G522), .O(gate153inter8));
  nand2 gate1088(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate1089(.a(s_77), .b(gate153inter3), .O(gate153inter10));
  nor2  gate1090(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate1091(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate1092(.a(gate153inter12), .b(gate153inter1), .O(G570));

  xor2  gate2479(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate2480(.a(gate154inter0), .b(s_276), .O(gate154inter1));
  and2  gate2481(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate2482(.a(s_276), .O(gate154inter3));
  inv1  gate2483(.a(s_277), .O(gate154inter4));
  nand2 gate2484(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate2485(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate2486(.a(G429), .O(gate154inter7));
  inv1  gate2487(.a(G522), .O(gate154inter8));
  nand2 gate2488(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate2489(.a(s_277), .b(gate154inter3), .O(gate154inter10));
  nor2  gate2490(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate2491(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate2492(.a(gate154inter12), .b(gate154inter1), .O(G571));

  xor2  gate1093(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate1094(.a(gate155inter0), .b(s_78), .O(gate155inter1));
  and2  gate1095(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate1096(.a(s_78), .O(gate155inter3));
  inv1  gate1097(.a(s_79), .O(gate155inter4));
  nand2 gate1098(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1099(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1100(.a(G432), .O(gate155inter7));
  inv1  gate1101(.a(G525), .O(gate155inter8));
  nand2 gate1102(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1103(.a(s_79), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1104(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1105(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1106(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate2591(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate2592(.a(gate159inter0), .b(s_292), .O(gate159inter1));
  and2  gate2593(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate2594(.a(s_292), .O(gate159inter3));
  inv1  gate2595(.a(s_293), .O(gate159inter4));
  nand2 gate2596(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate2597(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate2598(.a(G444), .O(gate159inter7));
  inv1  gate2599(.a(G531), .O(gate159inter8));
  nand2 gate2600(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate2601(.a(s_293), .b(gate159inter3), .O(gate159inter10));
  nor2  gate2602(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate2603(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate2604(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate2689(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate2690(.a(gate162inter0), .b(s_306), .O(gate162inter1));
  and2  gate2691(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate2692(.a(s_306), .O(gate162inter3));
  inv1  gate2693(.a(s_307), .O(gate162inter4));
  nand2 gate2694(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate2695(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate2696(.a(G453), .O(gate162inter7));
  inv1  gate2697(.a(G534), .O(gate162inter8));
  nand2 gate2698(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate2699(.a(s_307), .b(gate162inter3), .O(gate162inter10));
  nor2  gate2700(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate2701(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate2702(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate2997(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate2998(.a(gate165inter0), .b(s_350), .O(gate165inter1));
  and2  gate2999(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate3000(.a(s_350), .O(gate165inter3));
  inv1  gate3001(.a(s_351), .O(gate165inter4));
  nand2 gate3002(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate3003(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate3004(.a(G462), .O(gate165inter7));
  inv1  gate3005(.a(G540), .O(gate165inter8));
  nand2 gate3006(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate3007(.a(s_351), .b(gate165inter3), .O(gate165inter10));
  nor2  gate3008(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate3009(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate3010(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );

  xor2  gate2843(.a(G546), .b(G474), .O(gate169inter0));
  nand2 gate2844(.a(gate169inter0), .b(s_328), .O(gate169inter1));
  and2  gate2845(.a(G546), .b(G474), .O(gate169inter2));
  inv1  gate2846(.a(s_328), .O(gate169inter3));
  inv1  gate2847(.a(s_329), .O(gate169inter4));
  nand2 gate2848(.a(gate169inter4), .b(gate169inter3), .O(gate169inter5));
  nor2  gate2849(.a(gate169inter5), .b(gate169inter2), .O(gate169inter6));
  inv1  gate2850(.a(G474), .O(gate169inter7));
  inv1  gate2851(.a(G546), .O(gate169inter8));
  nand2 gate2852(.a(gate169inter8), .b(gate169inter7), .O(gate169inter9));
  nand2 gate2853(.a(s_329), .b(gate169inter3), .O(gate169inter10));
  nor2  gate2854(.a(gate169inter10), .b(gate169inter9), .O(gate169inter11));
  nor2  gate2855(.a(gate169inter11), .b(gate169inter6), .O(gate169inter12));
  nand2 gate2856(.a(gate169inter12), .b(gate169inter1), .O(G586));
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate1219(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate1220(.a(gate175inter0), .b(s_96), .O(gate175inter1));
  and2  gate1221(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate1222(.a(s_96), .O(gate175inter3));
  inv1  gate1223(.a(s_97), .O(gate175inter4));
  nand2 gate1224(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1225(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1226(.a(G492), .O(gate175inter7));
  inv1  gate1227(.a(G555), .O(gate175inter8));
  nand2 gate1228(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1229(.a(s_97), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1230(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1231(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1232(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );

  xor2  gate2745(.a(G558), .b(G498), .O(gate177inter0));
  nand2 gate2746(.a(gate177inter0), .b(s_314), .O(gate177inter1));
  and2  gate2747(.a(G558), .b(G498), .O(gate177inter2));
  inv1  gate2748(.a(s_314), .O(gate177inter3));
  inv1  gate2749(.a(s_315), .O(gate177inter4));
  nand2 gate2750(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate2751(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate2752(.a(G498), .O(gate177inter7));
  inv1  gate2753(.a(G558), .O(gate177inter8));
  nand2 gate2754(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate2755(.a(s_315), .b(gate177inter3), .O(gate177inter10));
  nor2  gate2756(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate2757(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate2758(.a(gate177inter12), .b(gate177inter1), .O(G594));
nand2 gate178( .a(G501), .b(G558), .O(G595) );

  xor2  gate1513(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate1514(.a(gate179inter0), .b(s_138), .O(gate179inter1));
  and2  gate1515(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate1516(.a(s_138), .O(gate179inter3));
  inv1  gate1517(.a(s_139), .O(gate179inter4));
  nand2 gate1518(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate1519(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate1520(.a(G504), .O(gate179inter7));
  inv1  gate1521(.a(G561), .O(gate179inter8));
  nand2 gate1522(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate1523(.a(s_139), .b(gate179inter3), .O(gate179inter10));
  nor2  gate1524(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate1525(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate1526(.a(gate179inter12), .b(gate179inter1), .O(G596));
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate1737(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate1738(.a(gate183inter0), .b(s_170), .O(gate183inter1));
  and2  gate1739(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate1740(.a(s_170), .O(gate183inter3));
  inv1  gate1741(.a(s_171), .O(gate183inter4));
  nand2 gate1742(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate1743(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate1744(.a(G516), .O(gate183inter7));
  inv1  gate1745(.a(G567), .O(gate183inter8));
  nand2 gate1746(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate1747(.a(s_171), .b(gate183inter3), .O(gate183inter10));
  nor2  gate1748(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate1749(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate1750(.a(gate183inter12), .b(gate183inter1), .O(G600));

  xor2  gate2507(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate2508(.a(gate184inter0), .b(s_280), .O(gate184inter1));
  and2  gate2509(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate2510(.a(s_280), .O(gate184inter3));
  inv1  gate2511(.a(s_281), .O(gate184inter4));
  nand2 gate2512(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate2513(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate2514(.a(G519), .O(gate184inter7));
  inv1  gate2515(.a(G567), .O(gate184inter8));
  nand2 gate2516(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate2517(.a(s_281), .b(gate184inter3), .O(gate184inter10));
  nor2  gate2518(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate2519(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate2520(.a(gate184inter12), .b(gate184inter1), .O(G601));

  xor2  gate2815(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate2816(.a(gate185inter0), .b(s_324), .O(gate185inter1));
  and2  gate2817(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate2818(.a(s_324), .O(gate185inter3));
  inv1  gate2819(.a(s_325), .O(gate185inter4));
  nand2 gate2820(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate2821(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate2822(.a(G570), .O(gate185inter7));
  inv1  gate2823(.a(G571), .O(gate185inter8));
  nand2 gate2824(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate2825(.a(s_325), .b(gate185inter3), .O(gate185inter10));
  nor2  gate2826(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate2827(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate2828(.a(gate185inter12), .b(gate185inter1), .O(G602));

  xor2  gate2549(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate2550(.a(gate186inter0), .b(s_286), .O(gate186inter1));
  and2  gate2551(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate2552(.a(s_286), .O(gate186inter3));
  inv1  gate2553(.a(s_287), .O(gate186inter4));
  nand2 gate2554(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate2555(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate2556(.a(G572), .O(gate186inter7));
  inv1  gate2557(.a(G573), .O(gate186inter8));
  nand2 gate2558(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate2559(.a(s_287), .b(gate186inter3), .O(gate186inter10));
  nor2  gate2560(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate2561(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate2562(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate589(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate590(.a(gate188inter0), .b(s_6), .O(gate188inter1));
  and2  gate591(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate592(.a(s_6), .O(gate188inter3));
  inv1  gate593(.a(s_7), .O(gate188inter4));
  nand2 gate594(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate595(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate596(.a(G576), .O(gate188inter7));
  inv1  gate597(.a(G577), .O(gate188inter8));
  nand2 gate598(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate599(.a(s_7), .b(gate188inter3), .O(gate188inter10));
  nor2  gate600(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate601(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate602(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate2185(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate2186(.a(gate191inter0), .b(s_234), .O(gate191inter1));
  and2  gate2187(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate2188(.a(s_234), .O(gate191inter3));
  inv1  gate2189(.a(s_235), .O(gate191inter4));
  nand2 gate2190(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate2191(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate2192(.a(G582), .O(gate191inter7));
  inv1  gate2193(.a(G583), .O(gate191inter8));
  nand2 gate2194(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate2195(.a(s_235), .b(gate191inter3), .O(gate191inter10));
  nor2  gate2196(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate2197(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate2198(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate2731(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate2732(.a(gate193inter0), .b(s_312), .O(gate193inter1));
  and2  gate2733(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate2734(.a(s_312), .O(gate193inter3));
  inv1  gate2735(.a(s_313), .O(gate193inter4));
  nand2 gate2736(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate2737(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate2738(.a(G586), .O(gate193inter7));
  inv1  gate2739(.a(G587), .O(gate193inter8));
  nand2 gate2740(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate2741(.a(s_313), .b(gate193inter3), .O(gate193inter10));
  nor2  gate2742(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate2743(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate2744(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate897(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate898(.a(gate196inter0), .b(s_50), .O(gate196inter1));
  and2  gate899(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate900(.a(s_50), .O(gate196inter3));
  inv1  gate901(.a(s_51), .O(gate196inter4));
  nand2 gate902(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate903(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate904(.a(G592), .O(gate196inter7));
  inv1  gate905(.a(G593), .O(gate196inter8));
  nand2 gate906(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate907(.a(s_51), .b(gate196inter3), .O(gate196inter10));
  nor2  gate908(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate909(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate910(.a(gate196inter12), .b(gate196inter1), .O(G651));

  xor2  gate1793(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate1794(.a(gate197inter0), .b(s_178), .O(gate197inter1));
  and2  gate1795(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate1796(.a(s_178), .O(gate197inter3));
  inv1  gate1797(.a(s_179), .O(gate197inter4));
  nand2 gate1798(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate1799(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate1800(.a(G594), .O(gate197inter7));
  inv1  gate1801(.a(G595), .O(gate197inter8));
  nand2 gate1802(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate1803(.a(s_179), .b(gate197inter3), .O(gate197inter10));
  nor2  gate1804(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate1805(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate1806(.a(gate197inter12), .b(gate197inter1), .O(G654));
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate1275(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate1276(.a(gate201inter0), .b(s_104), .O(gate201inter1));
  and2  gate1277(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate1278(.a(s_104), .O(gate201inter3));
  inv1  gate1279(.a(s_105), .O(gate201inter4));
  nand2 gate1280(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate1281(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate1282(.a(G602), .O(gate201inter7));
  inv1  gate1283(.a(G607), .O(gate201inter8));
  nand2 gate1284(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate1285(.a(s_105), .b(gate201inter3), .O(gate201inter10));
  nor2  gate1286(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate1287(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate1288(.a(gate201inter12), .b(gate201inter1), .O(G666));

  xor2  gate1751(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate1752(.a(gate202inter0), .b(s_172), .O(gate202inter1));
  and2  gate1753(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate1754(.a(s_172), .O(gate202inter3));
  inv1  gate1755(.a(s_173), .O(gate202inter4));
  nand2 gate1756(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate1757(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate1758(.a(G612), .O(gate202inter7));
  inv1  gate1759(.a(G617), .O(gate202inter8));
  nand2 gate1760(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate1761(.a(s_173), .b(gate202inter3), .O(gate202inter10));
  nor2  gate1762(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate1763(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate1764(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate1261(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate1262(.a(gate206inter0), .b(s_102), .O(gate206inter1));
  and2  gate1263(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate1264(.a(s_102), .O(gate206inter3));
  inv1  gate1265(.a(s_103), .O(gate206inter4));
  nand2 gate1266(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate1267(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate1268(.a(G632), .O(gate206inter7));
  inv1  gate1269(.a(G637), .O(gate206inter8));
  nand2 gate1270(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate1271(.a(s_103), .b(gate206inter3), .O(gate206inter10));
  nor2  gate1272(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate1273(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate1274(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate2423(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate2424(.a(gate211inter0), .b(s_268), .O(gate211inter1));
  and2  gate2425(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate2426(.a(s_268), .O(gate211inter3));
  inv1  gate2427(.a(s_269), .O(gate211inter4));
  nand2 gate2428(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate2429(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate2430(.a(G612), .O(gate211inter7));
  inv1  gate2431(.a(G669), .O(gate211inter8));
  nand2 gate2432(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate2433(.a(s_269), .b(gate211inter3), .O(gate211inter10));
  nor2  gate2434(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate2435(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate2436(.a(gate211inter12), .b(gate211inter1), .O(G692));

  xor2  gate1947(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate1948(.a(gate212inter0), .b(s_200), .O(gate212inter1));
  and2  gate1949(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate1950(.a(s_200), .O(gate212inter3));
  inv1  gate1951(.a(s_201), .O(gate212inter4));
  nand2 gate1952(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate1953(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate1954(.a(G617), .O(gate212inter7));
  inv1  gate1955(.a(G669), .O(gate212inter8));
  nand2 gate1956(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate1957(.a(s_201), .b(gate212inter3), .O(gate212inter10));
  nor2  gate1958(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate1959(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate1960(.a(gate212inter12), .b(gate212inter1), .O(G693));

  xor2  gate1681(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate1682(.a(gate213inter0), .b(s_162), .O(gate213inter1));
  and2  gate1683(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate1684(.a(s_162), .O(gate213inter3));
  inv1  gate1685(.a(s_163), .O(gate213inter4));
  nand2 gate1686(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate1687(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate1688(.a(G602), .O(gate213inter7));
  inv1  gate1689(.a(G672), .O(gate213inter8));
  nand2 gate1690(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate1691(.a(s_163), .b(gate213inter3), .O(gate213inter10));
  nor2  gate1692(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate1693(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate1694(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate1023(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate1024(.a(gate216inter0), .b(s_68), .O(gate216inter1));
  and2  gate1025(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate1026(.a(s_68), .O(gate216inter3));
  inv1  gate1027(.a(s_69), .O(gate216inter4));
  nand2 gate1028(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate1029(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate1030(.a(G617), .O(gate216inter7));
  inv1  gate1031(.a(G675), .O(gate216inter8));
  nand2 gate1032(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate1033(.a(s_69), .b(gate216inter3), .O(gate216inter10));
  nor2  gate1034(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate1035(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate1036(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate1975(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate1976(.a(gate220inter0), .b(s_204), .O(gate220inter1));
  and2  gate1977(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate1978(.a(s_204), .O(gate220inter3));
  inv1  gate1979(.a(s_205), .O(gate220inter4));
  nand2 gate1980(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate1981(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate1982(.a(G637), .O(gate220inter7));
  inv1  gate1983(.a(G681), .O(gate220inter8));
  nand2 gate1984(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate1985(.a(s_205), .b(gate220inter3), .O(gate220inter10));
  nor2  gate1986(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate1987(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate1988(.a(gate220inter12), .b(gate220inter1), .O(G701));
nand2 gate221( .a(G622), .b(G684), .O(G702) );

  xor2  gate631(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate632(.a(gate222inter0), .b(s_12), .O(gate222inter1));
  and2  gate633(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate634(.a(s_12), .O(gate222inter3));
  inv1  gate635(.a(s_13), .O(gate222inter4));
  nand2 gate636(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate637(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate638(.a(G632), .O(gate222inter7));
  inv1  gate639(.a(G684), .O(gate222inter8));
  nand2 gate640(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate641(.a(s_13), .b(gate222inter3), .O(gate222inter10));
  nor2  gate642(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate643(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate644(.a(gate222inter12), .b(gate222inter1), .O(G703));

  xor2  gate2003(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate2004(.a(gate223inter0), .b(s_208), .O(gate223inter1));
  and2  gate2005(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate2006(.a(s_208), .O(gate223inter3));
  inv1  gate2007(.a(s_209), .O(gate223inter4));
  nand2 gate2008(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate2009(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate2010(.a(G627), .O(gate223inter7));
  inv1  gate2011(.a(G687), .O(gate223inter8));
  nand2 gate2012(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate2013(.a(s_209), .b(gate223inter3), .O(gate223inter10));
  nor2  gate2014(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate2015(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate2016(.a(gate223inter12), .b(gate223inter1), .O(G704));

  xor2  gate1331(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate1332(.a(gate224inter0), .b(s_112), .O(gate224inter1));
  and2  gate1333(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate1334(.a(s_112), .O(gate224inter3));
  inv1  gate1335(.a(s_113), .O(gate224inter4));
  nand2 gate1336(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate1337(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate1338(.a(G637), .O(gate224inter7));
  inv1  gate1339(.a(G687), .O(gate224inter8));
  nand2 gate1340(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate1341(.a(s_113), .b(gate224inter3), .O(gate224inter10));
  nor2  gate1342(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate1343(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate1344(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate2353(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate2354(.a(gate227inter0), .b(s_258), .O(gate227inter1));
  and2  gate2355(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate2356(.a(s_258), .O(gate227inter3));
  inv1  gate2357(.a(s_259), .O(gate227inter4));
  nand2 gate2358(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate2359(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate2360(.a(G694), .O(gate227inter7));
  inv1  gate2361(.a(G695), .O(gate227inter8));
  nand2 gate2362(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate2363(.a(s_259), .b(gate227inter3), .O(gate227inter10));
  nor2  gate2364(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate2365(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate2366(.a(gate227inter12), .b(gate227inter1), .O(G712));
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate2899(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate2900(.a(gate233inter0), .b(s_336), .O(gate233inter1));
  and2  gate2901(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate2902(.a(s_336), .O(gate233inter3));
  inv1  gate2903(.a(s_337), .O(gate233inter4));
  nand2 gate2904(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate2905(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate2906(.a(G242), .O(gate233inter7));
  inv1  gate2907(.a(G718), .O(gate233inter8));
  nand2 gate2908(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate2909(.a(s_337), .b(gate233inter3), .O(gate233inter10));
  nor2  gate2910(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate2911(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate2912(.a(gate233inter12), .b(gate233inter1), .O(G730));

  xor2  gate1723(.a(G721), .b(G245), .O(gate234inter0));
  nand2 gate1724(.a(gate234inter0), .b(s_168), .O(gate234inter1));
  and2  gate1725(.a(G721), .b(G245), .O(gate234inter2));
  inv1  gate1726(.a(s_168), .O(gate234inter3));
  inv1  gate1727(.a(s_169), .O(gate234inter4));
  nand2 gate1728(.a(gate234inter4), .b(gate234inter3), .O(gate234inter5));
  nor2  gate1729(.a(gate234inter5), .b(gate234inter2), .O(gate234inter6));
  inv1  gate1730(.a(G245), .O(gate234inter7));
  inv1  gate1731(.a(G721), .O(gate234inter8));
  nand2 gate1732(.a(gate234inter8), .b(gate234inter7), .O(gate234inter9));
  nand2 gate1733(.a(s_169), .b(gate234inter3), .O(gate234inter10));
  nor2  gate1734(.a(gate234inter10), .b(gate234inter9), .O(gate234inter11));
  nor2  gate1735(.a(gate234inter11), .b(gate234inter6), .O(gate234inter12));
  nand2 gate1736(.a(gate234inter12), .b(gate234inter1), .O(G733));
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate1499(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate1500(.a(gate236inter0), .b(s_136), .O(gate236inter1));
  and2  gate1501(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate1502(.a(s_136), .O(gate236inter3));
  inv1  gate1503(.a(s_137), .O(gate236inter4));
  nand2 gate1504(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate1505(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate1506(.a(G251), .O(gate236inter7));
  inv1  gate1507(.a(G727), .O(gate236inter8));
  nand2 gate1508(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate1509(.a(s_137), .b(gate236inter3), .O(gate236inter10));
  nor2  gate1510(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate1511(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate1512(.a(gate236inter12), .b(gate236inter1), .O(G739));

  xor2  gate1233(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate1234(.a(gate237inter0), .b(s_98), .O(gate237inter1));
  and2  gate1235(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate1236(.a(s_98), .O(gate237inter3));
  inv1  gate1237(.a(s_99), .O(gate237inter4));
  nand2 gate1238(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1239(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1240(.a(G254), .O(gate237inter7));
  inv1  gate1241(.a(G706), .O(gate237inter8));
  nand2 gate1242(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1243(.a(s_99), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1244(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1245(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1246(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );

  xor2  gate2129(.a(G712), .b(G260), .O(gate239inter0));
  nand2 gate2130(.a(gate239inter0), .b(s_226), .O(gate239inter1));
  and2  gate2131(.a(G712), .b(G260), .O(gate239inter2));
  inv1  gate2132(.a(s_226), .O(gate239inter3));
  inv1  gate2133(.a(s_227), .O(gate239inter4));
  nand2 gate2134(.a(gate239inter4), .b(gate239inter3), .O(gate239inter5));
  nor2  gate2135(.a(gate239inter5), .b(gate239inter2), .O(gate239inter6));
  inv1  gate2136(.a(G260), .O(gate239inter7));
  inv1  gate2137(.a(G712), .O(gate239inter8));
  nand2 gate2138(.a(gate239inter8), .b(gate239inter7), .O(gate239inter9));
  nand2 gate2139(.a(s_227), .b(gate239inter3), .O(gate239inter10));
  nor2  gate2140(.a(gate239inter10), .b(gate239inter9), .O(gate239inter11));
  nor2  gate2141(.a(gate239inter11), .b(gate239inter6), .O(gate239inter12));
  nand2 gate2142(.a(gate239inter12), .b(gate239inter1), .O(G748));
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );

  xor2  gate1891(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1892(.a(gate243inter0), .b(s_192), .O(gate243inter1));
  and2  gate1893(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1894(.a(s_192), .O(gate243inter3));
  inv1  gate1895(.a(s_193), .O(gate243inter4));
  nand2 gate1896(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1897(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1898(.a(G245), .O(gate243inter7));
  inv1  gate1899(.a(G733), .O(gate243inter8));
  nand2 gate1900(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1901(.a(s_193), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1902(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1903(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1904(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );

  xor2  gate2171(.a(G736), .b(G248), .O(gate245inter0));
  nand2 gate2172(.a(gate245inter0), .b(s_232), .O(gate245inter1));
  and2  gate2173(.a(G736), .b(G248), .O(gate245inter2));
  inv1  gate2174(.a(s_232), .O(gate245inter3));
  inv1  gate2175(.a(s_233), .O(gate245inter4));
  nand2 gate2176(.a(gate245inter4), .b(gate245inter3), .O(gate245inter5));
  nor2  gate2177(.a(gate245inter5), .b(gate245inter2), .O(gate245inter6));
  inv1  gate2178(.a(G248), .O(gate245inter7));
  inv1  gate2179(.a(G736), .O(gate245inter8));
  nand2 gate2180(.a(gate245inter8), .b(gate245inter7), .O(gate245inter9));
  nand2 gate2181(.a(s_233), .b(gate245inter3), .O(gate245inter10));
  nor2  gate2182(.a(gate245inter10), .b(gate245inter9), .O(gate245inter11));
  nor2  gate2183(.a(gate245inter11), .b(gate245inter6), .O(gate245inter12));
  nand2 gate2184(.a(gate245inter12), .b(gate245inter1), .O(G758));

  xor2  gate547(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate548(.a(gate246inter0), .b(s_0), .O(gate246inter1));
  and2  gate549(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate550(.a(s_0), .O(gate246inter3));
  inv1  gate551(.a(s_1), .O(gate246inter4));
  nand2 gate552(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate553(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate554(.a(G724), .O(gate246inter7));
  inv1  gate555(.a(G736), .O(gate246inter8));
  nand2 gate556(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate557(.a(s_1), .b(gate246inter3), .O(gate246inter10));
  nor2  gate558(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate559(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate560(.a(gate246inter12), .b(gate246inter1), .O(G759));

  xor2  gate1849(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate1850(.a(gate247inter0), .b(s_186), .O(gate247inter1));
  and2  gate1851(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate1852(.a(s_186), .O(gate247inter3));
  inv1  gate1853(.a(s_187), .O(gate247inter4));
  nand2 gate1854(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate1855(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate1856(.a(G251), .O(gate247inter7));
  inv1  gate1857(.a(G739), .O(gate247inter8));
  nand2 gate1858(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate1859(.a(s_187), .b(gate247inter3), .O(gate247inter10));
  nor2  gate1860(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate1861(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate1862(.a(gate247inter12), .b(gate247inter1), .O(G760));

  xor2  gate1541(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate1542(.a(gate248inter0), .b(s_142), .O(gate248inter1));
  and2  gate1543(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate1544(.a(s_142), .O(gate248inter3));
  inv1  gate1545(.a(s_143), .O(gate248inter4));
  nand2 gate1546(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate1547(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate1548(.a(G727), .O(gate248inter7));
  inv1  gate1549(.a(G739), .O(gate248inter8));
  nand2 gate1550(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate1551(.a(s_143), .b(gate248inter3), .O(gate248inter10));
  nor2  gate1552(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate1553(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate1554(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );

  xor2  gate1359(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate1360(.a(gate251inter0), .b(s_116), .O(gate251inter1));
  and2  gate1361(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate1362(.a(s_116), .O(gate251inter3));
  inv1  gate1363(.a(s_117), .O(gate251inter4));
  nand2 gate1364(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate1365(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate1366(.a(G257), .O(gate251inter7));
  inv1  gate1367(.a(G745), .O(gate251inter8));
  nand2 gate1368(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate1369(.a(s_117), .b(gate251inter3), .O(gate251inter10));
  nor2  gate1370(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate1371(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate1372(.a(gate251inter12), .b(gate251inter1), .O(G764));
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate2297(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate2298(.a(gate253inter0), .b(s_250), .O(gate253inter1));
  and2  gate2299(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate2300(.a(s_250), .O(gate253inter3));
  inv1  gate2301(.a(s_251), .O(gate253inter4));
  nand2 gate2302(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate2303(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate2304(.a(G260), .O(gate253inter7));
  inv1  gate2305(.a(G748), .O(gate253inter8));
  nand2 gate2306(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate2307(.a(s_251), .b(gate253inter3), .O(gate253inter10));
  nor2  gate2308(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate2309(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate2310(.a(gate253inter12), .b(gate253inter1), .O(G766));

  xor2  gate855(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate856(.a(gate254inter0), .b(s_44), .O(gate254inter1));
  and2  gate857(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate858(.a(s_44), .O(gate254inter3));
  inv1  gate859(.a(s_45), .O(gate254inter4));
  nand2 gate860(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate861(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate862(.a(G712), .O(gate254inter7));
  inv1  gate863(.a(G748), .O(gate254inter8));
  nand2 gate864(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate865(.a(s_45), .b(gate254inter3), .O(gate254inter10));
  nor2  gate866(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate867(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate868(.a(gate254inter12), .b(gate254inter1), .O(G767));
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate2927(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate2928(.a(gate258inter0), .b(s_340), .O(gate258inter1));
  and2  gate2929(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate2930(.a(s_340), .O(gate258inter3));
  inv1  gate2931(.a(s_341), .O(gate258inter4));
  nand2 gate2932(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate2933(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate2934(.a(G756), .O(gate258inter7));
  inv1  gate2935(.a(G757), .O(gate258inter8));
  nand2 gate2936(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate2937(.a(s_341), .b(gate258inter3), .O(gate258inter10));
  nor2  gate2938(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate2939(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate2940(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );

  xor2  gate2367(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate2368(.a(gate261inter0), .b(s_260), .O(gate261inter1));
  and2  gate2369(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate2370(.a(s_260), .O(gate261inter3));
  inv1  gate2371(.a(s_261), .O(gate261inter4));
  nand2 gate2372(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate2373(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate2374(.a(G762), .O(gate261inter7));
  inv1  gate2375(.a(G763), .O(gate261inter8));
  nand2 gate2376(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate2377(.a(s_261), .b(gate261inter3), .O(gate261inter10));
  nor2  gate2378(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate2379(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate2380(.a(gate261inter12), .b(gate261inter1), .O(G782));

  xor2  gate827(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate828(.a(gate262inter0), .b(s_40), .O(gate262inter1));
  and2  gate829(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate830(.a(s_40), .O(gate262inter3));
  inv1  gate831(.a(s_41), .O(gate262inter4));
  nand2 gate832(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate833(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate834(.a(G764), .O(gate262inter7));
  inv1  gate835(.a(G765), .O(gate262inter8));
  nand2 gate836(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate837(.a(s_41), .b(gate262inter3), .O(gate262inter10));
  nor2  gate838(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate839(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate840(.a(gate262inter12), .b(gate262inter1), .O(G785));

  xor2  gate743(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate744(.a(gate263inter0), .b(s_28), .O(gate263inter1));
  and2  gate745(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate746(.a(s_28), .O(gate263inter3));
  inv1  gate747(.a(s_29), .O(gate263inter4));
  nand2 gate748(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate749(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate750(.a(G766), .O(gate263inter7));
  inv1  gate751(.a(G767), .O(gate263inter8));
  nand2 gate752(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate753(.a(s_29), .b(gate263inter3), .O(gate263inter10));
  nor2  gate754(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate755(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate756(.a(gate263inter12), .b(gate263inter1), .O(G788));

  xor2  gate981(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate982(.a(gate264inter0), .b(s_62), .O(gate264inter1));
  and2  gate983(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate984(.a(s_62), .O(gate264inter3));
  inv1  gate985(.a(s_63), .O(gate264inter4));
  nand2 gate986(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate987(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate988(.a(G768), .O(gate264inter7));
  inv1  gate989(.a(G769), .O(gate264inter8));
  nand2 gate990(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate991(.a(s_63), .b(gate264inter3), .O(gate264inter10));
  nor2  gate992(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate993(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate994(.a(gate264inter12), .b(gate264inter1), .O(G791));

  xor2  gate1835(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate1836(.a(gate265inter0), .b(s_184), .O(gate265inter1));
  and2  gate1837(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate1838(.a(s_184), .O(gate265inter3));
  inv1  gate1839(.a(s_185), .O(gate265inter4));
  nand2 gate1840(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate1841(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate1842(.a(G642), .O(gate265inter7));
  inv1  gate1843(.a(G770), .O(gate265inter8));
  nand2 gate1844(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate1845(.a(s_185), .b(gate265inter3), .O(gate265inter10));
  nor2  gate1846(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate1847(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate1848(.a(gate265inter12), .b(gate265inter1), .O(G794));
nand2 gate266( .a(G645), .b(G773), .O(G797) );

  xor2  gate1289(.a(G776), .b(G648), .O(gate267inter0));
  nand2 gate1290(.a(gate267inter0), .b(s_106), .O(gate267inter1));
  and2  gate1291(.a(G776), .b(G648), .O(gate267inter2));
  inv1  gate1292(.a(s_106), .O(gate267inter3));
  inv1  gate1293(.a(s_107), .O(gate267inter4));
  nand2 gate1294(.a(gate267inter4), .b(gate267inter3), .O(gate267inter5));
  nor2  gate1295(.a(gate267inter5), .b(gate267inter2), .O(gate267inter6));
  inv1  gate1296(.a(G648), .O(gate267inter7));
  inv1  gate1297(.a(G776), .O(gate267inter8));
  nand2 gate1298(.a(gate267inter8), .b(gate267inter7), .O(gate267inter9));
  nand2 gate1299(.a(s_107), .b(gate267inter3), .O(gate267inter10));
  nor2  gate1300(.a(gate267inter10), .b(gate267inter9), .O(gate267inter11));
  nor2  gate1301(.a(gate267inter11), .b(gate267inter6), .O(gate267inter12));
  nand2 gate1302(.a(gate267inter12), .b(gate267inter1), .O(G800));
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );

  xor2  gate2493(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate2494(.a(gate271inter0), .b(s_278), .O(gate271inter1));
  and2  gate2495(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate2496(.a(s_278), .O(gate271inter3));
  inv1  gate2497(.a(s_279), .O(gate271inter4));
  nand2 gate2498(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate2499(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate2500(.a(G660), .O(gate271inter7));
  inv1  gate2501(.a(G788), .O(gate271inter8));
  nand2 gate2502(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate2503(.a(s_279), .b(gate271inter3), .O(gate271inter10));
  nor2  gate2504(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate2505(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate2506(.a(gate271inter12), .b(gate271inter1), .O(G812));

  xor2  gate1527(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate1528(.a(gate272inter0), .b(s_140), .O(gate272inter1));
  and2  gate1529(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate1530(.a(s_140), .O(gate272inter3));
  inv1  gate1531(.a(s_141), .O(gate272inter4));
  nand2 gate1532(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate1533(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate1534(.a(G663), .O(gate272inter7));
  inv1  gate1535(.a(G791), .O(gate272inter8));
  nand2 gate1536(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate1537(.a(s_141), .b(gate272inter3), .O(gate272inter10));
  nor2  gate1538(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate1539(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate1540(.a(gate272inter12), .b(gate272inter1), .O(G815));

  xor2  gate1303(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate1304(.a(gate273inter0), .b(s_108), .O(gate273inter1));
  and2  gate1305(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate1306(.a(s_108), .O(gate273inter3));
  inv1  gate1307(.a(s_109), .O(gate273inter4));
  nand2 gate1308(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate1309(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate1310(.a(G642), .O(gate273inter7));
  inv1  gate1311(.a(G794), .O(gate273inter8));
  nand2 gate1312(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate1313(.a(s_109), .b(gate273inter3), .O(gate273inter10));
  nor2  gate1314(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate1315(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate1316(.a(gate273inter12), .b(gate273inter1), .O(G818));
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );

  xor2  gate1569(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate1570(.a(gate277inter0), .b(s_146), .O(gate277inter1));
  and2  gate1571(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate1572(.a(s_146), .O(gate277inter3));
  inv1  gate1573(.a(s_147), .O(gate277inter4));
  nand2 gate1574(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate1575(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate1576(.a(G648), .O(gate277inter7));
  inv1  gate1577(.a(G800), .O(gate277inter8));
  nand2 gate1578(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate1579(.a(s_147), .b(gate277inter3), .O(gate277inter10));
  nor2  gate1580(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate1581(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate1582(.a(gate277inter12), .b(gate277inter1), .O(G822));
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );

  xor2  gate1471(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate1472(.a(gate281inter0), .b(s_132), .O(gate281inter1));
  and2  gate1473(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate1474(.a(s_132), .O(gate281inter3));
  inv1  gate1475(.a(s_133), .O(gate281inter4));
  nand2 gate1476(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate1477(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate1478(.a(G654), .O(gate281inter7));
  inv1  gate1479(.a(G806), .O(gate281inter8));
  nand2 gate1480(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate1481(.a(s_133), .b(gate281inter3), .O(gate281inter10));
  nor2  gate1482(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate1483(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate1484(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );

  xor2  gate2311(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate2312(.a(gate284inter0), .b(s_252), .O(gate284inter1));
  and2  gate2313(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate2314(.a(s_252), .O(gate284inter3));
  inv1  gate2315(.a(s_253), .O(gate284inter4));
  nand2 gate2316(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate2317(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate2318(.a(G785), .O(gate284inter7));
  inv1  gate2319(.a(G809), .O(gate284inter8));
  nand2 gate2320(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate2321(.a(s_253), .b(gate284inter3), .O(gate284inter10));
  nor2  gate2322(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate2323(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate2324(.a(gate284inter12), .b(gate284inter1), .O(G829));

  xor2  gate1779(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate1780(.a(gate285inter0), .b(s_176), .O(gate285inter1));
  and2  gate1781(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate1782(.a(s_176), .O(gate285inter3));
  inv1  gate1783(.a(s_177), .O(gate285inter4));
  nand2 gate1784(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate1785(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate1786(.a(G660), .O(gate285inter7));
  inv1  gate1787(.a(G812), .O(gate285inter8));
  nand2 gate1788(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate1789(.a(s_177), .b(gate285inter3), .O(gate285inter10));
  nor2  gate1790(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate1791(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate1792(.a(gate285inter12), .b(gate285inter1), .O(G830));

  xor2  gate799(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate800(.a(gate286inter0), .b(s_36), .O(gate286inter1));
  and2  gate801(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate802(.a(s_36), .O(gate286inter3));
  inv1  gate803(.a(s_37), .O(gate286inter4));
  nand2 gate804(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate805(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate806(.a(G788), .O(gate286inter7));
  inv1  gate807(.a(G812), .O(gate286inter8));
  nand2 gate808(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate809(.a(s_37), .b(gate286inter3), .O(gate286inter10));
  nor2  gate810(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate811(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate812(.a(gate286inter12), .b(gate286inter1), .O(G831));

  xor2  gate2535(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate2536(.a(gate287inter0), .b(s_284), .O(gate287inter1));
  and2  gate2537(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate2538(.a(s_284), .O(gate287inter3));
  inv1  gate2539(.a(s_285), .O(gate287inter4));
  nand2 gate2540(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate2541(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate2542(.a(G663), .O(gate287inter7));
  inv1  gate2543(.a(G815), .O(gate287inter8));
  nand2 gate2544(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate2545(.a(s_285), .b(gate287inter3), .O(gate287inter10));
  nor2  gate2546(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate2547(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate2548(.a(gate287inter12), .b(gate287inter1), .O(G832));

  xor2  gate2857(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate2858(.a(gate288inter0), .b(s_330), .O(gate288inter1));
  and2  gate2859(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate2860(.a(s_330), .O(gate288inter3));
  inv1  gate2861(.a(s_331), .O(gate288inter4));
  nand2 gate2862(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate2863(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate2864(.a(G791), .O(gate288inter7));
  inv1  gate2865(.a(G815), .O(gate288inter8));
  nand2 gate2866(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate2867(.a(s_331), .b(gate288inter3), .O(gate288inter10));
  nor2  gate2868(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate2869(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate2870(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate2941(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate2942(.a(gate292inter0), .b(s_342), .O(gate292inter1));
  and2  gate2943(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate2944(.a(s_342), .O(gate292inter3));
  inv1  gate2945(.a(s_343), .O(gate292inter4));
  nand2 gate2946(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate2947(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate2948(.a(G824), .O(gate292inter7));
  inv1  gate2949(.a(G825), .O(gate292inter8));
  nand2 gate2950(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate2951(.a(s_343), .b(gate292inter3), .O(gate292inter10));
  nor2  gate2952(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate2953(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate2954(.a(gate292inter12), .b(gate292inter1), .O(G873));

  xor2  gate715(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate716(.a(gate293inter0), .b(s_24), .O(gate293inter1));
  and2  gate717(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate718(.a(s_24), .O(gate293inter3));
  inv1  gate719(.a(s_25), .O(gate293inter4));
  nand2 gate720(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate721(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate722(.a(G828), .O(gate293inter7));
  inv1  gate723(.a(G829), .O(gate293inter8));
  nand2 gate724(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate725(.a(s_25), .b(gate293inter3), .O(gate293inter10));
  nor2  gate726(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate727(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate728(.a(gate293inter12), .b(gate293inter1), .O(G886));

  xor2  gate953(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate954(.a(gate294inter0), .b(s_58), .O(gate294inter1));
  and2  gate955(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate956(.a(s_58), .O(gate294inter3));
  inv1  gate957(.a(s_59), .O(gate294inter4));
  nand2 gate958(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate959(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate960(.a(G832), .O(gate294inter7));
  inv1  gate961(.a(G833), .O(gate294inter8));
  nand2 gate962(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate963(.a(s_59), .b(gate294inter3), .O(gate294inter10));
  nor2  gate964(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate965(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate966(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate1317(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate1318(.a(gate393inter0), .b(s_110), .O(gate393inter1));
  and2  gate1319(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate1320(.a(s_110), .O(gate393inter3));
  inv1  gate1321(.a(s_111), .O(gate393inter4));
  nand2 gate1322(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate1323(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate1324(.a(G7), .O(gate393inter7));
  inv1  gate1325(.a(G1054), .O(gate393inter8));
  nand2 gate1326(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate1327(.a(s_111), .b(gate393inter3), .O(gate393inter10));
  nor2  gate1328(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate1329(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate1330(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );

  xor2  gate2031(.a(G1069), .b(G12), .O(gate398inter0));
  nand2 gate2032(.a(gate398inter0), .b(s_212), .O(gate398inter1));
  and2  gate2033(.a(G1069), .b(G12), .O(gate398inter2));
  inv1  gate2034(.a(s_212), .O(gate398inter3));
  inv1  gate2035(.a(s_213), .O(gate398inter4));
  nand2 gate2036(.a(gate398inter4), .b(gate398inter3), .O(gate398inter5));
  nor2  gate2037(.a(gate398inter5), .b(gate398inter2), .O(gate398inter6));
  inv1  gate2038(.a(G12), .O(gate398inter7));
  inv1  gate2039(.a(G1069), .O(gate398inter8));
  nand2 gate2040(.a(gate398inter8), .b(gate398inter7), .O(gate398inter9));
  nand2 gate2041(.a(s_213), .b(gate398inter3), .O(gate398inter10));
  nor2  gate2042(.a(gate398inter10), .b(gate398inter9), .O(gate398inter11));
  nor2  gate2043(.a(gate398inter11), .b(gate398inter6), .O(gate398inter12));
  nand2 gate2044(.a(gate398inter12), .b(gate398inter1), .O(G1165));

  xor2  gate2661(.a(G1072), .b(G13), .O(gate399inter0));
  nand2 gate2662(.a(gate399inter0), .b(s_302), .O(gate399inter1));
  and2  gate2663(.a(G1072), .b(G13), .O(gate399inter2));
  inv1  gate2664(.a(s_302), .O(gate399inter3));
  inv1  gate2665(.a(s_303), .O(gate399inter4));
  nand2 gate2666(.a(gate399inter4), .b(gate399inter3), .O(gate399inter5));
  nor2  gate2667(.a(gate399inter5), .b(gate399inter2), .O(gate399inter6));
  inv1  gate2668(.a(G13), .O(gate399inter7));
  inv1  gate2669(.a(G1072), .O(gate399inter8));
  nand2 gate2670(.a(gate399inter8), .b(gate399inter7), .O(gate399inter9));
  nand2 gate2671(.a(s_303), .b(gate399inter3), .O(gate399inter10));
  nor2  gate2672(.a(gate399inter10), .b(gate399inter9), .O(gate399inter11));
  nor2  gate2673(.a(gate399inter11), .b(gate399inter6), .O(gate399inter12));
  nand2 gate2674(.a(gate399inter12), .b(gate399inter1), .O(G1168));
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );

  xor2  gate2283(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate2284(.a(gate401inter0), .b(s_248), .O(gate401inter1));
  and2  gate2285(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate2286(.a(s_248), .O(gate401inter3));
  inv1  gate2287(.a(s_249), .O(gate401inter4));
  nand2 gate2288(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate2289(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate2290(.a(G15), .O(gate401inter7));
  inv1  gate2291(.a(G1078), .O(gate401inter8));
  nand2 gate2292(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate2293(.a(s_249), .b(gate401inter3), .O(gate401inter10));
  nor2  gate2294(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate2295(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate2296(.a(gate401inter12), .b(gate401inter1), .O(G1174));
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate2255(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate2256(.a(gate403inter0), .b(s_244), .O(gate403inter1));
  and2  gate2257(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate2258(.a(s_244), .O(gate403inter3));
  inv1  gate2259(.a(s_245), .O(gate403inter4));
  nand2 gate2260(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate2261(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate2262(.a(G17), .O(gate403inter7));
  inv1  gate2263(.a(G1084), .O(gate403inter8));
  nand2 gate2264(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate2265(.a(s_245), .b(gate403inter3), .O(gate403inter10));
  nor2  gate2266(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate2267(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate2268(.a(gate403inter12), .b(gate403inter1), .O(G1180));
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );

  xor2  gate561(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate562(.a(gate410inter0), .b(s_2), .O(gate410inter1));
  and2  gate563(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate564(.a(s_2), .O(gate410inter3));
  inv1  gate565(.a(s_3), .O(gate410inter4));
  nand2 gate566(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate567(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate568(.a(G24), .O(gate410inter7));
  inv1  gate569(.a(G1105), .O(gate410inter8));
  nand2 gate570(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate571(.a(s_3), .b(gate410inter3), .O(gate410inter10));
  nor2  gate572(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate573(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate574(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate995(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate996(.a(gate415inter0), .b(s_64), .O(gate415inter1));
  and2  gate997(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate998(.a(s_64), .O(gate415inter3));
  inv1  gate999(.a(s_65), .O(gate415inter4));
  nand2 gate1000(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate1001(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate1002(.a(G29), .O(gate415inter7));
  inv1  gate1003(.a(G1120), .O(gate415inter8));
  nand2 gate1004(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate1005(.a(s_65), .b(gate415inter3), .O(gate415inter10));
  nor2  gate1006(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate1007(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate1008(.a(gate415inter12), .b(gate415inter1), .O(G1216));

  xor2  gate1037(.a(G1123), .b(G30), .O(gate416inter0));
  nand2 gate1038(.a(gate416inter0), .b(s_70), .O(gate416inter1));
  and2  gate1039(.a(G1123), .b(G30), .O(gate416inter2));
  inv1  gate1040(.a(s_70), .O(gate416inter3));
  inv1  gate1041(.a(s_71), .O(gate416inter4));
  nand2 gate1042(.a(gate416inter4), .b(gate416inter3), .O(gate416inter5));
  nor2  gate1043(.a(gate416inter5), .b(gate416inter2), .O(gate416inter6));
  inv1  gate1044(.a(G30), .O(gate416inter7));
  inv1  gate1045(.a(G1123), .O(gate416inter8));
  nand2 gate1046(.a(gate416inter8), .b(gate416inter7), .O(gate416inter9));
  nand2 gate1047(.a(s_71), .b(gate416inter3), .O(gate416inter10));
  nor2  gate1048(.a(gate416inter10), .b(gate416inter9), .O(gate416inter11));
  nor2  gate1049(.a(gate416inter11), .b(gate416inter6), .O(gate416inter12));
  nand2 gate1050(.a(gate416inter12), .b(gate416inter1), .O(G1219));

  xor2  gate2913(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate2914(.a(gate417inter0), .b(s_338), .O(gate417inter1));
  and2  gate2915(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate2916(.a(s_338), .O(gate417inter3));
  inv1  gate2917(.a(s_339), .O(gate417inter4));
  nand2 gate2918(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate2919(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate2920(.a(G31), .O(gate417inter7));
  inv1  gate2921(.a(G1126), .O(gate417inter8));
  nand2 gate2922(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate2923(.a(s_339), .b(gate417inter3), .O(gate417inter10));
  nor2  gate2924(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate2925(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate2926(.a(gate417inter12), .b(gate417inter1), .O(G1222));

  xor2  gate2885(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate2886(.a(gate418inter0), .b(s_334), .O(gate418inter1));
  and2  gate2887(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate2888(.a(s_334), .O(gate418inter3));
  inv1  gate2889(.a(s_335), .O(gate418inter4));
  nand2 gate2890(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate2891(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate2892(.a(G32), .O(gate418inter7));
  inv1  gate2893(.a(G1129), .O(gate418inter8));
  nand2 gate2894(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate2895(.a(s_335), .b(gate418inter3), .O(gate418inter10));
  nor2  gate2896(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate2897(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate2898(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate1583(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate1584(.a(gate422inter0), .b(s_148), .O(gate422inter1));
  and2  gate1585(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate1586(.a(s_148), .O(gate422inter3));
  inv1  gate1587(.a(s_149), .O(gate422inter4));
  nand2 gate1588(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate1589(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate1590(.a(G1039), .O(gate422inter7));
  inv1  gate1591(.a(G1135), .O(gate422inter8));
  nand2 gate1592(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate1593(.a(s_149), .b(gate422inter3), .O(gate422inter10));
  nor2  gate1594(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate1595(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate1596(.a(gate422inter12), .b(gate422inter1), .O(G1231));

  xor2  gate1065(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate1066(.a(gate423inter0), .b(s_74), .O(gate423inter1));
  and2  gate1067(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate1068(.a(s_74), .O(gate423inter3));
  inv1  gate1069(.a(s_75), .O(gate423inter4));
  nand2 gate1070(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate1071(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate1072(.a(G3), .O(gate423inter7));
  inv1  gate1073(.a(G1138), .O(gate423inter8));
  nand2 gate1074(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate1075(.a(s_75), .b(gate423inter3), .O(gate423inter10));
  nor2  gate1076(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate1077(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate1078(.a(gate423inter12), .b(gate423inter1), .O(G1232));

  xor2  gate1667(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate1668(.a(gate424inter0), .b(s_160), .O(gate424inter1));
  and2  gate1669(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate1670(.a(s_160), .O(gate424inter3));
  inv1  gate1671(.a(s_161), .O(gate424inter4));
  nand2 gate1672(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate1673(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate1674(.a(G1042), .O(gate424inter7));
  inv1  gate1675(.a(G1138), .O(gate424inter8));
  nand2 gate1676(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate1677(.a(s_161), .b(gate424inter3), .O(gate424inter10));
  nor2  gate1678(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate1679(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate1680(.a(gate424inter12), .b(gate424inter1), .O(G1233));

  xor2  gate1597(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate1598(.a(gate425inter0), .b(s_150), .O(gate425inter1));
  and2  gate1599(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate1600(.a(s_150), .O(gate425inter3));
  inv1  gate1601(.a(s_151), .O(gate425inter4));
  nand2 gate1602(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate1603(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate1604(.a(G4), .O(gate425inter7));
  inv1  gate1605(.a(G1141), .O(gate425inter8));
  nand2 gate1606(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate1607(.a(s_151), .b(gate425inter3), .O(gate425inter10));
  nor2  gate1608(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate1609(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate1610(.a(gate425inter12), .b(gate425inter1), .O(G1234));
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate2213(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate2214(.a(gate430inter0), .b(s_238), .O(gate430inter1));
  and2  gate2215(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate2216(.a(s_238), .O(gate430inter3));
  inv1  gate2217(.a(s_239), .O(gate430inter4));
  nand2 gate2218(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate2219(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate2220(.a(G1051), .O(gate430inter7));
  inv1  gate2221(.a(G1147), .O(gate430inter8));
  nand2 gate2222(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate2223(.a(s_239), .b(gate430inter3), .O(gate430inter10));
  nor2  gate2224(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate2225(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate2226(.a(gate430inter12), .b(gate430inter1), .O(G1239));

  xor2  gate2101(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate2102(.a(gate431inter0), .b(s_222), .O(gate431inter1));
  and2  gate2103(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate2104(.a(s_222), .O(gate431inter3));
  inv1  gate2105(.a(s_223), .O(gate431inter4));
  nand2 gate2106(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate2107(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate2108(.a(G7), .O(gate431inter7));
  inv1  gate2109(.a(G1150), .O(gate431inter8));
  nand2 gate2110(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate2111(.a(s_223), .b(gate431inter3), .O(gate431inter10));
  nor2  gate2112(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate2113(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate2114(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate785(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate786(.a(gate433inter0), .b(s_34), .O(gate433inter1));
  and2  gate787(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate788(.a(s_34), .O(gate433inter3));
  inv1  gate789(.a(s_35), .O(gate433inter4));
  nand2 gate790(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate791(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate792(.a(G8), .O(gate433inter7));
  inv1  gate793(.a(G1153), .O(gate433inter8));
  nand2 gate794(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate795(.a(s_35), .b(gate433inter3), .O(gate433inter10));
  nor2  gate796(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate797(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate798(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate2437(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate2438(.a(gate435inter0), .b(s_270), .O(gate435inter1));
  and2  gate2439(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate2440(.a(s_270), .O(gate435inter3));
  inv1  gate2441(.a(s_271), .O(gate435inter4));
  nand2 gate2442(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate2443(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate2444(.a(G9), .O(gate435inter7));
  inv1  gate2445(.a(G1156), .O(gate435inter8));
  nand2 gate2446(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate2447(.a(s_271), .b(gate435inter3), .O(gate435inter10));
  nor2  gate2448(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate2449(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate2450(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate1653(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate1654(.a(gate439inter0), .b(s_158), .O(gate439inter1));
  and2  gate1655(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate1656(.a(s_158), .O(gate439inter3));
  inv1  gate1657(.a(s_159), .O(gate439inter4));
  nand2 gate1658(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate1659(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate1660(.a(G11), .O(gate439inter7));
  inv1  gate1661(.a(G1162), .O(gate439inter8));
  nand2 gate1662(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate1663(.a(s_159), .b(gate439inter3), .O(gate439inter10));
  nor2  gate1664(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate1665(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate1666(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate2829(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate2830(.a(gate442inter0), .b(s_326), .O(gate442inter1));
  and2  gate2831(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate2832(.a(s_326), .O(gate442inter3));
  inv1  gate2833(.a(s_327), .O(gate442inter4));
  nand2 gate2834(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate2835(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate2836(.a(G1069), .O(gate442inter7));
  inv1  gate2837(.a(G1165), .O(gate442inter8));
  nand2 gate2838(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate2839(.a(s_327), .b(gate442inter3), .O(gate442inter10));
  nor2  gate2840(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate2841(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate2842(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );

  xor2  gate2087(.a(G1174), .b(G1078), .O(gate448inter0));
  nand2 gate2088(.a(gate448inter0), .b(s_220), .O(gate448inter1));
  and2  gate2089(.a(G1174), .b(G1078), .O(gate448inter2));
  inv1  gate2090(.a(s_220), .O(gate448inter3));
  inv1  gate2091(.a(s_221), .O(gate448inter4));
  nand2 gate2092(.a(gate448inter4), .b(gate448inter3), .O(gate448inter5));
  nor2  gate2093(.a(gate448inter5), .b(gate448inter2), .O(gate448inter6));
  inv1  gate2094(.a(G1078), .O(gate448inter7));
  inv1  gate2095(.a(G1174), .O(gate448inter8));
  nand2 gate2096(.a(gate448inter8), .b(gate448inter7), .O(gate448inter9));
  nand2 gate2097(.a(s_221), .b(gate448inter3), .O(gate448inter10));
  nor2  gate2098(.a(gate448inter10), .b(gate448inter9), .O(gate448inter11));
  nor2  gate2099(.a(gate448inter11), .b(gate448inter6), .O(gate448inter12));
  nand2 gate2100(.a(gate448inter12), .b(gate448inter1), .O(G1257));
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );

  xor2  gate1919(.a(G1177), .b(G1081), .O(gate450inter0));
  nand2 gate1920(.a(gate450inter0), .b(s_196), .O(gate450inter1));
  and2  gate1921(.a(G1177), .b(G1081), .O(gate450inter2));
  inv1  gate1922(.a(s_196), .O(gate450inter3));
  inv1  gate1923(.a(s_197), .O(gate450inter4));
  nand2 gate1924(.a(gate450inter4), .b(gate450inter3), .O(gate450inter5));
  nor2  gate1925(.a(gate450inter5), .b(gate450inter2), .O(gate450inter6));
  inv1  gate1926(.a(G1081), .O(gate450inter7));
  inv1  gate1927(.a(G1177), .O(gate450inter8));
  nand2 gate1928(.a(gate450inter8), .b(gate450inter7), .O(gate450inter9));
  nand2 gate1929(.a(s_197), .b(gate450inter3), .O(gate450inter10));
  nor2  gate1930(.a(gate450inter10), .b(gate450inter9), .O(gate450inter11));
  nor2  gate1931(.a(gate450inter11), .b(gate450inter6), .O(gate450inter12));
  nand2 gate1932(.a(gate450inter12), .b(gate450inter1), .O(G1259));

  xor2  gate2227(.a(G1180), .b(G17), .O(gate451inter0));
  nand2 gate2228(.a(gate451inter0), .b(s_240), .O(gate451inter1));
  and2  gate2229(.a(G1180), .b(G17), .O(gate451inter2));
  inv1  gate2230(.a(s_240), .O(gate451inter3));
  inv1  gate2231(.a(s_241), .O(gate451inter4));
  nand2 gate2232(.a(gate451inter4), .b(gate451inter3), .O(gate451inter5));
  nor2  gate2233(.a(gate451inter5), .b(gate451inter2), .O(gate451inter6));
  inv1  gate2234(.a(G17), .O(gate451inter7));
  inv1  gate2235(.a(G1180), .O(gate451inter8));
  nand2 gate2236(.a(gate451inter8), .b(gate451inter7), .O(gate451inter9));
  nand2 gate2237(.a(s_241), .b(gate451inter3), .O(gate451inter10));
  nor2  gate2238(.a(gate451inter10), .b(gate451inter9), .O(gate451inter11));
  nor2  gate2239(.a(gate451inter11), .b(gate451inter6), .O(gate451inter12));
  nand2 gate2240(.a(gate451inter12), .b(gate451inter1), .O(G1260));
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate1695(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate1696(.a(gate453inter0), .b(s_164), .O(gate453inter1));
  and2  gate1697(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate1698(.a(s_164), .O(gate453inter3));
  inv1  gate1699(.a(s_165), .O(gate453inter4));
  nand2 gate1700(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate1701(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate1702(.a(G18), .O(gate453inter7));
  inv1  gate1703(.a(G1183), .O(gate453inter8));
  nand2 gate1704(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate1705(.a(s_165), .b(gate453inter3), .O(gate453inter10));
  nor2  gate1706(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate1707(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate1708(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate939(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate940(.a(gate457inter0), .b(s_56), .O(gate457inter1));
  and2  gate941(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate942(.a(s_56), .O(gate457inter3));
  inv1  gate943(.a(s_57), .O(gate457inter4));
  nand2 gate944(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate945(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate946(.a(G20), .O(gate457inter7));
  inv1  gate947(.a(G1189), .O(gate457inter8));
  nand2 gate948(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate949(.a(s_57), .b(gate457inter3), .O(gate457inter10));
  nor2  gate950(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate951(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate952(.a(gate457inter12), .b(gate457inter1), .O(G1266));

  xor2  gate2073(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate2074(.a(gate458inter0), .b(s_218), .O(gate458inter1));
  and2  gate2075(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate2076(.a(s_218), .O(gate458inter3));
  inv1  gate2077(.a(s_219), .O(gate458inter4));
  nand2 gate2078(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate2079(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate2080(.a(G1093), .O(gate458inter7));
  inv1  gate2081(.a(G1189), .O(gate458inter8));
  nand2 gate2082(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate2083(.a(s_219), .b(gate458inter3), .O(gate458inter10));
  nor2  gate2084(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate2085(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate2086(.a(gate458inter12), .b(gate458inter1), .O(G1267));

  xor2  gate1373(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate1374(.a(gate459inter0), .b(s_118), .O(gate459inter1));
  and2  gate1375(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate1376(.a(s_118), .O(gate459inter3));
  inv1  gate1377(.a(s_119), .O(gate459inter4));
  nand2 gate1378(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate1379(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate1380(.a(G21), .O(gate459inter7));
  inv1  gate1381(.a(G1192), .O(gate459inter8));
  nand2 gate1382(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate1383(.a(s_119), .b(gate459inter3), .O(gate459inter10));
  nor2  gate1384(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate1385(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate1386(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate1149(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate1150(.a(gate461inter0), .b(s_86), .O(gate461inter1));
  and2  gate1151(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate1152(.a(s_86), .O(gate461inter3));
  inv1  gate1153(.a(s_87), .O(gate461inter4));
  nand2 gate1154(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate1155(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate1156(.a(G22), .O(gate461inter7));
  inv1  gate1157(.a(G1195), .O(gate461inter8));
  nand2 gate1158(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate1159(.a(s_87), .b(gate461inter3), .O(gate461inter10));
  nor2  gate1160(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate1161(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate1162(.a(gate461inter12), .b(gate461inter1), .O(G1270));

  xor2  gate575(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate576(.a(gate462inter0), .b(s_4), .O(gate462inter1));
  and2  gate577(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate578(.a(s_4), .O(gate462inter3));
  inv1  gate579(.a(s_5), .O(gate462inter4));
  nand2 gate580(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate581(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate582(.a(G1099), .O(gate462inter7));
  inv1  gate583(.a(G1195), .O(gate462inter8));
  nand2 gate584(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate585(.a(s_5), .b(gate462inter3), .O(gate462inter10));
  nor2  gate586(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate587(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate588(.a(gate462inter12), .b(gate462inter1), .O(G1271));

  xor2  gate1639(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate1640(.a(gate463inter0), .b(s_156), .O(gate463inter1));
  and2  gate1641(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate1642(.a(s_156), .O(gate463inter3));
  inv1  gate1643(.a(s_157), .O(gate463inter4));
  nand2 gate1644(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate1645(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate1646(.a(G23), .O(gate463inter7));
  inv1  gate1647(.a(G1198), .O(gate463inter8));
  nand2 gate1648(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate1649(.a(s_157), .b(gate463inter3), .O(gate463inter10));
  nor2  gate1650(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate1651(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate1652(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate1401(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate1402(.a(gate465inter0), .b(s_122), .O(gate465inter1));
  and2  gate1403(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate1404(.a(s_122), .O(gate465inter3));
  inv1  gate1405(.a(s_123), .O(gate465inter4));
  nand2 gate1406(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate1407(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate1408(.a(G24), .O(gate465inter7));
  inv1  gate1409(.a(G1201), .O(gate465inter8));
  nand2 gate1410(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate1411(.a(s_123), .b(gate465inter3), .O(gate465inter10));
  nor2  gate1412(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate1413(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate1414(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );

  xor2  gate2871(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate2872(.a(gate468inter0), .b(s_332), .O(gate468inter1));
  and2  gate2873(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate2874(.a(s_332), .O(gate468inter3));
  inv1  gate2875(.a(s_333), .O(gate468inter4));
  nand2 gate2876(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate2877(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate2878(.a(G1108), .O(gate468inter7));
  inv1  gate2879(.a(G1204), .O(gate468inter8));
  nand2 gate2880(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate2881(.a(s_333), .b(gate468inter3), .O(gate468inter10));
  nor2  gate2882(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate2883(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate2884(.a(gate468inter12), .b(gate468inter1), .O(G1277));

  xor2  gate1961(.a(G1207), .b(G26), .O(gate469inter0));
  nand2 gate1962(.a(gate469inter0), .b(s_202), .O(gate469inter1));
  and2  gate1963(.a(G1207), .b(G26), .O(gate469inter2));
  inv1  gate1964(.a(s_202), .O(gate469inter3));
  inv1  gate1965(.a(s_203), .O(gate469inter4));
  nand2 gate1966(.a(gate469inter4), .b(gate469inter3), .O(gate469inter5));
  nor2  gate1967(.a(gate469inter5), .b(gate469inter2), .O(gate469inter6));
  inv1  gate1968(.a(G26), .O(gate469inter7));
  inv1  gate1969(.a(G1207), .O(gate469inter8));
  nand2 gate1970(.a(gate469inter8), .b(gate469inter7), .O(gate469inter9));
  nand2 gate1971(.a(s_203), .b(gate469inter3), .O(gate469inter10));
  nor2  gate1972(.a(gate469inter10), .b(gate469inter9), .O(gate469inter11));
  nor2  gate1973(.a(gate469inter11), .b(gate469inter6), .O(gate469inter12));
  nand2 gate1974(.a(gate469inter12), .b(gate469inter1), .O(G1278));
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate673(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate674(.a(gate471inter0), .b(s_18), .O(gate471inter1));
  and2  gate675(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate676(.a(s_18), .O(gate471inter3));
  inv1  gate677(.a(s_19), .O(gate471inter4));
  nand2 gate678(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate679(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate680(.a(G27), .O(gate471inter7));
  inv1  gate681(.a(G1210), .O(gate471inter8));
  nand2 gate682(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate683(.a(s_19), .b(gate471inter3), .O(gate471inter10));
  nor2  gate684(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate685(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate686(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );

  xor2  gate2157(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate2158(.a(gate479inter0), .b(s_230), .O(gate479inter1));
  and2  gate2159(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate2160(.a(s_230), .O(gate479inter3));
  inv1  gate2161(.a(s_231), .O(gate479inter4));
  nand2 gate2162(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate2163(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate2164(.a(G31), .O(gate479inter7));
  inv1  gate2165(.a(G1222), .O(gate479inter8));
  nand2 gate2166(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate2167(.a(s_231), .b(gate479inter3), .O(gate479inter10));
  nor2  gate2168(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate2169(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate2170(.a(gate479inter12), .b(gate479inter1), .O(G1288));

  xor2  gate771(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate772(.a(gate480inter0), .b(s_32), .O(gate480inter1));
  and2  gate773(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate774(.a(s_32), .O(gate480inter3));
  inv1  gate775(.a(s_33), .O(gate480inter4));
  nand2 gate776(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate777(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate778(.a(G1126), .O(gate480inter7));
  inv1  gate779(.a(G1222), .O(gate480inter8));
  nand2 gate780(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate781(.a(s_33), .b(gate480inter3), .O(gate480inter10));
  nor2  gate782(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate783(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate784(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate2339(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate2340(.a(gate482inter0), .b(s_256), .O(gate482inter1));
  and2  gate2341(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate2342(.a(s_256), .O(gate482inter3));
  inv1  gate2343(.a(s_257), .O(gate482inter4));
  nand2 gate2344(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate2345(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate2346(.a(G1129), .O(gate482inter7));
  inv1  gate2347(.a(G1225), .O(gate482inter8));
  nand2 gate2348(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate2349(.a(s_257), .b(gate482inter3), .O(gate482inter10));
  nor2  gate2350(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate2351(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate2352(.a(gate482inter12), .b(gate482inter1), .O(G1291));

  xor2  gate2759(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate2760(.a(gate483inter0), .b(s_316), .O(gate483inter1));
  and2  gate2761(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate2762(.a(s_316), .O(gate483inter3));
  inv1  gate2763(.a(s_317), .O(gate483inter4));
  nand2 gate2764(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate2765(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate2766(.a(G1228), .O(gate483inter7));
  inv1  gate2767(.a(G1229), .O(gate483inter8));
  nand2 gate2768(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate2769(.a(s_317), .b(gate483inter3), .O(gate483inter10));
  nor2  gate2770(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate2771(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate2772(.a(gate483inter12), .b(gate483inter1), .O(G1292));

  xor2  gate841(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate842(.a(gate484inter0), .b(s_42), .O(gate484inter1));
  and2  gate843(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate844(.a(s_42), .O(gate484inter3));
  inv1  gate845(.a(s_43), .O(gate484inter4));
  nand2 gate846(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate847(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate848(.a(G1230), .O(gate484inter7));
  inv1  gate849(.a(G1231), .O(gate484inter8));
  nand2 gate850(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate851(.a(s_43), .b(gate484inter3), .O(gate484inter10));
  nor2  gate852(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate853(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate854(.a(gate484inter12), .b(gate484inter1), .O(G1293));

  xor2  gate2605(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate2606(.a(gate485inter0), .b(s_294), .O(gate485inter1));
  and2  gate2607(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate2608(.a(s_294), .O(gate485inter3));
  inv1  gate2609(.a(s_295), .O(gate485inter4));
  nand2 gate2610(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate2611(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate2612(.a(G1232), .O(gate485inter7));
  inv1  gate2613(.a(G1233), .O(gate485inter8));
  nand2 gate2614(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate2615(.a(s_295), .b(gate485inter3), .O(gate485inter10));
  nor2  gate2616(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate2617(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate2618(.a(gate485inter12), .b(gate485inter1), .O(G1294));

  xor2  gate1107(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate1108(.a(gate486inter0), .b(s_80), .O(gate486inter1));
  and2  gate1109(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate1110(.a(s_80), .O(gate486inter3));
  inv1  gate1111(.a(s_81), .O(gate486inter4));
  nand2 gate1112(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate1113(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate1114(.a(G1234), .O(gate486inter7));
  inv1  gate1115(.a(G1235), .O(gate486inter8));
  nand2 gate1116(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate1117(.a(s_81), .b(gate486inter3), .O(gate486inter10));
  nor2  gate1118(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate1119(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate1120(.a(gate486inter12), .b(gate486inter1), .O(G1295));

  xor2  gate2241(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate2242(.a(gate487inter0), .b(s_242), .O(gate487inter1));
  and2  gate2243(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate2244(.a(s_242), .O(gate487inter3));
  inv1  gate2245(.a(s_243), .O(gate487inter4));
  nand2 gate2246(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate2247(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate2248(.a(G1236), .O(gate487inter7));
  inv1  gate2249(.a(G1237), .O(gate487inter8));
  nand2 gate2250(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate2251(.a(s_243), .b(gate487inter3), .O(gate487inter10));
  nor2  gate2252(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate2253(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate2254(.a(gate487inter12), .b(gate487inter1), .O(G1296));

  xor2  gate2801(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate2802(.a(gate488inter0), .b(s_322), .O(gate488inter1));
  and2  gate2803(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate2804(.a(s_322), .O(gate488inter3));
  inv1  gate2805(.a(s_323), .O(gate488inter4));
  nand2 gate2806(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate2807(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate2808(.a(G1238), .O(gate488inter7));
  inv1  gate2809(.a(G1239), .O(gate488inter8));
  nand2 gate2810(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate2811(.a(s_323), .b(gate488inter3), .O(gate488inter10));
  nor2  gate2812(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate2813(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate2814(.a(gate488inter12), .b(gate488inter1), .O(G1297));
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate2969(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate2970(.a(gate490inter0), .b(s_346), .O(gate490inter1));
  and2  gate2971(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate2972(.a(s_346), .O(gate490inter3));
  inv1  gate2973(.a(s_347), .O(gate490inter4));
  nand2 gate2974(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate2975(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate2976(.a(G1242), .O(gate490inter7));
  inv1  gate2977(.a(G1243), .O(gate490inter8));
  nand2 gate2978(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate2979(.a(s_347), .b(gate490inter3), .O(gate490inter10));
  nor2  gate2980(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate2981(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate2982(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate2563(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate2564(.a(gate492inter0), .b(s_288), .O(gate492inter1));
  and2  gate2565(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate2566(.a(s_288), .O(gate492inter3));
  inv1  gate2567(.a(s_289), .O(gate492inter4));
  nand2 gate2568(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate2569(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate2570(.a(G1246), .O(gate492inter7));
  inv1  gate2571(.a(G1247), .O(gate492inter8));
  nand2 gate2572(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate2573(.a(s_289), .b(gate492inter3), .O(gate492inter10));
  nor2  gate2574(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate2575(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate2576(.a(gate492inter12), .b(gate492inter1), .O(G1301));
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );

  xor2  gate1135(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate1136(.a(gate495inter0), .b(s_84), .O(gate495inter1));
  and2  gate1137(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate1138(.a(s_84), .O(gate495inter3));
  inv1  gate1139(.a(s_85), .O(gate495inter4));
  nand2 gate1140(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate1141(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate1142(.a(G1252), .O(gate495inter7));
  inv1  gate1143(.a(G1253), .O(gate495inter8));
  nand2 gate1144(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate1145(.a(s_85), .b(gate495inter3), .O(gate495inter10));
  nor2  gate1146(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate1147(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate1148(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate2059(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate2060(.a(gate501inter0), .b(s_216), .O(gate501inter1));
  and2  gate2061(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate2062(.a(s_216), .O(gate501inter3));
  inv1  gate2063(.a(s_217), .O(gate501inter4));
  nand2 gate2064(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate2065(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate2066(.a(G1264), .O(gate501inter7));
  inv1  gate2067(.a(G1265), .O(gate501inter8));
  nand2 gate2068(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate2069(.a(s_217), .b(gate501inter3), .O(gate501inter10));
  nor2  gate2070(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate2071(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate2072(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );

  xor2  gate659(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate660(.a(gate505inter0), .b(s_16), .O(gate505inter1));
  and2  gate661(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate662(.a(s_16), .O(gate505inter3));
  inv1  gate663(.a(s_17), .O(gate505inter4));
  nand2 gate664(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate665(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate666(.a(G1272), .O(gate505inter7));
  inv1  gate667(.a(G1273), .O(gate505inter8));
  nand2 gate668(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate669(.a(s_17), .b(gate505inter3), .O(gate505inter10));
  nor2  gate670(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate671(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate672(.a(gate505inter12), .b(gate505inter1), .O(G1314));
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate2143(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate2144(.a(gate508inter0), .b(s_228), .O(gate508inter1));
  and2  gate2145(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate2146(.a(s_228), .O(gate508inter3));
  inv1  gate2147(.a(s_229), .O(gate508inter4));
  nand2 gate2148(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate2149(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate2150(.a(G1278), .O(gate508inter7));
  inv1  gate2151(.a(G1279), .O(gate508inter8));
  nand2 gate2152(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate2153(.a(s_229), .b(gate508inter3), .O(gate508inter10));
  nor2  gate2154(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate2155(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate2156(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate1625(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate1626(.a(gate510inter0), .b(s_154), .O(gate510inter1));
  and2  gate1627(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate1628(.a(s_154), .O(gate510inter3));
  inv1  gate1629(.a(s_155), .O(gate510inter4));
  nand2 gate1630(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate1631(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate1632(.a(G1282), .O(gate510inter7));
  inv1  gate1633(.a(G1283), .O(gate510inter8));
  nand2 gate1634(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate1635(.a(s_155), .b(gate510inter3), .O(gate510inter10));
  nor2  gate1636(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate1637(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate1638(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate2633(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate2634(.a(gate514inter0), .b(s_298), .O(gate514inter1));
  and2  gate2635(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate2636(.a(s_298), .O(gate514inter3));
  inv1  gate2637(.a(s_299), .O(gate514inter4));
  nand2 gate2638(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate2639(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate2640(.a(G1290), .O(gate514inter7));
  inv1  gate2641(.a(G1291), .O(gate514inter8));
  nand2 gate2642(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate2643(.a(s_299), .b(gate514inter3), .O(gate514inter10));
  nor2  gate2644(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate2645(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate2646(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule