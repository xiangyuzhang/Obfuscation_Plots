module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate163inter0, gate163inter1, gate163inter2, gate163inter3, gate163inter4, gate163inter5, gate163inter6, gate163inter7, gate163inter8, gate163inter9, gate163inter10, gate163inter11, gate163inter12, gate392inter0, gate392inter1, gate392inter2, gate392inter3, gate392inter4, gate392inter5, gate392inter6, gate392inter7, gate392inter8, gate392inter9, gate392inter10, gate392inter11, gate392inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate161inter0, gate161inter1, gate161inter2, gate161inter3, gate161inter4, gate161inter5, gate161inter6, gate161inter7, gate161inter8, gate161inter9, gate161inter10, gate161inter11, gate161inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate253inter0, gate253inter1, gate253inter2, gate253inter3, gate253inter4, gate253inter5, gate253inter6, gate253inter7, gate253inter8, gate253inter9, gate253inter10, gate253inter11, gate253inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate474inter0, gate474inter1, gate474inter2, gate474inter3, gate474inter4, gate474inter5, gate474inter6, gate474inter7, gate474inter8, gate474inter9, gate474inter10, gate474inter11, gate474inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate214inter0, gate214inter1, gate214inter2, gate214inter3, gate214inter4, gate214inter5, gate214inter6, gate214inter7, gate214inter8, gate214inter9, gate214inter10, gate214inter11, gate214inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate468inter0, gate468inter1, gate468inter2, gate468inter3, gate468inter4, gate468inter5, gate468inter6, gate468inter7, gate468inter8, gate468inter9, gate468inter10, gate468inter11, gate468inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate1191(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate1192(.a(gate9inter0), .b(s_92), .O(gate9inter1));
  and2  gate1193(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate1194(.a(s_92), .O(gate9inter3));
  inv1  gate1195(.a(s_93), .O(gate9inter4));
  nand2 gate1196(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate1197(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate1198(.a(G1), .O(gate9inter7));
  inv1  gate1199(.a(G2), .O(gate9inter8));
  nand2 gate1200(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate1201(.a(s_93), .b(gate9inter3), .O(gate9inter10));
  nor2  gate1202(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate1203(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate1204(.a(gate9inter12), .b(gate9inter1), .O(G266));
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate701(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate702(.a(gate22inter0), .b(s_22), .O(gate22inter1));
  and2  gate703(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate704(.a(s_22), .O(gate22inter3));
  inv1  gate705(.a(s_23), .O(gate22inter4));
  nand2 gate706(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate707(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate708(.a(G27), .O(gate22inter7));
  inv1  gate709(.a(G28), .O(gate22inter8));
  nand2 gate710(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate711(.a(s_23), .b(gate22inter3), .O(gate22inter10));
  nor2  gate712(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate713(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate714(.a(gate22inter12), .b(gate22inter1), .O(G305));
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );

  xor2  gate771(.a(G5), .b(G1), .O(gate25inter0));
  nand2 gate772(.a(gate25inter0), .b(s_32), .O(gate25inter1));
  and2  gate773(.a(G5), .b(G1), .O(gate25inter2));
  inv1  gate774(.a(s_32), .O(gate25inter3));
  inv1  gate775(.a(s_33), .O(gate25inter4));
  nand2 gate776(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate777(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate778(.a(G1), .O(gate25inter7));
  inv1  gate779(.a(G5), .O(gate25inter8));
  nand2 gate780(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate781(.a(s_33), .b(gate25inter3), .O(gate25inter10));
  nor2  gate782(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate783(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate784(.a(gate25inter12), .b(gate25inter1), .O(G314));
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate729(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate730(.a(gate27inter0), .b(s_26), .O(gate27inter1));
  and2  gate731(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate732(.a(s_26), .O(gate27inter3));
  inv1  gate733(.a(s_27), .O(gate27inter4));
  nand2 gate734(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate735(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate736(.a(G2), .O(gate27inter7));
  inv1  gate737(.a(G6), .O(gate27inter8));
  nand2 gate738(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate739(.a(s_27), .b(gate27inter3), .O(gate27inter10));
  nor2  gate740(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate741(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate742(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );

  xor2  gate1065(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate1066(.a(gate38inter0), .b(s_74), .O(gate38inter1));
  and2  gate1067(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate1068(.a(s_74), .O(gate38inter3));
  inv1  gate1069(.a(s_75), .O(gate38inter4));
  nand2 gate1070(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate1071(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate1072(.a(G27), .O(gate38inter7));
  inv1  gate1073(.a(G31), .O(gate38inter8));
  nand2 gate1074(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate1075(.a(s_75), .b(gate38inter3), .O(gate38inter10));
  nor2  gate1076(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate1077(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate1078(.a(gate38inter12), .b(gate38inter1), .O(G353));
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );

  xor2  gate967(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate968(.a(gate52inter0), .b(s_60), .O(gate52inter1));
  and2  gate969(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate970(.a(s_60), .O(gate52inter3));
  inv1  gate971(.a(s_61), .O(gate52inter4));
  nand2 gate972(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate973(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate974(.a(G12), .O(gate52inter7));
  inv1  gate975(.a(G281), .O(gate52inter8));
  nand2 gate976(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate977(.a(s_61), .b(gate52inter3), .O(gate52inter10));
  nor2  gate978(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate979(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate980(.a(gate52inter12), .b(gate52inter1), .O(G373));
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate883(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate884(.a(gate59inter0), .b(s_48), .O(gate59inter1));
  and2  gate885(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate886(.a(s_48), .O(gate59inter3));
  inv1  gate887(.a(s_49), .O(gate59inter4));
  nand2 gate888(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate889(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate890(.a(G19), .O(gate59inter7));
  inv1  gate891(.a(G293), .O(gate59inter8));
  nand2 gate892(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate893(.a(s_49), .b(gate59inter3), .O(gate59inter10));
  nor2  gate894(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate895(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate896(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate995(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate996(.a(gate67inter0), .b(s_64), .O(gate67inter1));
  and2  gate997(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate998(.a(s_64), .O(gate67inter3));
  inv1  gate999(.a(s_65), .O(gate67inter4));
  nand2 gate1000(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate1001(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate1002(.a(G27), .O(gate67inter7));
  inv1  gate1003(.a(G305), .O(gate67inter8));
  nand2 gate1004(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate1005(.a(s_65), .b(gate67inter3), .O(gate67inter10));
  nor2  gate1006(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate1007(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate1008(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );

  xor2  gate1415(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate1416(.a(gate72inter0), .b(s_124), .O(gate72inter1));
  and2  gate1417(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate1418(.a(s_124), .O(gate72inter3));
  inv1  gate1419(.a(s_125), .O(gate72inter4));
  nand2 gate1420(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate1421(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate1422(.a(G32), .O(gate72inter7));
  inv1  gate1423(.a(G311), .O(gate72inter8));
  nand2 gate1424(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate1425(.a(s_125), .b(gate72inter3), .O(gate72inter10));
  nor2  gate1426(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate1427(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate1428(.a(gate72inter12), .b(gate72inter1), .O(G393));
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );

  xor2  gate1163(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate1164(.a(gate89inter0), .b(s_88), .O(gate89inter1));
  and2  gate1165(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate1166(.a(s_88), .O(gate89inter3));
  inv1  gate1167(.a(s_89), .O(gate89inter4));
  nand2 gate1168(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate1169(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate1170(.a(G17), .O(gate89inter7));
  inv1  gate1171(.a(G338), .O(gate89inter8));
  nand2 gate1172(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate1173(.a(s_89), .b(gate89inter3), .O(gate89inter10));
  nor2  gate1174(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate1175(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate1176(.a(gate89inter12), .b(gate89inter1), .O(G410));

  xor2  gate617(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate618(.a(gate90inter0), .b(s_10), .O(gate90inter1));
  and2  gate619(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate620(.a(s_10), .O(gate90inter3));
  inv1  gate621(.a(s_11), .O(gate90inter4));
  nand2 gate622(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate623(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate624(.a(G21), .O(gate90inter7));
  inv1  gate625(.a(G338), .O(gate90inter8));
  nand2 gate626(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate627(.a(s_11), .b(gate90inter3), .O(gate90inter10));
  nor2  gate628(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate629(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate630(.a(gate90inter12), .b(gate90inter1), .O(G411));
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate925(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate926(.a(gate98inter0), .b(s_54), .O(gate98inter1));
  and2  gate927(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate928(.a(s_54), .O(gate98inter3));
  inv1  gate929(.a(s_55), .O(gate98inter4));
  nand2 gate930(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate931(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate932(.a(G23), .O(gate98inter7));
  inv1  gate933(.a(G350), .O(gate98inter8));
  nand2 gate934(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate935(.a(s_55), .b(gate98inter3), .O(gate98inter10));
  nor2  gate936(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate937(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate938(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate715(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate716(.a(gate106inter0), .b(s_24), .O(gate106inter1));
  and2  gate717(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate718(.a(s_24), .O(gate106inter3));
  inv1  gate719(.a(s_25), .O(gate106inter4));
  nand2 gate720(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate721(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate722(.a(G364), .O(gate106inter7));
  inv1  gate723(.a(G365), .O(gate106inter8));
  nand2 gate724(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate725(.a(s_25), .b(gate106inter3), .O(gate106inter10));
  nor2  gate726(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate727(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate728(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );

  xor2  gate1093(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate1094(.a(gate117inter0), .b(s_78), .O(gate117inter1));
  and2  gate1095(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate1096(.a(s_78), .O(gate117inter3));
  inv1  gate1097(.a(s_79), .O(gate117inter4));
  nand2 gate1098(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate1099(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate1100(.a(G386), .O(gate117inter7));
  inv1  gate1101(.a(G387), .O(gate117inter8));
  nand2 gate1102(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate1103(.a(s_79), .b(gate117inter3), .O(gate117inter10));
  nor2  gate1104(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate1105(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate1106(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate1205(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate1206(.a(gate125inter0), .b(s_94), .O(gate125inter1));
  and2  gate1207(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate1208(.a(s_94), .O(gate125inter3));
  inv1  gate1209(.a(s_95), .O(gate125inter4));
  nand2 gate1210(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate1211(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate1212(.a(G402), .O(gate125inter7));
  inv1  gate1213(.a(G403), .O(gate125inter8));
  nand2 gate1214(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate1215(.a(s_95), .b(gate125inter3), .O(gate125inter10));
  nor2  gate1216(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate1217(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate1218(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate743(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate744(.a(gate142inter0), .b(s_28), .O(gate142inter1));
  and2  gate745(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate746(.a(s_28), .O(gate142inter3));
  inv1  gate747(.a(s_29), .O(gate142inter4));
  nand2 gate748(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate749(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate750(.a(G456), .O(gate142inter7));
  inv1  gate751(.a(G459), .O(gate142inter8));
  nand2 gate752(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate753(.a(s_29), .b(gate142inter3), .O(gate142inter10));
  nor2  gate754(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate755(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate756(.a(gate142inter12), .b(gate142inter1), .O(G537));

  xor2  gate1247(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate1248(.a(gate143inter0), .b(s_100), .O(gate143inter1));
  and2  gate1249(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate1250(.a(s_100), .O(gate143inter3));
  inv1  gate1251(.a(s_101), .O(gate143inter4));
  nand2 gate1252(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate1253(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate1254(.a(G462), .O(gate143inter7));
  inv1  gate1255(.a(G465), .O(gate143inter8));
  nand2 gate1256(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate1257(.a(s_101), .b(gate143inter3), .O(gate143inter10));
  nor2  gate1258(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate1259(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate1260(.a(gate143inter12), .b(gate143inter1), .O(G540));
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );

  xor2  gate1317(.a(G513), .b(G510), .O(gate151inter0));
  nand2 gate1318(.a(gate151inter0), .b(s_110), .O(gate151inter1));
  and2  gate1319(.a(G513), .b(G510), .O(gate151inter2));
  inv1  gate1320(.a(s_110), .O(gate151inter3));
  inv1  gate1321(.a(s_111), .O(gate151inter4));
  nand2 gate1322(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate1323(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate1324(.a(G510), .O(gate151inter7));
  inv1  gate1325(.a(G513), .O(gate151inter8));
  nand2 gate1326(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate1327(.a(s_111), .b(gate151inter3), .O(gate151inter10));
  nor2  gate1328(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate1329(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate1330(.a(gate151inter12), .b(gate151inter1), .O(G564));
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );

  xor2  gate1219(.a(G525), .b(G432), .O(gate155inter0));
  nand2 gate1220(.a(gate155inter0), .b(s_96), .O(gate155inter1));
  and2  gate1221(.a(G525), .b(G432), .O(gate155inter2));
  inv1  gate1222(.a(s_96), .O(gate155inter3));
  inv1  gate1223(.a(s_97), .O(gate155inter4));
  nand2 gate1224(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate1225(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate1226(.a(G432), .O(gate155inter7));
  inv1  gate1227(.a(G525), .O(gate155inter8));
  nand2 gate1228(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate1229(.a(s_97), .b(gate155inter3), .O(gate155inter10));
  nor2  gate1230(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate1231(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate1232(.a(gate155inter12), .b(gate155inter1), .O(G572));
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );

  xor2  gate757(.a(G534), .b(G450), .O(gate161inter0));
  nand2 gate758(.a(gate161inter0), .b(s_30), .O(gate161inter1));
  and2  gate759(.a(G534), .b(G450), .O(gate161inter2));
  inv1  gate760(.a(s_30), .O(gate161inter3));
  inv1  gate761(.a(s_31), .O(gate161inter4));
  nand2 gate762(.a(gate161inter4), .b(gate161inter3), .O(gate161inter5));
  nor2  gate763(.a(gate161inter5), .b(gate161inter2), .O(gate161inter6));
  inv1  gate764(.a(G450), .O(gate161inter7));
  inv1  gate765(.a(G534), .O(gate161inter8));
  nand2 gate766(.a(gate161inter8), .b(gate161inter7), .O(gate161inter9));
  nand2 gate767(.a(s_31), .b(gate161inter3), .O(gate161inter10));
  nor2  gate768(.a(gate161inter10), .b(gate161inter9), .O(gate161inter11));
  nor2  gate769(.a(gate161inter11), .b(gate161inter6), .O(gate161inter12));
  nand2 gate770(.a(gate161inter12), .b(gate161inter1), .O(G578));
nand2 gate162( .a(G453), .b(G534), .O(G579) );

  xor2  gate575(.a(G537), .b(G456), .O(gate163inter0));
  nand2 gate576(.a(gate163inter0), .b(s_4), .O(gate163inter1));
  and2  gate577(.a(G537), .b(G456), .O(gate163inter2));
  inv1  gate578(.a(s_4), .O(gate163inter3));
  inv1  gate579(.a(s_5), .O(gate163inter4));
  nand2 gate580(.a(gate163inter4), .b(gate163inter3), .O(gate163inter5));
  nor2  gate581(.a(gate163inter5), .b(gate163inter2), .O(gate163inter6));
  inv1  gate582(.a(G456), .O(gate163inter7));
  inv1  gate583(.a(G537), .O(gate163inter8));
  nand2 gate584(.a(gate163inter8), .b(gate163inter7), .O(gate163inter9));
  nand2 gate585(.a(s_5), .b(gate163inter3), .O(gate163inter10));
  nor2  gate586(.a(gate163inter10), .b(gate163inter9), .O(gate163inter11));
  nor2  gate587(.a(gate163inter11), .b(gate163inter6), .O(gate163inter12));
  nand2 gate588(.a(gate163inter12), .b(gate163inter1), .O(G580));
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate687(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate688(.a(gate172inter0), .b(s_20), .O(gate172inter1));
  and2  gate689(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate690(.a(s_20), .O(gate172inter3));
  inv1  gate691(.a(s_21), .O(gate172inter4));
  nand2 gate692(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate693(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate694(.a(G483), .O(gate172inter7));
  inv1  gate695(.a(G549), .O(gate172inter8));
  nand2 gate696(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate697(.a(s_21), .b(gate172inter3), .O(gate172inter10));
  nor2  gate698(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate699(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate700(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );

  xor2  gate1401(.a(G561), .b(G507), .O(gate180inter0));
  nand2 gate1402(.a(gate180inter0), .b(s_122), .O(gate180inter1));
  and2  gate1403(.a(G561), .b(G507), .O(gate180inter2));
  inv1  gate1404(.a(s_122), .O(gate180inter3));
  inv1  gate1405(.a(s_123), .O(gate180inter4));
  nand2 gate1406(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate1407(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate1408(.a(G507), .O(gate180inter7));
  inv1  gate1409(.a(G561), .O(gate180inter8));
  nand2 gate1410(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate1411(.a(s_123), .b(gate180inter3), .O(gate180inter10));
  nor2  gate1412(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate1413(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate1414(.a(gate180inter12), .b(gate180inter1), .O(G597));
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate561(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate562(.a(gate186inter0), .b(s_2), .O(gate186inter1));
  and2  gate563(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate564(.a(s_2), .O(gate186inter3));
  inv1  gate565(.a(s_3), .O(gate186inter4));
  nand2 gate566(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate567(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate568(.a(G572), .O(gate186inter7));
  inv1  gate569(.a(G573), .O(gate186inter8));
  nand2 gate570(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate571(.a(s_3), .b(gate186inter3), .O(gate186inter10));
  nor2  gate572(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate573(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate574(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate1289(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate1290(.a(gate198inter0), .b(s_106), .O(gate198inter1));
  and2  gate1291(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate1292(.a(s_106), .O(gate198inter3));
  inv1  gate1293(.a(s_107), .O(gate198inter4));
  nand2 gate1294(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate1295(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate1296(.a(G596), .O(gate198inter7));
  inv1  gate1297(.a(G597), .O(gate198inter8));
  nand2 gate1298(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate1299(.a(s_107), .b(gate198inter3), .O(gate198inter10));
  nor2  gate1300(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate1301(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate1302(.a(gate198inter12), .b(gate198inter1), .O(G657));

  xor2  gate869(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate870(.a(gate199inter0), .b(s_46), .O(gate199inter1));
  and2  gate871(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate872(.a(s_46), .O(gate199inter3));
  inv1  gate873(.a(s_47), .O(gate199inter4));
  nand2 gate874(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate875(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate876(.a(G598), .O(gate199inter7));
  inv1  gate877(.a(G599), .O(gate199inter8));
  nand2 gate878(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate879(.a(s_47), .b(gate199inter3), .O(gate199inter10));
  nor2  gate880(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate881(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate882(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate1345(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate1346(.a(gate201inter0), .b(s_114), .O(gate201inter1));
  and2  gate1347(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate1348(.a(s_114), .O(gate201inter3));
  inv1  gate1349(.a(s_115), .O(gate201inter4));
  nand2 gate1350(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate1351(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate1352(.a(G602), .O(gate201inter7));
  inv1  gate1353(.a(G607), .O(gate201inter8));
  nand2 gate1354(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate1355(.a(s_115), .b(gate201inter3), .O(gate201inter10));
  nor2  gate1356(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate1357(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate1358(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate1233(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate1234(.a(gate206inter0), .b(s_98), .O(gate206inter1));
  and2  gate1235(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate1236(.a(s_98), .O(gate206inter3));
  inv1  gate1237(.a(s_99), .O(gate206inter4));
  nand2 gate1238(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate1239(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate1240(.a(G632), .O(gate206inter7));
  inv1  gate1241(.a(G637), .O(gate206inter8));
  nand2 gate1242(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate1243(.a(s_99), .b(gate206inter3), .O(gate206inter10));
  nor2  gate1244(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate1245(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate1246(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );

  xor2  gate827(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate828(.a(gate213inter0), .b(s_40), .O(gate213inter1));
  and2  gate829(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate830(.a(s_40), .O(gate213inter3));
  inv1  gate831(.a(s_41), .O(gate213inter4));
  nand2 gate832(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate833(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate834(.a(G602), .O(gate213inter7));
  inv1  gate835(.a(G672), .O(gate213inter8));
  nand2 gate836(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate837(.a(s_41), .b(gate213inter3), .O(gate213inter10));
  nor2  gate838(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate839(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate840(.a(gate213inter12), .b(gate213inter1), .O(G694));

  xor2  gate1261(.a(G672), .b(G612), .O(gate214inter0));
  nand2 gate1262(.a(gate214inter0), .b(s_102), .O(gate214inter1));
  and2  gate1263(.a(G672), .b(G612), .O(gate214inter2));
  inv1  gate1264(.a(s_102), .O(gate214inter3));
  inv1  gate1265(.a(s_103), .O(gate214inter4));
  nand2 gate1266(.a(gate214inter4), .b(gate214inter3), .O(gate214inter5));
  nor2  gate1267(.a(gate214inter5), .b(gate214inter2), .O(gate214inter6));
  inv1  gate1268(.a(G612), .O(gate214inter7));
  inv1  gate1269(.a(G672), .O(gate214inter8));
  nand2 gate1270(.a(gate214inter8), .b(gate214inter7), .O(gate214inter9));
  nand2 gate1271(.a(s_103), .b(gate214inter3), .O(gate214inter10));
  nor2  gate1272(.a(gate214inter10), .b(gate214inter9), .O(gate214inter11));
  nor2  gate1273(.a(gate214inter11), .b(gate214inter6), .O(gate214inter12));
  nand2 gate1274(.a(gate214inter12), .b(gate214inter1), .O(G695));
nand2 gate215( .a(G607), .b(G675), .O(G696) );

  xor2  gate1177(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate1178(.a(gate216inter0), .b(s_90), .O(gate216inter1));
  and2  gate1179(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate1180(.a(s_90), .O(gate216inter3));
  inv1  gate1181(.a(s_91), .O(gate216inter4));
  nand2 gate1182(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate1183(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate1184(.a(G617), .O(gate216inter7));
  inv1  gate1185(.a(G675), .O(gate216inter8));
  nand2 gate1186(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate1187(.a(s_91), .b(gate216inter3), .O(gate216inter10));
  nor2  gate1188(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate1189(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate1190(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );

  xor2  gate1275(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate1276(.a(gate230inter0), .b(s_104), .O(gate230inter1));
  and2  gate1277(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate1278(.a(s_104), .O(gate230inter3));
  inv1  gate1279(.a(s_105), .O(gate230inter4));
  nand2 gate1280(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate1281(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate1282(.a(G700), .O(gate230inter7));
  inv1  gate1283(.a(G701), .O(gate230inter8));
  nand2 gate1284(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate1285(.a(s_105), .b(gate230inter3), .O(gate230inter10));
  nor2  gate1286(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate1287(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate1288(.a(gate230inter12), .b(gate230inter1), .O(G721));
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );

  xor2  gate1037(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate1038(.a(gate235inter0), .b(s_70), .O(gate235inter1));
  and2  gate1039(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate1040(.a(s_70), .O(gate235inter3));
  inv1  gate1041(.a(s_71), .O(gate235inter4));
  nand2 gate1042(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate1043(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate1044(.a(G248), .O(gate235inter7));
  inv1  gate1045(.a(G724), .O(gate235inter8));
  nand2 gate1046(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate1047(.a(s_71), .b(gate235inter3), .O(gate235inter10));
  nor2  gate1048(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate1049(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate1050(.a(gate235inter12), .b(gate235inter1), .O(G736));
nand2 gate236( .a(G251), .b(G727), .O(G739) );

  xor2  gate855(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate856(.a(gate237inter0), .b(s_44), .O(gate237inter1));
  and2  gate857(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate858(.a(s_44), .O(gate237inter3));
  inv1  gate859(.a(s_45), .O(gate237inter4));
  nand2 gate860(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate861(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate862(.a(G254), .O(gate237inter7));
  inv1  gate863(.a(G706), .O(gate237inter8));
  nand2 gate864(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate865(.a(s_45), .b(gate237inter3), .O(gate237inter10));
  nor2  gate866(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate867(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate868(.a(gate237inter12), .b(gate237inter1), .O(G742));

  xor2  gate841(.a(G709), .b(G257), .O(gate238inter0));
  nand2 gate842(.a(gate238inter0), .b(s_42), .O(gate238inter1));
  and2  gate843(.a(G709), .b(G257), .O(gate238inter2));
  inv1  gate844(.a(s_42), .O(gate238inter3));
  inv1  gate845(.a(s_43), .O(gate238inter4));
  nand2 gate846(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate847(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate848(.a(G257), .O(gate238inter7));
  inv1  gate849(.a(G709), .O(gate238inter8));
  nand2 gate850(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate851(.a(s_43), .b(gate238inter3), .O(gate238inter10));
  nor2  gate852(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate853(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate854(.a(gate238inter12), .b(gate238inter1), .O(G745));
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate953(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate954(.a(gate241inter0), .b(s_58), .O(gate241inter1));
  and2  gate955(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate956(.a(s_58), .O(gate241inter3));
  inv1  gate957(.a(s_59), .O(gate241inter4));
  nand2 gate958(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate959(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate960(.a(G242), .O(gate241inter7));
  inv1  gate961(.a(G730), .O(gate241inter8));
  nand2 gate962(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate963(.a(s_59), .b(gate241inter3), .O(gate241inter10));
  nor2  gate964(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate965(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate966(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );

  xor2  gate547(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate548(.a(gate246inter0), .b(s_0), .O(gate246inter1));
  and2  gate549(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate550(.a(s_0), .O(gate246inter3));
  inv1  gate551(.a(s_1), .O(gate246inter4));
  nand2 gate552(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate553(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate554(.a(G724), .O(gate246inter7));
  inv1  gate555(.a(G736), .O(gate246inter8));
  nand2 gate556(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate557(.a(s_1), .b(gate246inter3), .O(gate246inter10));
  nor2  gate558(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate559(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate560(.a(gate246inter12), .b(gate246inter1), .O(G759));
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );

  xor2  gate911(.a(G748), .b(G260), .O(gate253inter0));
  nand2 gate912(.a(gate253inter0), .b(s_52), .O(gate253inter1));
  and2  gate913(.a(G748), .b(G260), .O(gate253inter2));
  inv1  gate914(.a(s_52), .O(gate253inter3));
  inv1  gate915(.a(s_53), .O(gate253inter4));
  nand2 gate916(.a(gate253inter4), .b(gate253inter3), .O(gate253inter5));
  nor2  gate917(.a(gate253inter5), .b(gate253inter2), .O(gate253inter6));
  inv1  gate918(.a(G260), .O(gate253inter7));
  inv1  gate919(.a(G748), .O(gate253inter8));
  nand2 gate920(.a(gate253inter8), .b(gate253inter7), .O(gate253inter9));
  nand2 gate921(.a(s_53), .b(gate253inter3), .O(gate253inter10));
  nor2  gate922(.a(gate253inter10), .b(gate253inter9), .O(gate253inter11));
  nor2  gate923(.a(gate253inter11), .b(gate253inter6), .O(gate253inter12));
  nand2 gate924(.a(gate253inter12), .b(gate253inter1), .O(G766));
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate1457(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate1458(.a(gate257inter0), .b(s_130), .O(gate257inter1));
  and2  gate1459(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate1460(.a(s_130), .O(gate257inter3));
  inv1  gate1461(.a(s_131), .O(gate257inter4));
  nand2 gate1462(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate1463(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate1464(.a(G754), .O(gate257inter7));
  inv1  gate1465(.a(G755), .O(gate257inter8));
  nand2 gate1466(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate1467(.a(s_131), .b(gate257inter3), .O(gate257inter10));
  nor2  gate1468(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate1469(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate1470(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate1079(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate1080(.a(gate262inter0), .b(s_76), .O(gate262inter1));
  and2  gate1081(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate1082(.a(s_76), .O(gate262inter3));
  inv1  gate1083(.a(s_77), .O(gate262inter4));
  nand2 gate1084(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate1085(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate1086(.a(G764), .O(gate262inter7));
  inv1  gate1087(.a(G765), .O(gate262inter8));
  nand2 gate1088(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate1089(.a(s_77), .b(gate262inter3), .O(gate262inter10));
  nor2  gate1090(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate1091(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate1092(.a(gate262inter12), .b(gate262inter1), .O(G785));
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );

  xor2  gate1387(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate1388(.a(gate277inter0), .b(s_120), .O(gate277inter1));
  and2  gate1389(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate1390(.a(s_120), .O(gate277inter3));
  inv1  gate1391(.a(s_121), .O(gate277inter4));
  nand2 gate1392(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate1393(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate1394(.a(G648), .O(gate277inter7));
  inv1  gate1395(.a(G800), .O(gate277inter8));
  nand2 gate1396(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate1397(.a(s_121), .b(gate277inter3), .O(gate277inter10));
  nor2  gate1398(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate1399(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate1400(.a(gate277inter12), .b(gate277inter1), .O(G822));
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate1429(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate1430(.a(gate292inter0), .b(s_126), .O(gate292inter1));
  and2  gate1431(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate1432(.a(s_126), .O(gate292inter3));
  inv1  gate1433(.a(s_127), .O(gate292inter4));
  nand2 gate1434(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate1435(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate1436(.a(G824), .O(gate292inter7));
  inv1  gate1437(.a(G825), .O(gate292inter8));
  nand2 gate1438(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate1439(.a(s_127), .b(gate292inter3), .O(gate292inter10));
  nor2  gate1440(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate1441(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate1442(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );

  xor2  gate1051(.a(G833), .b(G832), .O(gate294inter0));
  nand2 gate1052(.a(gate294inter0), .b(s_72), .O(gate294inter1));
  and2  gate1053(.a(G833), .b(G832), .O(gate294inter2));
  inv1  gate1054(.a(s_72), .O(gate294inter3));
  inv1  gate1055(.a(s_73), .O(gate294inter4));
  nand2 gate1056(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate1057(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate1058(.a(G832), .O(gate294inter7));
  inv1  gate1059(.a(G833), .O(gate294inter8));
  nand2 gate1060(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate1061(.a(s_73), .b(gate294inter3), .O(gate294inter10));
  nor2  gate1062(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate1063(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate1064(.a(gate294inter12), .b(gate294inter1), .O(G899));
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate1149(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate1150(.a(gate296inter0), .b(s_86), .O(gate296inter1));
  and2  gate1151(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate1152(.a(s_86), .O(gate296inter3));
  inv1  gate1153(.a(s_87), .O(gate296inter4));
  nand2 gate1154(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate1155(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate1156(.a(G826), .O(gate296inter7));
  inv1  gate1157(.a(G827), .O(gate296inter8));
  nand2 gate1158(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate1159(.a(s_87), .b(gate296inter3), .O(gate296inter10));
  nor2  gate1160(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate1161(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate1162(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate1009(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate1010(.a(gate388inter0), .b(s_66), .O(gate388inter1));
  and2  gate1011(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate1012(.a(s_66), .O(gate388inter3));
  inv1  gate1013(.a(s_67), .O(gate388inter4));
  nand2 gate1014(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate1015(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate1016(.a(G2), .O(gate388inter7));
  inv1  gate1017(.a(G1039), .O(gate388inter8));
  nand2 gate1018(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate1019(.a(s_67), .b(gate388inter3), .O(gate388inter10));
  nor2  gate1020(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate1021(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate1022(.a(gate388inter12), .b(gate388inter1), .O(G1135));
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate813(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate814(.a(gate391inter0), .b(s_38), .O(gate391inter1));
  and2  gate815(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate816(.a(s_38), .O(gate391inter3));
  inv1  gate817(.a(s_39), .O(gate391inter4));
  nand2 gate818(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate819(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate820(.a(G5), .O(gate391inter7));
  inv1  gate821(.a(G1048), .O(gate391inter8));
  nand2 gate822(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate823(.a(s_39), .b(gate391inter3), .O(gate391inter10));
  nor2  gate824(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate825(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate826(.a(gate391inter12), .b(gate391inter1), .O(G1144));

  xor2  gate589(.a(G1051), .b(G6), .O(gate392inter0));
  nand2 gate590(.a(gate392inter0), .b(s_6), .O(gate392inter1));
  and2  gate591(.a(G1051), .b(G6), .O(gate392inter2));
  inv1  gate592(.a(s_6), .O(gate392inter3));
  inv1  gate593(.a(s_7), .O(gate392inter4));
  nand2 gate594(.a(gate392inter4), .b(gate392inter3), .O(gate392inter5));
  nor2  gate595(.a(gate392inter5), .b(gate392inter2), .O(gate392inter6));
  inv1  gate596(.a(G6), .O(gate392inter7));
  inv1  gate597(.a(G1051), .O(gate392inter8));
  nand2 gate598(.a(gate392inter8), .b(gate392inter7), .O(gate392inter9));
  nand2 gate599(.a(s_7), .b(gate392inter3), .O(gate392inter10));
  nor2  gate600(.a(gate392inter10), .b(gate392inter9), .O(gate392inter11));
  nor2  gate601(.a(gate392inter11), .b(gate392inter6), .O(gate392inter12));
  nand2 gate602(.a(gate392inter12), .b(gate392inter1), .O(G1147));
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate1359(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate1360(.a(gate394inter0), .b(s_116), .O(gate394inter1));
  and2  gate1361(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate1362(.a(s_116), .O(gate394inter3));
  inv1  gate1363(.a(s_117), .O(gate394inter4));
  nand2 gate1364(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate1365(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate1366(.a(G8), .O(gate394inter7));
  inv1  gate1367(.a(G1057), .O(gate394inter8));
  nand2 gate1368(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate1369(.a(s_117), .b(gate394inter3), .O(gate394inter10));
  nor2  gate1370(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate1371(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate1372(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate897(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate898(.a(gate397inter0), .b(s_50), .O(gate397inter1));
  and2  gate899(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate900(.a(s_50), .O(gate397inter3));
  inv1  gate901(.a(s_51), .O(gate397inter4));
  nand2 gate902(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate903(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate904(.a(G11), .O(gate397inter7));
  inv1  gate905(.a(G1066), .O(gate397inter8));
  nand2 gate906(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate907(.a(s_51), .b(gate397inter3), .O(gate397inter10));
  nor2  gate908(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate909(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate910(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );

  xor2  gate1303(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate1304(.a(gate412inter0), .b(s_108), .O(gate412inter1));
  and2  gate1305(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate1306(.a(s_108), .O(gate412inter3));
  inv1  gate1307(.a(s_109), .O(gate412inter4));
  nand2 gate1308(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate1309(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate1310(.a(G26), .O(gate412inter7));
  inv1  gate1311(.a(G1111), .O(gate412inter8));
  nand2 gate1312(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate1313(.a(s_109), .b(gate412inter3), .O(gate412inter10));
  nor2  gate1314(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate1315(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate1316(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );

  xor2  gate631(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate632(.a(gate418inter0), .b(s_12), .O(gate418inter1));
  and2  gate633(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate634(.a(s_12), .O(gate418inter3));
  inv1  gate635(.a(s_13), .O(gate418inter4));
  nand2 gate636(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate637(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate638(.a(G32), .O(gate418inter7));
  inv1  gate639(.a(G1129), .O(gate418inter8));
  nand2 gate640(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate641(.a(s_13), .b(gate418inter3), .O(gate418inter10));
  nor2  gate642(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate643(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate644(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate1331(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1332(.a(gate420inter0), .b(s_112), .O(gate420inter1));
  and2  gate1333(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1334(.a(s_112), .O(gate420inter3));
  inv1  gate1335(.a(s_113), .O(gate420inter4));
  nand2 gate1336(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1337(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1338(.a(G1036), .O(gate420inter7));
  inv1  gate1339(.a(G1132), .O(gate420inter8));
  nand2 gate1340(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1341(.a(s_113), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1342(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1343(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1344(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );

  xor2  gate1373(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate1374(.a(gate424inter0), .b(s_118), .O(gate424inter1));
  and2  gate1375(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate1376(.a(s_118), .O(gate424inter3));
  inv1  gate1377(.a(s_119), .O(gate424inter4));
  nand2 gate1378(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate1379(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate1380(.a(G1042), .O(gate424inter7));
  inv1  gate1381(.a(G1138), .O(gate424inter8));
  nand2 gate1382(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate1383(.a(s_119), .b(gate424inter3), .O(gate424inter10));
  nor2  gate1384(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate1385(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate1386(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate1107(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate1108(.a(gate433inter0), .b(s_80), .O(gate433inter1));
  and2  gate1109(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate1110(.a(s_80), .O(gate433inter3));
  inv1  gate1111(.a(s_81), .O(gate433inter4));
  nand2 gate1112(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate1113(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate1114(.a(G8), .O(gate433inter7));
  inv1  gate1115(.a(G1153), .O(gate433inter8));
  nand2 gate1116(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate1117(.a(s_81), .b(gate433inter3), .O(gate433inter10));
  nor2  gate1118(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate1119(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate1120(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );

  xor2  gate1121(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate1122(.a(gate446inter0), .b(s_82), .O(gate446inter1));
  and2  gate1123(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate1124(.a(s_82), .O(gate446inter3));
  inv1  gate1125(.a(s_83), .O(gate446inter4));
  nand2 gate1126(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate1127(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate1128(.a(G1075), .O(gate446inter7));
  inv1  gate1129(.a(G1171), .O(gate446inter8));
  nand2 gate1130(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate1131(.a(s_83), .b(gate446inter3), .O(gate446inter10));
  nor2  gate1132(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate1133(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate1134(.a(gate446inter12), .b(gate446inter1), .O(G1255));
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate1023(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate1024(.a(gate457inter0), .b(s_68), .O(gate457inter1));
  and2  gate1025(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate1026(.a(s_68), .O(gate457inter3));
  inv1  gate1027(.a(s_69), .O(gate457inter4));
  nand2 gate1028(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate1029(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate1030(.a(G20), .O(gate457inter7));
  inv1  gate1031(.a(G1189), .O(gate457inter8));
  nand2 gate1032(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate1033(.a(s_69), .b(gate457inter3), .O(gate457inter10));
  nor2  gate1034(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate1035(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate1036(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate785(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate786(.a(gate459inter0), .b(s_34), .O(gate459inter1));
  and2  gate787(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate788(.a(s_34), .O(gate459inter3));
  inv1  gate789(.a(s_35), .O(gate459inter4));
  nand2 gate790(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate791(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate792(.a(G21), .O(gate459inter7));
  inv1  gate793(.a(G1192), .O(gate459inter8));
  nand2 gate794(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate795(.a(s_35), .b(gate459inter3), .O(gate459inter10));
  nor2  gate796(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate797(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate798(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate1135(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate1136(.a(gate463inter0), .b(s_84), .O(gate463inter1));
  and2  gate1137(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate1138(.a(s_84), .O(gate463inter3));
  inv1  gate1139(.a(s_85), .O(gate463inter4));
  nand2 gate1140(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate1141(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate1142(.a(G23), .O(gate463inter7));
  inv1  gate1143(.a(G1198), .O(gate463inter8));
  nand2 gate1144(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate1145(.a(s_85), .b(gate463inter3), .O(gate463inter10));
  nor2  gate1146(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate1147(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate1148(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate673(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate674(.a(gate465inter0), .b(s_18), .O(gate465inter1));
  and2  gate675(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate676(.a(s_18), .O(gate465inter3));
  inv1  gate677(.a(s_19), .O(gate465inter4));
  nand2 gate678(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate679(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate680(.a(G24), .O(gate465inter7));
  inv1  gate681(.a(G1201), .O(gate465inter8));
  nand2 gate682(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate683(.a(s_19), .b(gate465inter3), .O(gate465inter10));
  nor2  gate684(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate685(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate686(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );

  xor2  gate1443(.a(G1204), .b(G1108), .O(gate468inter0));
  nand2 gate1444(.a(gate468inter0), .b(s_128), .O(gate468inter1));
  and2  gate1445(.a(G1204), .b(G1108), .O(gate468inter2));
  inv1  gate1446(.a(s_128), .O(gate468inter3));
  inv1  gate1447(.a(s_129), .O(gate468inter4));
  nand2 gate1448(.a(gate468inter4), .b(gate468inter3), .O(gate468inter5));
  nor2  gate1449(.a(gate468inter5), .b(gate468inter2), .O(gate468inter6));
  inv1  gate1450(.a(G1108), .O(gate468inter7));
  inv1  gate1451(.a(G1204), .O(gate468inter8));
  nand2 gate1452(.a(gate468inter8), .b(gate468inter7), .O(gate468inter9));
  nand2 gate1453(.a(s_129), .b(gate468inter3), .O(gate468inter10));
  nor2  gate1454(.a(gate468inter10), .b(gate468inter9), .O(gate468inter11));
  nor2  gate1455(.a(gate468inter11), .b(gate468inter6), .O(gate468inter12));
  nand2 gate1456(.a(gate468inter12), .b(gate468inter1), .O(G1277));
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );

  xor2  gate939(.a(G1213), .b(G1117), .O(gate474inter0));
  nand2 gate940(.a(gate474inter0), .b(s_56), .O(gate474inter1));
  and2  gate941(.a(G1213), .b(G1117), .O(gate474inter2));
  inv1  gate942(.a(s_56), .O(gate474inter3));
  inv1  gate943(.a(s_57), .O(gate474inter4));
  nand2 gate944(.a(gate474inter4), .b(gate474inter3), .O(gate474inter5));
  nor2  gate945(.a(gate474inter5), .b(gate474inter2), .O(gate474inter6));
  inv1  gate946(.a(G1117), .O(gate474inter7));
  inv1  gate947(.a(G1213), .O(gate474inter8));
  nand2 gate948(.a(gate474inter8), .b(gate474inter7), .O(gate474inter9));
  nand2 gate949(.a(s_57), .b(gate474inter3), .O(gate474inter10));
  nor2  gate950(.a(gate474inter10), .b(gate474inter9), .O(gate474inter11));
  nor2  gate951(.a(gate474inter11), .b(gate474inter6), .O(gate474inter12));
  nand2 gate952(.a(gate474inter12), .b(gate474inter1), .O(G1283));
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate645(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate646(.a(gate480inter0), .b(s_14), .O(gate480inter1));
  and2  gate647(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate648(.a(s_14), .O(gate480inter3));
  inv1  gate649(.a(s_15), .O(gate480inter4));
  nand2 gate650(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate651(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate652(.a(G1126), .O(gate480inter7));
  inv1  gate653(.a(G1222), .O(gate480inter8));
  nand2 gate654(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate655(.a(s_15), .b(gate480inter3), .O(gate480inter10));
  nor2  gate656(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate657(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate658(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );

  xor2  gate799(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate800(.a(gate484inter0), .b(s_36), .O(gate484inter1));
  and2  gate801(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate802(.a(s_36), .O(gate484inter3));
  inv1  gate803(.a(s_37), .O(gate484inter4));
  nand2 gate804(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate805(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate806(.a(G1230), .O(gate484inter7));
  inv1  gate807(.a(G1231), .O(gate484inter8));
  nand2 gate808(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate809(.a(s_37), .b(gate484inter3), .O(gate484inter10));
  nor2  gate810(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate811(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate812(.a(gate484inter12), .b(gate484inter1), .O(G1293));
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate981(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate982(.a(gate487inter0), .b(s_62), .O(gate487inter1));
  and2  gate983(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate984(.a(s_62), .O(gate487inter3));
  inv1  gate985(.a(s_63), .O(gate487inter4));
  nand2 gate986(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate987(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate988(.a(G1236), .O(gate487inter7));
  inv1  gate989(.a(G1237), .O(gate487inter8));
  nand2 gate990(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate991(.a(s_63), .b(gate487inter3), .O(gate487inter10));
  nor2  gate992(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate993(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate994(.a(gate487inter12), .b(gate487inter1), .O(G1296));
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );

  xor2  gate659(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate660(.a(gate498inter0), .b(s_16), .O(gate498inter1));
  and2  gate661(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate662(.a(s_16), .O(gate498inter3));
  inv1  gate663(.a(s_17), .O(gate498inter4));
  nand2 gate664(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate665(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate666(.a(G1258), .O(gate498inter7));
  inv1  gate667(.a(G1259), .O(gate498inter8));
  nand2 gate668(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate669(.a(s_17), .b(gate498inter3), .O(gate498inter10));
  nor2  gate670(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate671(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate672(.a(gate498inter12), .b(gate498inter1), .O(G1307));
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate603(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate604(.a(gate500inter0), .b(s_8), .O(gate500inter1));
  and2  gate605(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate606(.a(s_8), .O(gate500inter3));
  inv1  gate607(.a(s_9), .O(gate500inter4));
  nand2 gate608(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate609(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate610(.a(G1262), .O(gate500inter7));
  inv1  gate611(.a(G1263), .O(gate500inter8));
  nand2 gate612(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate613(.a(s_9), .b(gate500inter3), .O(gate500inter10));
  nor2  gate614(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate615(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate616(.a(gate500inter12), .b(gate500inter1), .O(G1309));
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule