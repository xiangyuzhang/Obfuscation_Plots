module c499 (N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
             N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
             N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
             N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
             N137,N724,N725,N726,N727,N728,N729,N730,N731,N732,
             N733,N734,N735,N736,N737,N738,N739,N740,N741,N742,
             N743,N744,N745,N746,N747,N748,N749,N750,N751,N752,
             N753,N754,N755);
input N1,N5,N9,N13,N17,N21,N25,N29,N33,N37,
      N41,N45,N49,N53,N57,N61,N65,N69,N73,N77,
      N81,N85,N89,N93,N97,N101,N105,N109,N113,N117,
      N121,N125,N129,N130,N131,N132,N133,N134,N135,N136,
      N137;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51;
output N724,N725,N726,N727,N728,N729,N730,N731,N732,N733,
       N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
       N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
       N754,N755;
wire N250,N251,N252,N253,N254,N255,N256,N257,N258,N259,
     N260,N261,N262,N263,N264,N265,N266,N267,N268,N269,
     N270,N271,N272,N273,N274,N275,N276,N277,N278,N279,
     N280,N281,N282,N283,N284,N285,N286,N287,N288,N289,
     N290,N293,N296,N299,N302,N305,N308,N311,N314,N315,
     N316,N317,N318,N319,N320,N321,N338,N339,N340,N341,
     N342,N343,N344,N345,N346,N347,N348,N349,N350,N351,
     N352,N353,N354,N367,N380,N393,N406,N419,N432,N445,
     N554,N555,N556,N557,N558,N559,N560,N561,N562,N563,
     N564,N565,N566,N567,N568,N569,N570,N571,N572,N573,
     N574,N575,N576,N577,N578,N579,N580,N581,N582,N583,
     N584,N585,N586,N587,N588,N589,N590,N591,N592,N593,
     N594,N595,N596,N597,N598,N599,N600,N601,N602,N607,
     N620,N625,N630,N635,N640,N645,N650,N655,N692,N693,
     N694,N695,N696,N697,N698,N699,N700,N701,N702,N703,
     N704,N705,N706,N707,N708,N709,N710,N711,N712,N713,
     N714,N715,N716,N717,N718,N719,N720,N721,N722,N723, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate8inter0, gate8inter1, gate8inter2, gate8inter3, gate8inter4, gate8inter5, gate8inter6, gate8inter7, gate8inter8, gate8inter9, gate8inter10, gate8inter11, gate8inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate35inter0, gate35inter1, gate35inter2, gate35inter3, gate35inter4, gate35inter5, gate35inter6, gate35inter7, gate35inter8, gate35inter9, gate35inter10, gate35inter11, gate35inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate14inter0, gate14inter1, gate14inter2, gate14inter3, gate14inter4, gate14inter5, gate14inter6, gate14inter7, gate14inter8, gate14inter9, gate14inter10, gate14inter11, gate14inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate190inter0, gate190inter1, gate190inter2, gate190inter3, gate190inter4, gate190inter5, gate190inter6, gate190inter7, gate190inter8, gate190inter9, gate190inter10, gate190inter11, gate190inter12, gate189inter0, gate189inter1, gate189inter2, gate189inter3, gate189inter4, gate189inter5, gate189inter6, gate189inter7, gate189inter8, gate189inter9, gate189inter10, gate189inter11, gate189inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate171inter0, gate171inter1, gate171inter2, gate171inter3, gate171inter4, gate171inter5, gate171inter6, gate171inter7, gate171inter8, gate171inter9, gate171inter10, gate171inter11, gate171inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate25inter0, gate25inter1, gate25inter2, gate25inter3, gate25inter4, gate25inter5, gate25inter6, gate25inter7, gate25inter8, gate25inter9, gate25inter10, gate25inter11, gate25inter12;


xor2 gate1( .a(N1), .b(N5), .O(N250) );
xor2 gate2( .a(N9), .b(N13), .O(N251) );
xor2 gate3( .a(N17), .b(N21), .O(N252) );
xor2 gate4( .a(N25), .b(N29), .O(N253) );
xor2 gate5( .a(N33), .b(N37), .O(N254) );
xor2 gate6( .a(N41), .b(N45), .O(N255) );
xor2 gate7( .a(N49), .b(N53), .O(N256) );

  xor2  gate287(.a(N61), .b(N57), .O(gate8inter0));
  nand2 gate288(.a(gate8inter0), .b(s_12), .O(gate8inter1));
  and2  gate289(.a(N61), .b(N57), .O(gate8inter2));
  inv1  gate290(.a(s_12), .O(gate8inter3));
  inv1  gate291(.a(s_13), .O(gate8inter4));
  nand2 gate292(.a(gate8inter4), .b(gate8inter3), .O(gate8inter5));
  nor2  gate293(.a(gate8inter5), .b(gate8inter2), .O(gate8inter6));
  inv1  gate294(.a(N57), .O(gate8inter7));
  inv1  gate295(.a(N61), .O(gate8inter8));
  nand2 gate296(.a(gate8inter8), .b(gate8inter7), .O(gate8inter9));
  nand2 gate297(.a(s_13), .b(gate8inter3), .O(gate8inter10));
  nor2  gate298(.a(gate8inter10), .b(gate8inter9), .O(gate8inter11));
  nor2  gate299(.a(gate8inter11), .b(gate8inter6), .O(gate8inter12));
  nand2 gate300(.a(gate8inter12), .b(gate8inter1), .O(N257));
xor2 gate9( .a(N65), .b(N69), .O(N258) );
xor2 gate10( .a(N73), .b(N77), .O(N259) );
xor2 gate11( .a(N81), .b(N85), .O(N260) );
xor2 gate12( .a(N89), .b(N93), .O(N261) );
xor2 gate13( .a(N97), .b(N101), .O(N262) );

  xor2  gate357(.a(N109), .b(N105), .O(gate14inter0));
  nand2 gate358(.a(gate14inter0), .b(s_22), .O(gate14inter1));
  and2  gate359(.a(N109), .b(N105), .O(gate14inter2));
  inv1  gate360(.a(s_22), .O(gate14inter3));
  inv1  gate361(.a(s_23), .O(gate14inter4));
  nand2 gate362(.a(gate14inter4), .b(gate14inter3), .O(gate14inter5));
  nor2  gate363(.a(gate14inter5), .b(gate14inter2), .O(gate14inter6));
  inv1  gate364(.a(N105), .O(gate14inter7));
  inv1  gate365(.a(N109), .O(gate14inter8));
  nand2 gate366(.a(gate14inter8), .b(gate14inter7), .O(gate14inter9));
  nand2 gate367(.a(s_23), .b(gate14inter3), .O(gate14inter10));
  nor2  gate368(.a(gate14inter10), .b(gate14inter9), .O(gate14inter11));
  nor2  gate369(.a(gate14inter11), .b(gate14inter6), .O(gate14inter12));
  nand2 gate370(.a(gate14inter12), .b(gate14inter1), .O(N263));
xor2 gate15( .a(N113), .b(N117), .O(N264) );
xor2 gate16( .a(N121), .b(N125), .O(N265) );
and2 gate17( .a(N129), .b(N137), .O(N266) );
and2 gate18( .a(N130), .b(N137), .O(N267) );
and2 gate19( .a(N131), .b(N137), .O(N268) );
and2 gate20( .a(N132), .b(N137), .O(N269) );
and2 gate21( .a(N133), .b(N137), .O(N270) );
and2 gate22( .a(N134), .b(N137), .O(N271) );
and2 gate23( .a(N135), .b(N137), .O(N272) );
and2 gate24( .a(N136), .b(N137), .O(N273) );

  xor2  gate553(.a(N17), .b(N1), .O(gate25inter0));
  nand2 gate554(.a(gate25inter0), .b(s_50), .O(gate25inter1));
  and2  gate555(.a(N17), .b(N1), .O(gate25inter2));
  inv1  gate556(.a(s_50), .O(gate25inter3));
  inv1  gate557(.a(s_51), .O(gate25inter4));
  nand2 gate558(.a(gate25inter4), .b(gate25inter3), .O(gate25inter5));
  nor2  gate559(.a(gate25inter5), .b(gate25inter2), .O(gate25inter6));
  inv1  gate560(.a(N1), .O(gate25inter7));
  inv1  gate561(.a(N17), .O(gate25inter8));
  nand2 gate562(.a(gate25inter8), .b(gate25inter7), .O(gate25inter9));
  nand2 gate563(.a(s_51), .b(gate25inter3), .O(gate25inter10));
  nor2  gate564(.a(gate25inter10), .b(gate25inter9), .O(gate25inter11));
  nor2  gate565(.a(gate25inter11), .b(gate25inter6), .O(gate25inter12));
  nand2 gate566(.a(gate25inter12), .b(gate25inter1), .O(N274));
xor2 gate26( .a(N33), .b(N49), .O(N275) );
xor2 gate27( .a(N5), .b(N21), .O(N276) );
xor2 gate28( .a(N37), .b(N53), .O(N277) );

  xor2  gate259(.a(N25), .b(N9), .O(gate29inter0));
  nand2 gate260(.a(gate29inter0), .b(s_8), .O(gate29inter1));
  and2  gate261(.a(N25), .b(N9), .O(gate29inter2));
  inv1  gate262(.a(s_8), .O(gate29inter3));
  inv1  gate263(.a(s_9), .O(gate29inter4));
  nand2 gate264(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate265(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate266(.a(N9), .O(gate29inter7));
  inv1  gate267(.a(N25), .O(gate29inter8));
  nand2 gate268(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate269(.a(s_9), .b(gate29inter3), .O(gate29inter10));
  nor2  gate270(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate271(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate272(.a(gate29inter12), .b(gate29inter1), .O(N278));
xor2 gate30( .a(N41), .b(N57), .O(N279) );
xor2 gate31( .a(N13), .b(N29), .O(N280) );
xor2 gate32( .a(N45), .b(N61), .O(N281) );
xor2 gate33( .a(N65), .b(N81), .O(N282) );
xor2 gate34( .a(N97), .b(N113), .O(N283) );

  xor2  gate329(.a(N85), .b(N69), .O(gate35inter0));
  nand2 gate330(.a(gate35inter0), .b(s_18), .O(gate35inter1));
  and2  gate331(.a(N85), .b(N69), .O(gate35inter2));
  inv1  gate332(.a(s_18), .O(gate35inter3));
  inv1  gate333(.a(s_19), .O(gate35inter4));
  nand2 gate334(.a(gate35inter4), .b(gate35inter3), .O(gate35inter5));
  nor2  gate335(.a(gate35inter5), .b(gate35inter2), .O(gate35inter6));
  inv1  gate336(.a(N69), .O(gate35inter7));
  inv1  gate337(.a(N85), .O(gate35inter8));
  nand2 gate338(.a(gate35inter8), .b(gate35inter7), .O(gate35inter9));
  nand2 gate339(.a(s_19), .b(gate35inter3), .O(gate35inter10));
  nor2  gate340(.a(gate35inter10), .b(gate35inter9), .O(gate35inter11));
  nor2  gate341(.a(gate35inter11), .b(gate35inter6), .O(gate35inter12));
  nand2 gate342(.a(gate35inter12), .b(gate35inter1), .O(N284));
xor2 gate36( .a(N101), .b(N117), .O(N285) );
xor2 gate37( .a(N73), .b(N89), .O(N286) );

  xor2  gate497(.a(N121), .b(N105), .O(gate38inter0));
  nand2 gate498(.a(gate38inter0), .b(s_42), .O(gate38inter1));
  and2  gate499(.a(N121), .b(N105), .O(gate38inter2));
  inv1  gate500(.a(s_42), .O(gate38inter3));
  inv1  gate501(.a(s_43), .O(gate38inter4));
  nand2 gate502(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate503(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate504(.a(N105), .O(gate38inter7));
  inv1  gate505(.a(N121), .O(gate38inter8));
  nand2 gate506(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate507(.a(s_43), .b(gate38inter3), .O(gate38inter10));
  nor2  gate508(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate509(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate510(.a(gate38inter12), .b(gate38inter1), .O(N287));

  xor2  gate483(.a(N93), .b(N77), .O(gate39inter0));
  nand2 gate484(.a(gate39inter0), .b(s_40), .O(gate39inter1));
  and2  gate485(.a(N93), .b(N77), .O(gate39inter2));
  inv1  gate486(.a(s_40), .O(gate39inter3));
  inv1  gate487(.a(s_41), .O(gate39inter4));
  nand2 gate488(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate489(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate490(.a(N77), .O(gate39inter7));
  inv1  gate491(.a(N93), .O(gate39inter8));
  nand2 gate492(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate493(.a(s_41), .b(gate39inter3), .O(gate39inter10));
  nor2  gate494(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate495(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate496(.a(gate39inter12), .b(gate39inter1), .O(N288));

  xor2  gate441(.a(N125), .b(N109), .O(gate40inter0));
  nand2 gate442(.a(gate40inter0), .b(s_34), .O(gate40inter1));
  and2  gate443(.a(N125), .b(N109), .O(gate40inter2));
  inv1  gate444(.a(s_34), .O(gate40inter3));
  inv1  gate445(.a(s_35), .O(gate40inter4));
  nand2 gate446(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate447(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate448(.a(N109), .O(gate40inter7));
  inv1  gate449(.a(N125), .O(gate40inter8));
  nand2 gate450(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate451(.a(s_35), .b(gate40inter3), .O(gate40inter10));
  nor2  gate452(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate453(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate454(.a(gate40inter12), .b(gate40inter1), .O(N289));
xor2 gate41( .a(N250), .b(N251), .O(N290) );
xor2 gate42( .a(N252), .b(N253), .O(N293) );
xor2 gate43( .a(N254), .b(N255), .O(N296) );
xor2 gate44( .a(N256), .b(N257), .O(N299) );
xor2 gate45( .a(N258), .b(N259), .O(N302) );

  xor2  gate343(.a(N261), .b(N260), .O(gate46inter0));
  nand2 gate344(.a(gate46inter0), .b(s_20), .O(gate46inter1));
  and2  gate345(.a(N261), .b(N260), .O(gate46inter2));
  inv1  gate346(.a(s_20), .O(gate46inter3));
  inv1  gate347(.a(s_21), .O(gate46inter4));
  nand2 gate348(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate349(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate350(.a(N260), .O(gate46inter7));
  inv1  gate351(.a(N261), .O(gate46inter8));
  nand2 gate352(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate353(.a(s_21), .b(gate46inter3), .O(gate46inter10));
  nor2  gate354(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate355(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate356(.a(gate46inter12), .b(gate46inter1), .O(N305));
xor2 gate47( .a(N262), .b(N263), .O(N308) );
xor2 gate48( .a(N264), .b(N265), .O(N311) );
xor2 gate49( .a(N274), .b(N275), .O(N314) );
xor2 gate50( .a(N276), .b(N277), .O(N315) );
xor2 gate51( .a(N278), .b(N279), .O(N316) );
xor2 gate52( .a(N280), .b(N281), .O(N317) );
xor2 gate53( .a(N282), .b(N283), .O(N318) );
xor2 gate54( .a(N284), .b(N285), .O(N319) );
xor2 gate55( .a(N286), .b(N287), .O(N320) );
xor2 gate56( .a(N288), .b(N289), .O(N321) );
xor2 gate57( .a(N290), .b(N293), .O(N338) );
xor2 gate58( .a(N296), .b(N299), .O(N339) );

  xor2  gate301(.a(N296), .b(N290), .O(gate59inter0));
  nand2 gate302(.a(gate59inter0), .b(s_14), .O(gate59inter1));
  and2  gate303(.a(N296), .b(N290), .O(gate59inter2));
  inv1  gate304(.a(s_14), .O(gate59inter3));
  inv1  gate305(.a(s_15), .O(gate59inter4));
  nand2 gate306(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate307(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate308(.a(N290), .O(gate59inter7));
  inv1  gate309(.a(N296), .O(gate59inter8));
  nand2 gate310(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate311(.a(s_15), .b(gate59inter3), .O(gate59inter10));
  nor2  gate312(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate313(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate314(.a(gate59inter12), .b(gate59inter1), .O(N340));

  xor2  gate245(.a(N299), .b(N293), .O(gate60inter0));
  nand2 gate246(.a(gate60inter0), .b(s_6), .O(gate60inter1));
  and2  gate247(.a(N299), .b(N293), .O(gate60inter2));
  inv1  gate248(.a(s_6), .O(gate60inter3));
  inv1  gate249(.a(s_7), .O(gate60inter4));
  nand2 gate250(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate251(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate252(.a(N293), .O(gate60inter7));
  inv1  gate253(.a(N299), .O(gate60inter8));
  nand2 gate254(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate255(.a(s_7), .b(gate60inter3), .O(gate60inter10));
  nor2  gate256(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate257(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate258(.a(gate60inter12), .b(gate60inter1), .O(N341));
xor2 gate61( .a(N302), .b(N305), .O(N342) );
xor2 gate62( .a(N308), .b(N311), .O(N343) );

  xor2  gate231(.a(N308), .b(N302), .O(gate63inter0));
  nand2 gate232(.a(gate63inter0), .b(s_4), .O(gate63inter1));
  and2  gate233(.a(N308), .b(N302), .O(gate63inter2));
  inv1  gate234(.a(s_4), .O(gate63inter3));
  inv1  gate235(.a(s_5), .O(gate63inter4));
  nand2 gate236(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate237(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate238(.a(N302), .O(gate63inter7));
  inv1  gate239(.a(N308), .O(gate63inter8));
  nand2 gate240(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate241(.a(s_5), .b(gate63inter3), .O(gate63inter10));
  nor2  gate242(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate243(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate244(.a(gate63inter12), .b(gate63inter1), .O(N344));
xor2 gate64( .a(N305), .b(N311), .O(N345) );
xor2 gate65( .a(N266), .b(N342), .O(N346) );
xor2 gate66( .a(N267), .b(N343), .O(N347) );
xor2 gate67( .a(N268), .b(N344), .O(N348) );
xor2 gate68( .a(N269), .b(N345), .O(N349) );
xor2 gate69( .a(N270), .b(N338), .O(N350) );
xor2 gate70( .a(N271), .b(N339), .O(N351) );

  xor2  gate413(.a(N340), .b(N272), .O(gate71inter0));
  nand2 gate414(.a(gate71inter0), .b(s_30), .O(gate71inter1));
  and2  gate415(.a(N340), .b(N272), .O(gate71inter2));
  inv1  gate416(.a(s_30), .O(gate71inter3));
  inv1  gate417(.a(s_31), .O(gate71inter4));
  nand2 gate418(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate419(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate420(.a(N272), .O(gate71inter7));
  inv1  gate421(.a(N340), .O(gate71inter8));
  nand2 gate422(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate423(.a(s_31), .b(gate71inter3), .O(gate71inter10));
  nor2  gate424(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate425(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate426(.a(gate71inter12), .b(gate71inter1), .O(N352));
xor2 gate72( .a(N273), .b(N341), .O(N353) );

  xor2  gate371(.a(N346), .b(N314), .O(gate73inter0));
  nand2 gate372(.a(gate73inter0), .b(s_24), .O(gate73inter1));
  and2  gate373(.a(N346), .b(N314), .O(gate73inter2));
  inv1  gate374(.a(s_24), .O(gate73inter3));
  inv1  gate375(.a(s_25), .O(gate73inter4));
  nand2 gate376(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate377(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate378(.a(N314), .O(gate73inter7));
  inv1  gate379(.a(N346), .O(gate73inter8));
  nand2 gate380(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate381(.a(s_25), .b(gate73inter3), .O(gate73inter10));
  nor2  gate382(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate383(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate384(.a(gate73inter12), .b(gate73inter1), .O(N354));
xor2 gate74( .a(N315), .b(N347), .O(N367) );
xor2 gate75( .a(N316), .b(N348), .O(N380) );

  xor2  gate203(.a(N349), .b(N317), .O(gate76inter0));
  nand2 gate204(.a(gate76inter0), .b(s_0), .O(gate76inter1));
  and2  gate205(.a(N349), .b(N317), .O(gate76inter2));
  inv1  gate206(.a(s_0), .O(gate76inter3));
  inv1  gate207(.a(s_1), .O(gate76inter4));
  nand2 gate208(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate209(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate210(.a(N317), .O(gate76inter7));
  inv1  gate211(.a(N349), .O(gate76inter8));
  nand2 gate212(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate213(.a(s_1), .b(gate76inter3), .O(gate76inter10));
  nor2  gate214(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate215(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate216(.a(gate76inter12), .b(gate76inter1), .O(N393));
xor2 gate77( .a(N318), .b(N350), .O(N406) );
xor2 gate78( .a(N319), .b(N351), .O(N419) );

  xor2  gate455(.a(N352), .b(N320), .O(gate79inter0));
  nand2 gate456(.a(gate79inter0), .b(s_36), .O(gate79inter1));
  and2  gate457(.a(N352), .b(N320), .O(gate79inter2));
  inv1  gate458(.a(s_36), .O(gate79inter3));
  inv1  gate459(.a(s_37), .O(gate79inter4));
  nand2 gate460(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate461(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate462(.a(N320), .O(gate79inter7));
  inv1  gate463(.a(N352), .O(gate79inter8));
  nand2 gate464(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate465(.a(s_37), .b(gate79inter3), .O(gate79inter10));
  nor2  gate466(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate467(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate468(.a(gate79inter12), .b(gate79inter1), .O(N432));

  xor2  gate315(.a(N353), .b(N321), .O(gate80inter0));
  nand2 gate316(.a(gate80inter0), .b(s_16), .O(gate80inter1));
  and2  gate317(.a(N353), .b(N321), .O(gate80inter2));
  inv1  gate318(.a(s_16), .O(gate80inter3));
  inv1  gate319(.a(s_17), .O(gate80inter4));
  nand2 gate320(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate321(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate322(.a(N321), .O(gate80inter7));
  inv1  gate323(.a(N353), .O(gate80inter8));
  nand2 gate324(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate325(.a(s_17), .b(gate80inter3), .O(gate80inter10));
  nor2  gate326(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate327(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate328(.a(gate80inter12), .b(gate80inter1), .O(N445));
inv1 gate81( .a(N354), .O(N554) );
inv1 gate82( .a(N367), .O(N555) );
inv1 gate83( .a(N380), .O(N556) );
inv1 gate84( .a(N354), .O(N557) );
inv1 gate85( .a(N367), .O(N558) );
inv1 gate86( .a(N393), .O(N559) );
inv1 gate87( .a(N354), .O(N560) );
inv1 gate88( .a(N380), .O(N561) );
inv1 gate89( .a(N393), .O(N562) );
inv1 gate90( .a(N367), .O(N563) );
inv1 gate91( .a(N380), .O(N564) );
inv1 gate92( .a(N393), .O(N565) );
inv1 gate93( .a(N419), .O(N566) );
inv1 gate94( .a(N445), .O(N567) );
inv1 gate95( .a(N419), .O(N568) );
inv1 gate96( .a(N432), .O(N569) );
inv1 gate97( .a(N406), .O(N570) );
inv1 gate98( .a(N445), .O(N571) );
inv1 gate99( .a(N406), .O(N572) );
inv1 gate100( .a(N432), .O(N573) );
inv1 gate101( .a(N406), .O(N574) );
inv1 gate102( .a(N419), .O(N575) );
inv1 gate103( .a(N432), .O(N576) );
inv1 gate104( .a(N406), .O(N577) );
inv1 gate105( .a(N419), .O(N578) );
inv1 gate106( .a(N445), .O(N579) );
inv1 gate107( .a(N406), .O(N580) );
inv1 gate108( .a(N432), .O(N581) );
inv1 gate109( .a(N445), .O(N582) );
inv1 gate110( .a(N419), .O(N583) );
inv1 gate111( .a(N432), .O(N584) );
inv1 gate112( .a(N445), .O(N585) );
inv1 gate113( .a(N367), .O(N586) );
inv1 gate114( .a(N393), .O(N587) );
inv1 gate115( .a(N367), .O(N588) );
inv1 gate116( .a(N380), .O(N589) );
inv1 gate117( .a(N354), .O(N590) );
inv1 gate118( .a(N393), .O(N591) );
inv1 gate119( .a(N354), .O(N592) );
inv1 gate120( .a(N380), .O(N593) );
and4 gate121( .a(N554), .b(N555), .c(N556), .d(N393), .O(N594) );
and4 gate122( .a(N557), .b(N558), .c(N380), .d(N559), .O(N595) );
and4 gate123( .a(N560), .b(N367), .c(N561), .d(N562), .O(N596) );
and4 gate124( .a(N354), .b(N563), .c(N564), .d(N565), .O(N597) );
and4 gate125( .a(N574), .b(N575), .c(N576), .d(N445), .O(N598) );
and4 gate126( .a(N577), .b(N578), .c(N432), .d(N579), .O(N599) );
and4 gate127( .a(N580), .b(N419), .c(N581), .d(N582), .O(N600) );
and4 gate128( .a(N406), .b(N583), .c(N584), .d(N585), .O(N601) );
or4 gate129( .a(N594), .b(N595), .c(N596), .d(N597), .O(N602) );
or4 gate130( .a(N598), .b(N599), .c(N600), .d(N601), .O(N607) );
and5 gate131( .a(N406), .b(N566), .c(N432), .d(N567), .e(N602), .O(N620) );
and5 gate132( .a(N406), .b(N568), .c(N569), .d(N445), .e(N602), .O(N625) );
and5 gate133( .a(N570), .b(N419), .c(N432), .d(N571), .e(N602), .O(N630) );
and5 gate134( .a(N572), .b(N419), .c(N573), .d(N445), .e(N602), .O(N635) );
and5 gate135( .a(N354), .b(N586), .c(N380), .d(N587), .e(N607), .O(N640) );
and5 gate136( .a(N354), .b(N588), .c(N589), .d(N393), .e(N607), .O(N645) );
and5 gate137( .a(N590), .b(N367), .c(N380), .d(N591), .e(N607), .O(N650) );
and5 gate138( .a(N592), .b(N367), .c(N593), .d(N393), .e(N607), .O(N655) );
and2 gate139( .a(N354), .b(N620), .O(N692) );
and2 gate140( .a(N367), .b(N620), .O(N693) );
and2 gate141( .a(N380), .b(N620), .O(N694) );
and2 gate142( .a(N393), .b(N620), .O(N695) );
and2 gate143( .a(N354), .b(N625), .O(N696) );
and2 gate144( .a(N367), .b(N625), .O(N697) );
and2 gate145( .a(N380), .b(N625), .O(N698) );
and2 gate146( .a(N393), .b(N625), .O(N699) );
and2 gate147( .a(N354), .b(N630), .O(N700) );
and2 gate148( .a(N367), .b(N630), .O(N701) );
and2 gate149( .a(N380), .b(N630), .O(N702) );
and2 gate150( .a(N393), .b(N630), .O(N703) );
and2 gate151( .a(N354), .b(N635), .O(N704) );
and2 gate152( .a(N367), .b(N635), .O(N705) );
and2 gate153( .a(N380), .b(N635), .O(N706) );
and2 gate154( .a(N393), .b(N635), .O(N707) );
and2 gate155( .a(N406), .b(N640), .O(N708) );
and2 gate156( .a(N419), .b(N640), .O(N709) );
and2 gate157( .a(N432), .b(N640), .O(N710) );
and2 gate158( .a(N445), .b(N640), .O(N711) );
and2 gate159( .a(N406), .b(N645), .O(N712) );
and2 gate160( .a(N419), .b(N645), .O(N713) );
and2 gate161( .a(N432), .b(N645), .O(N714) );
and2 gate162( .a(N445), .b(N645), .O(N715) );
and2 gate163( .a(N406), .b(N650), .O(N716) );
and2 gate164( .a(N419), .b(N650), .O(N717) );
and2 gate165( .a(N432), .b(N650), .O(N718) );
and2 gate166( .a(N445), .b(N650), .O(N719) );
and2 gate167( .a(N406), .b(N655), .O(N720) );
and2 gate168( .a(N419), .b(N655), .O(N721) );
and2 gate169( .a(N432), .b(N655), .O(N722) );
and2 gate170( .a(N445), .b(N655), .O(N723) );

  xor2  gate511(.a(N692), .b(N1), .O(gate171inter0));
  nand2 gate512(.a(gate171inter0), .b(s_44), .O(gate171inter1));
  and2  gate513(.a(N692), .b(N1), .O(gate171inter2));
  inv1  gate514(.a(s_44), .O(gate171inter3));
  inv1  gate515(.a(s_45), .O(gate171inter4));
  nand2 gate516(.a(gate171inter4), .b(gate171inter3), .O(gate171inter5));
  nor2  gate517(.a(gate171inter5), .b(gate171inter2), .O(gate171inter6));
  inv1  gate518(.a(N1), .O(gate171inter7));
  inv1  gate519(.a(N692), .O(gate171inter8));
  nand2 gate520(.a(gate171inter8), .b(gate171inter7), .O(gate171inter9));
  nand2 gate521(.a(s_45), .b(gate171inter3), .O(gate171inter10));
  nor2  gate522(.a(gate171inter10), .b(gate171inter9), .O(gate171inter11));
  nor2  gate523(.a(gate171inter11), .b(gate171inter6), .O(gate171inter12));
  nand2 gate524(.a(gate171inter12), .b(gate171inter1), .O(N724));
xor2 gate172( .a(N5), .b(N693), .O(N725) );
xor2 gate173( .a(N9), .b(N694), .O(N726) );
xor2 gate174( .a(N13), .b(N695), .O(N727) );
xor2 gate175( .a(N17), .b(N696), .O(N728) );
xor2 gate176( .a(N21), .b(N697), .O(N729) );

  xor2  gate469(.a(N698), .b(N25), .O(gate177inter0));
  nand2 gate470(.a(gate177inter0), .b(s_38), .O(gate177inter1));
  and2  gate471(.a(N698), .b(N25), .O(gate177inter2));
  inv1  gate472(.a(s_38), .O(gate177inter3));
  inv1  gate473(.a(s_39), .O(gate177inter4));
  nand2 gate474(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate475(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate476(.a(N25), .O(gate177inter7));
  inv1  gate477(.a(N698), .O(gate177inter8));
  nand2 gate478(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate479(.a(s_39), .b(gate177inter3), .O(gate177inter10));
  nor2  gate480(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate481(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate482(.a(gate177inter12), .b(gate177inter1), .O(N730));

  xor2  gate273(.a(N699), .b(N29), .O(gate178inter0));
  nand2 gate274(.a(gate178inter0), .b(s_10), .O(gate178inter1));
  and2  gate275(.a(N699), .b(N29), .O(gate178inter2));
  inv1  gate276(.a(s_10), .O(gate178inter3));
  inv1  gate277(.a(s_11), .O(gate178inter4));
  nand2 gate278(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate279(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate280(.a(N29), .O(gate178inter7));
  inv1  gate281(.a(N699), .O(gate178inter8));
  nand2 gate282(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate283(.a(s_11), .b(gate178inter3), .O(gate178inter10));
  nor2  gate284(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate285(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate286(.a(gate178inter12), .b(gate178inter1), .O(N731));
xor2 gate179( .a(N33), .b(N700), .O(N732) );
xor2 gate180( .a(N37), .b(N701), .O(N733) );
xor2 gate181( .a(N41), .b(N702), .O(N734) );

  xor2  gate539(.a(N703), .b(N45), .O(gate182inter0));
  nand2 gate540(.a(gate182inter0), .b(s_48), .O(gate182inter1));
  and2  gate541(.a(N703), .b(N45), .O(gate182inter2));
  inv1  gate542(.a(s_48), .O(gate182inter3));
  inv1  gate543(.a(s_49), .O(gate182inter4));
  nand2 gate544(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate545(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate546(.a(N45), .O(gate182inter7));
  inv1  gate547(.a(N703), .O(gate182inter8));
  nand2 gate548(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate549(.a(s_49), .b(gate182inter3), .O(gate182inter10));
  nor2  gate550(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate551(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate552(.a(gate182inter12), .b(gate182inter1), .O(N735));
xor2 gate183( .a(N49), .b(N704), .O(N736) );

  xor2  gate427(.a(N705), .b(N53), .O(gate184inter0));
  nand2 gate428(.a(gate184inter0), .b(s_32), .O(gate184inter1));
  and2  gate429(.a(N705), .b(N53), .O(gate184inter2));
  inv1  gate430(.a(s_32), .O(gate184inter3));
  inv1  gate431(.a(s_33), .O(gate184inter4));
  nand2 gate432(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate433(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate434(.a(N53), .O(gate184inter7));
  inv1  gate435(.a(N705), .O(gate184inter8));
  nand2 gate436(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate437(.a(s_33), .b(gate184inter3), .O(gate184inter10));
  nor2  gate438(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate439(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate440(.a(gate184inter12), .b(gate184inter1), .O(N737));
xor2 gate185( .a(N57), .b(N706), .O(N738) );
xor2 gate186( .a(N61), .b(N707), .O(N739) );
xor2 gate187( .a(N65), .b(N708), .O(N740) );
xor2 gate188( .a(N69), .b(N709), .O(N741) );

  xor2  gate399(.a(N710), .b(N73), .O(gate189inter0));
  nand2 gate400(.a(gate189inter0), .b(s_28), .O(gate189inter1));
  and2  gate401(.a(N710), .b(N73), .O(gate189inter2));
  inv1  gate402(.a(s_28), .O(gate189inter3));
  inv1  gate403(.a(s_29), .O(gate189inter4));
  nand2 gate404(.a(gate189inter4), .b(gate189inter3), .O(gate189inter5));
  nor2  gate405(.a(gate189inter5), .b(gate189inter2), .O(gate189inter6));
  inv1  gate406(.a(N73), .O(gate189inter7));
  inv1  gate407(.a(N710), .O(gate189inter8));
  nand2 gate408(.a(gate189inter8), .b(gate189inter7), .O(gate189inter9));
  nand2 gate409(.a(s_29), .b(gate189inter3), .O(gate189inter10));
  nor2  gate410(.a(gate189inter10), .b(gate189inter9), .O(gate189inter11));
  nor2  gate411(.a(gate189inter11), .b(gate189inter6), .O(gate189inter12));
  nand2 gate412(.a(gate189inter12), .b(gate189inter1), .O(N742));

  xor2  gate385(.a(N711), .b(N77), .O(gate190inter0));
  nand2 gate386(.a(gate190inter0), .b(s_26), .O(gate190inter1));
  and2  gate387(.a(N711), .b(N77), .O(gate190inter2));
  inv1  gate388(.a(s_26), .O(gate190inter3));
  inv1  gate389(.a(s_27), .O(gate190inter4));
  nand2 gate390(.a(gate190inter4), .b(gate190inter3), .O(gate190inter5));
  nor2  gate391(.a(gate190inter5), .b(gate190inter2), .O(gate190inter6));
  inv1  gate392(.a(N77), .O(gate190inter7));
  inv1  gate393(.a(N711), .O(gate190inter8));
  nand2 gate394(.a(gate190inter8), .b(gate190inter7), .O(gate190inter9));
  nand2 gate395(.a(s_27), .b(gate190inter3), .O(gate190inter10));
  nor2  gate396(.a(gate190inter10), .b(gate190inter9), .O(gate190inter11));
  nor2  gate397(.a(gate190inter11), .b(gate190inter6), .O(gate190inter12));
  nand2 gate398(.a(gate190inter12), .b(gate190inter1), .O(N743));
xor2 gate191( .a(N81), .b(N712), .O(N744) );
xor2 gate192( .a(N85), .b(N713), .O(N745) );
xor2 gate193( .a(N89), .b(N714), .O(N746) );
xor2 gate194( .a(N93), .b(N715), .O(N747) );
xor2 gate195( .a(N97), .b(N716), .O(N748) );
xor2 gate196( .a(N101), .b(N717), .O(N749) );
xor2 gate197( .a(N105), .b(N718), .O(N750) );

  xor2  gate525(.a(N719), .b(N109), .O(gate198inter0));
  nand2 gate526(.a(gate198inter0), .b(s_46), .O(gate198inter1));
  and2  gate527(.a(N719), .b(N109), .O(gate198inter2));
  inv1  gate528(.a(s_46), .O(gate198inter3));
  inv1  gate529(.a(s_47), .O(gate198inter4));
  nand2 gate530(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate531(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate532(.a(N109), .O(gate198inter7));
  inv1  gate533(.a(N719), .O(gate198inter8));
  nand2 gate534(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate535(.a(s_47), .b(gate198inter3), .O(gate198inter10));
  nor2  gate536(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate537(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate538(.a(gate198inter12), .b(gate198inter1), .O(N751));
xor2 gate199( .a(N113), .b(N720), .O(N752) );
xor2 gate200( .a(N117), .b(N721), .O(N753) );

  xor2  gate217(.a(N722), .b(N121), .O(gate201inter0));
  nand2 gate218(.a(gate201inter0), .b(s_2), .O(gate201inter1));
  and2  gate219(.a(N722), .b(N121), .O(gate201inter2));
  inv1  gate220(.a(s_2), .O(gate201inter3));
  inv1  gate221(.a(s_3), .O(gate201inter4));
  nand2 gate222(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate223(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate224(.a(N121), .O(gate201inter7));
  inv1  gate225(.a(N722), .O(gate201inter8));
  nand2 gate226(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate227(.a(s_3), .b(gate201inter3), .O(gate201inter10));
  nor2  gate228(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate229(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate230(.a(gate201inter12), .b(gate201inter1), .O(N754));
xor2 gate202( .a(N125), .b(N723), .O(N755) );

endmodule