module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate213inter0, gate213inter1, gate213inter2, gate213inter3, gate213inter4, gate213inter5, gate213inter6, gate213inter7, gate213inter8, gate213inter9, gate213inter10, gate213inter11, gate213inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate11inter0, gate11inter1, gate11inter2, gate11inter3, gate11inter4, gate11inter5, gate11inter6, gate11inter7, gate11inter8, gate11inter9, gate11inter10, gate11inter11, gate11inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate505inter0, gate505inter1, gate505inter2, gate505inter3, gate505inter4, gate505inter5, gate505inter6, gate505inter7, gate505inter8, gate505inter9, gate505inter10, gate505inter11, gate505inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate196inter0, gate196inter1, gate196inter2, gate196inter3, gate196inter4, gate196inter5, gate196inter6, gate196inter7, gate196inter8, gate196inter9, gate196inter10, gate196inter11, gate196inter12, gate212inter0, gate212inter1, gate212inter2, gate212inter3, gate212inter4, gate212inter5, gate212inter6, gate212inter7, gate212inter8, gate212inter9, gate212inter10, gate212inter11, gate212inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate395inter0, gate395inter1, gate395inter2, gate395inter3, gate395inter4, gate395inter5, gate395inter6, gate395inter7, gate395inter8, gate395inter9, gate395inter10, gate395inter11, gate395inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate246inter0, gate246inter1, gate246inter2, gate246inter3, gate246inter4, gate246inter5, gate246inter6, gate246inter7, gate246inter8, gate246inter9, gate246inter10, gate246inter11, gate246inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate79inter0, gate79inter1, gate79inter2, gate79inter3, gate79inter4, gate79inter5, gate79inter6, gate79inter7, gate79inter8, gate79inter9, gate79inter10, gate79inter11, gate79inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate421inter0, gate421inter1, gate421inter2, gate421inter3, gate421inter4, gate421inter5, gate421inter6, gate421inter7, gate421inter8, gate421inter9, gate421inter10, gate421inter11, gate421inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );

  xor2  gate729(.a(G6), .b(G5), .O(gate11inter0));
  nand2 gate730(.a(gate11inter0), .b(s_26), .O(gate11inter1));
  and2  gate731(.a(G6), .b(G5), .O(gate11inter2));
  inv1  gate732(.a(s_26), .O(gate11inter3));
  inv1  gate733(.a(s_27), .O(gate11inter4));
  nand2 gate734(.a(gate11inter4), .b(gate11inter3), .O(gate11inter5));
  nor2  gate735(.a(gate11inter5), .b(gate11inter2), .O(gate11inter6));
  inv1  gate736(.a(G5), .O(gate11inter7));
  inv1  gate737(.a(G6), .O(gate11inter8));
  nand2 gate738(.a(gate11inter8), .b(gate11inter7), .O(gate11inter9));
  nand2 gate739(.a(s_27), .b(gate11inter3), .O(gate11inter10));
  nor2  gate740(.a(gate11inter10), .b(gate11inter9), .O(gate11inter11));
  nor2  gate741(.a(gate11inter11), .b(gate11inter6), .O(gate11inter12));
  nand2 gate742(.a(gate11inter12), .b(gate11inter1), .O(G272));
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );

  xor2  gate603(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate604(.a(gate17inter0), .b(s_8), .O(gate17inter1));
  and2  gate605(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate606(.a(s_8), .O(gate17inter3));
  inv1  gate607(.a(s_9), .O(gate17inter4));
  nand2 gate608(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate609(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate610(.a(G17), .O(gate17inter7));
  inv1  gate611(.a(G18), .O(gate17inter8));
  nand2 gate612(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate613(.a(s_9), .b(gate17inter3), .O(gate17inter10));
  nor2  gate614(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate615(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate616(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );

  xor2  gate659(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate660(.a(gate40inter0), .b(s_16), .O(gate40inter1));
  and2  gate661(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate662(.a(s_16), .O(gate40inter3));
  inv1  gate663(.a(s_17), .O(gate40inter4));
  nand2 gate664(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate665(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate666(.a(G28), .O(gate40inter7));
  inv1  gate667(.a(G32), .O(gate40inter8));
  nand2 gate668(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate669(.a(s_17), .b(gate40inter3), .O(gate40inter10));
  nor2  gate670(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate671(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate672(.a(gate40inter12), .b(gate40inter1), .O(G359));
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate953(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate954(.a(gate46inter0), .b(s_58), .O(gate46inter1));
  and2  gate955(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate956(.a(s_58), .O(gate46inter3));
  inv1  gate957(.a(s_59), .O(gate46inter4));
  nand2 gate958(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate959(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate960(.a(G6), .O(gate46inter7));
  inv1  gate961(.a(G272), .O(gate46inter8));
  nand2 gate962(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate963(.a(s_59), .b(gate46inter3), .O(gate46inter10));
  nor2  gate964(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate965(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate966(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate799(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate800(.a(gate54inter0), .b(s_36), .O(gate54inter1));
  and2  gate801(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate802(.a(s_36), .O(gate54inter3));
  inv1  gate803(.a(s_37), .O(gate54inter4));
  nand2 gate804(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate805(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate806(.a(G14), .O(gate54inter7));
  inv1  gate807(.a(G284), .O(gate54inter8));
  nand2 gate808(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate809(.a(s_37), .b(gate54inter3), .O(gate54inter10));
  nor2  gate810(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate811(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate812(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );

  xor2  gate1051(.a(G323), .b(G10), .O(gate79inter0));
  nand2 gate1052(.a(gate79inter0), .b(s_72), .O(gate79inter1));
  and2  gate1053(.a(G323), .b(G10), .O(gate79inter2));
  inv1  gate1054(.a(s_72), .O(gate79inter3));
  inv1  gate1055(.a(s_73), .O(gate79inter4));
  nand2 gate1056(.a(gate79inter4), .b(gate79inter3), .O(gate79inter5));
  nor2  gate1057(.a(gate79inter5), .b(gate79inter2), .O(gate79inter6));
  inv1  gate1058(.a(G10), .O(gate79inter7));
  inv1  gate1059(.a(G323), .O(gate79inter8));
  nand2 gate1060(.a(gate79inter8), .b(gate79inter7), .O(gate79inter9));
  nand2 gate1061(.a(s_73), .b(gate79inter3), .O(gate79inter10));
  nor2  gate1062(.a(gate79inter10), .b(gate79inter9), .O(gate79inter11));
  nor2  gate1063(.a(gate79inter11), .b(gate79inter6), .O(gate79inter12));
  nand2 gate1064(.a(gate79inter12), .b(gate79inter1), .O(G400));
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );

  xor2  gate575(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate576(.a(gate100inter0), .b(s_4), .O(gate100inter1));
  and2  gate577(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate578(.a(s_4), .O(gate100inter3));
  inv1  gate579(.a(s_5), .O(gate100inter4));
  nand2 gate580(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate581(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate582(.a(G31), .O(gate100inter7));
  inv1  gate583(.a(G353), .O(gate100inter8));
  nand2 gate584(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate585(.a(s_5), .b(gate100inter3), .O(gate100inter10));
  nor2  gate586(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate587(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate588(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );

  xor2  gate617(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate618(.a(gate106inter0), .b(s_10), .O(gate106inter1));
  and2  gate619(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate620(.a(s_10), .O(gate106inter3));
  inv1  gate621(.a(s_11), .O(gate106inter4));
  nand2 gate622(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate623(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate624(.a(G364), .O(gate106inter7));
  inv1  gate625(.a(G365), .O(gate106inter8));
  nand2 gate626(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate627(.a(s_11), .b(gate106inter3), .O(gate106inter10));
  nor2  gate628(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate629(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate630(.a(gate106inter12), .b(gate106inter1), .O(G429));

  xor2  gate883(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate884(.a(gate107inter0), .b(s_48), .O(gate107inter1));
  and2  gate885(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate886(.a(s_48), .O(gate107inter3));
  inv1  gate887(.a(s_49), .O(gate107inter4));
  nand2 gate888(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate889(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate890(.a(G366), .O(gate107inter7));
  inv1  gate891(.a(G367), .O(gate107inter8));
  nand2 gate892(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate893(.a(s_49), .b(gate107inter3), .O(gate107inter10));
  nor2  gate894(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate895(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate896(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );

  xor2  gate1107(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate1108(.a(gate115inter0), .b(s_80), .O(gate115inter1));
  and2  gate1109(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate1110(.a(s_80), .O(gate115inter3));
  inv1  gate1111(.a(s_81), .O(gate115inter4));
  nand2 gate1112(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate1113(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate1114(.a(G382), .O(gate115inter7));
  inv1  gate1115(.a(G383), .O(gate115inter8));
  nand2 gate1116(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate1117(.a(s_81), .b(gate115inter3), .O(gate115inter10));
  nor2  gate1118(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate1119(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate1120(.a(gate115inter12), .b(gate115inter1), .O(G456));
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );

  xor2  gate841(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate842(.a(gate120inter0), .b(s_42), .O(gate120inter1));
  and2  gate843(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate844(.a(s_42), .O(gate120inter3));
  inv1  gate845(.a(s_43), .O(gate120inter4));
  nand2 gate846(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate847(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate848(.a(G392), .O(gate120inter7));
  inv1  gate849(.a(G393), .O(gate120inter8));
  nand2 gate850(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate851(.a(s_43), .b(gate120inter3), .O(gate120inter10));
  nor2  gate852(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate853(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate854(.a(gate120inter12), .b(gate120inter1), .O(G471));
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );

  xor2  gate911(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate912(.a(gate131inter0), .b(s_52), .O(gate131inter1));
  and2  gate913(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate914(.a(s_52), .O(gate131inter3));
  inv1  gate915(.a(s_53), .O(gate131inter4));
  nand2 gate916(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate917(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate918(.a(G414), .O(gate131inter7));
  inv1  gate919(.a(G415), .O(gate131inter8));
  nand2 gate920(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate921(.a(s_53), .b(gate131inter3), .O(gate131inter10));
  nor2  gate922(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate923(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate924(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate561(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate562(.a(gate136inter0), .b(s_2), .O(gate136inter1));
  and2  gate563(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate564(.a(s_2), .O(gate136inter3));
  inv1  gate565(.a(s_3), .O(gate136inter4));
  nand2 gate566(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate567(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate568(.a(G424), .O(gate136inter7));
  inv1  gate569(.a(G425), .O(gate136inter8));
  nand2 gate570(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate571(.a(s_3), .b(gate136inter3), .O(gate136inter10));
  nor2  gate572(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate573(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate574(.a(gate136inter12), .b(gate136inter1), .O(G519));
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate1093(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1094(.a(gate148inter0), .b(s_78), .O(gate148inter1));
  and2  gate1095(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1096(.a(s_78), .O(gate148inter3));
  inv1  gate1097(.a(s_79), .O(gate148inter4));
  nand2 gate1098(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1099(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1100(.a(G492), .O(gate148inter7));
  inv1  gate1101(.a(G495), .O(gate148inter8));
  nand2 gate1102(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1103(.a(s_79), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1104(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1105(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1106(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );

  xor2  gate967(.a(G573), .b(G572), .O(gate186inter0));
  nand2 gate968(.a(gate186inter0), .b(s_60), .O(gate186inter1));
  and2  gate969(.a(G573), .b(G572), .O(gate186inter2));
  inv1  gate970(.a(s_60), .O(gate186inter3));
  inv1  gate971(.a(s_61), .O(gate186inter4));
  nand2 gate972(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate973(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate974(.a(G572), .O(gate186inter7));
  inv1  gate975(.a(G573), .O(gate186inter8));
  nand2 gate976(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate977(.a(s_61), .b(gate186inter3), .O(gate186inter10));
  nor2  gate978(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate979(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate980(.a(gate186inter12), .b(gate186inter1), .O(G607));
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );

  xor2  gate855(.a(G593), .b(G592), .O(gate196inter0));
  nand2 gate856(.a(gate196inter0), .b(s_44), .O(gate196inter1));
  and2  gate857(.a(G593), .b(G592), .O(gate196inter2));
  inv1  gate858(.a(s_44), .O(gate196inter3));
  inv1  gate859(.a(s_45), .O(gate196inter4));
  nand2 gate860(.a(gate196inter4), .b(gate196inter3), .O(gate196inter5));
  nor2  gate861(.a(gate196inter5), .b(gate196inter2), .O(gate196inter6));
  inv1  gate862(.a(G592), .O(gate196inter7));
  inv1  gate863(.a(G593), .O(gate196inter8));
  nand2 gate864(.a(gate196inter8), .b(gate196inter7), .O(gate196inter9));
  nand2 gate865(.a(s_45), .b(gate196inter3), .O(gate196inter10));
  nor2  gate866(.a(gate196inter10), .b(gate196inter9), .O(gate196inter11));
  nor2  gate867(.a(gate196inter11), .b(gate196inter6), .O(gate196inter12));
  nand2 gate868(.a(gate196inter12), .b(gate196inter1), .O(G651));
nand2 gate197( .a(G594), .b(G595), .O(G654) );
nand2 gate198( .a(G596), .b(G597), .O(G657) );
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );

  xor2  gate631(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate632(.a(gate201inter0), .b(s_12), .O(gate201inter1));
  and2  gate633(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate634(.a(s_12), .O(gate201inter3));
  inv1  gate635(.a(s_13), .O(gate201inter4));
  nand2 gate636(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate637(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate638(.a(G602), .O(gate201inter7));
  inv1  gate639(.a(G607), .O(gate201inter8));
  nand2 gate640(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate641(.a(s_13), .b(gate201inter3), .O(gate201inter10));
  nor2  gate642(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate643(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate644(.a(gate201inter12), .b(gate201inter1), .O(G666));
nand2 gate202( .a(G612), .b(G617), .O(G669) );
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate1079(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate1080(.a(gate206inter0), .b(s_76), .O(gate206inter1));
  and2  gate1081(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate1082(.a(s_76), .O(gate206inter3));
  inv1  gate1083(.a(s_77), .O(gate206inter4));
  nand2 gate1084(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate1085(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate1086(.a(G632), .O(gate206inter7));
  inv1  gate1087(.a(G637), .O(gate206inter8));
  nand2 gate1088(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate1089(.a(s_77), .b(gate206inter3), .O(gate206inter10));
  nor2  gate1090(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate1091(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate1092(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );

  xor2  gate547(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate548(.a(gate211inter0), .b(s_0), .O(gate211inter1));
  and2  gate549(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate550(.a(s_0), .O(gate211inter3));
  inv1  gate551(.a(s_1), .O(gate211inter4));
  nand2 gate552(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate553(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate554(.a(G612), .O(gate211inter7));
  inv1  gate555(.a(G669), .O(gate211inter8));
  nand2 gate556(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate557(.a(s_1), .b(gate211inter3), .O(gate211inter10));
  nor2  gate558(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate559(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate560(.a(gate211inter12), .b(gate211inter1), .O(G692));

  xor2  gate869(.a(G669), .b(G617), .O(gate212inter0));
  nand2 gate870(.a(gate212inter0), .b(s_46), .O(gate212inter1));
  and2  gate871(.a(G669), .b(G617), .O(gate212inter2));
  inv1  gate872(.a(s_46), .O(gate212inter3));
  inv1  gate873(.a(s_47), .O(gate212inter4));
  nand2 gate874(.a(gate212inter4), .b(gate212inter3), .O(gate212inter5));
  nor2  gate875(.a(gate212inter5), .b(gate212inter2), .O(gate212inter6));
  inv1  gate876(.a(G617), .O(gate212inter7));
  inv1  gate877(.a(G669), .O(gate212inter8));
  nand2 gate878(.a(gate212inter8), .b(gate212inter7), .O(gate212inter9));
  nand2 gate879(.a(s_47), .b(gate212inter3), .O(gate212inter10));
  nor2  gate880(.a(gate212inter10), .b(gate212inter9), .O(gate212inter11));
  nor2  gate881(.a(gate212inter11), .b(gate212inter6), .O(gate212inter12));
  nand2 gate882(.a(gate212inter12), .b(gate212inter1), .O(G693));

  xor2  gate645(.a(G672), .b(G602), .O(gate213inter0));
  nand2 gate646(.a(gate213inter0), .b(s_14), .O(gate213inter1));
  and2  gate647(.a(G672), .b(G602), .O(gate213inter2));
  inv1  gate648(.a(s_14), .O(gate213inter3));
  inv1  gate649(.a(s_15), .O(gate213inter4));
  nand2 gate650(.a(gate213inter4), .b(gate213inter3), .O(gate213inter5));
  nor2  gate651(.a(gate213inter5), .b(gate213inter2), .O(gate213inter6));
  inv1  gate652(.a(G602), .O(gate213inter7));
  inv1  gate653(.a(G672), .O(gate213inter8));
  nand2 gate654(.a(gate213inter8), .b(gate213inter7), .O(gate213inter9));
  nand2 gate655(.a(s_15), .b(gate213inter3), .O(gate213inter10));
  nor2  gate656(.a(gate213inter10), .b(gate213inter9), .O(gate213inter11));
  nor2  gate657(.a(gate213inter11), .b(gate213inter6), .O(gate213inter12));
  nand2 gate658(.a(gate213inter12), .b(gate213inter1), .O(G694));
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );

  xor2  gate673(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate674(.a(gate221inter0), .b(s_18), .O(gate221inter1));
  and2  gate675(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate676(.a(s_18), .O(gate221inter3));
  inv1  gate677(.a(s_19), .O(gate221inter4));
  nand2 gate678(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate679(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate680(.a(G622), .O(gate221inter7));
  inv1  gate681(.a(G684), .O(gate221inter8));
  nand2 gate682(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate683(.a(s_19), .b(gate221inter3), .O(gate221inter10));
  nor2  gate684(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate685(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate686(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );

  xor2  gate1023(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate1024(.a(gate223inter0), .b(s_68), .O(gate223inter1));
  and2  gate1025(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate1026(.a(s_68), .O(gate223inter3));
  inv1  gate1027(.a(s_69), .O(gate223inter4));
  nand2 gate1028(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate1029(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate1030(.a(G627), .O(gate223inter7));
  inv1  gate1031(.a(G687), .O(gate223inter8));
  nand2 gate1032(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate1033(.a(s_69), .b(gate223inter3), .O(gate223inter10));
  nor2  gate1034(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate1035(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate1036(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );

  xor2  gate939(.a(G736), .b(G724), .O(gate246inter0));
  nand2 gate940(.a(gate246inter0), .b(s_56), .O(gate246inter1));
  and2  gate941(.a(G736), .b(G724), .O(gate246inter2));
  inv1  gate942(.a(s_56), .O(gate246inter3));
  inv1  gate943(.a(s_57), .O(gate246inter4));
  nand2 gate944(.a(gate246inter4), .b(gate246inter3), .O(gate246inter5));
  nor2  gate945(.a(gate246inter5), .b(gate246inter2), .O(gate246inter6));
  inv1  gate946(.a(G724), .O(gate246inter7));
  inv1  gate947(.a(G736), .O(gate246inter8));
  nand2 gate948(.a(gate246inter8), .b(gate246inter7), .O(gate246inter9));
  nand2 gate949(.a(s_57), .b(gate246inter3), .O(gate246inter10));
  nor2  gate950(.a(gate246inter10), .b(gate246inter9), .O(gate246inter11));
  nor2  gate951(.a(gate246inter11), .b(gate246inter6), .O(gate246inter12));
  nand2 gate952(.a(gate246inter12), .b(gate246inter1), .O(G759));
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );

  xor2  gate1177(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate1178(.a(gate254inter0), .b(s_90), .O(gate254inter1));
  and2  gate1179(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate1180(.a(s_90), .O(gate254inter3));
  inv1  gate1181(.a(s_91), .O(gate254inter4));
  nand2 gate1182(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate1183(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate1184(.a(G712), .O(gate254inter7));
  inv1  gate1185(.a(G748), .O(gate254inter8));
  nand2 gate1186(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate1187(.a(s_91), .b(gate254inter3), .O(gate254inter10));
  nor2  gate1188(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate1189(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate1190(.a(gate254inter12), .b(gate254inter1), .O(G767));
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate995(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate996(.a(gate258inter0), .b(s_64), .O(gate258inter1));
  and2  gate997(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate998(.a(s_64), .O(gate258inter3));
  inv1  gate999(.a(s_65), .O(gate258inter4));
  nand2 gate1000(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate1001(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate1002(.a(G756), .O(gate258inter7));
  inv1  gate1003(.a(G757), .O(gate258inter8));
  nand2 gate1004(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate1005(.a(s_65), .b(gate258inter3), .O(gate258inter10));
  nor2  gate1006(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate1007(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate1008(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );

  xor2  gate827(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate828(.a(gate277inter0), .b(s_40), .O(gate277inter1));
  and2  gate829(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate830(.a(s_40), .O(gate277inter3));
  inv1  gate831(.a(s_41), .O(gate277inter4));
  nand2 gate832(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate833(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate834(.a(G648), .O(gate277inter7));
  inv1  gate835(.a(G800), .O(gate277inter8));
  nand2 gate836(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate837(.a(s_41), .b(gate277inter3), .O(gate277inter10));
  nor2  gate838(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate839(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate840(.a(gate277inter12), .b(gate277inter1), .O(G822));
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );

  xor2  gate687(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate688(.a(gate286inter0), .b(s_20), .O(gate286inter1));
  and2  gate689(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate690(.a(s_20), .O(gate286inter3));
  inv1  gate691(.a(s_21), .O(gate286inter4));
  nand2 gate692(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate693(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate694(.a(G788), .O(gate286inter7));
  inv1  gate695(.a(G812), .O(gate286inter8));
  nand2 gate696(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate697(.a(s_21), .b(gate286inter3), .O(gate286inter10));
  nor2  gate698(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate699(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate700(.a(gate286inter12), .b(gate286inter1), .O(G831));
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate1009(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate1010(.a(gate291inter0), .b(s_66), .O(gate291inter1));
  and2  gate1011(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate1012(.a(s_66), .O(gate291inter3));
  inv1  gate1013(.a(s_67), .O(gate291inter4));
  nand2 gate1014(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate1015(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate1016(.a(G822), .O(gate291inter7));
  inv1  gate1017(.a(G823), .O(gate291inter8));
  nand2 gate1018(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate1019(.a(s_67), .b(gate291inter3), .O(gate291inter10));
  nor2  gate1020(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate1021(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate1022(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );

  xor2  gate897(.a(G1060), .b(G9), .O(gate395inter0));
  nand2 gate898(.a(gate395inter0), .b(s_50), .O(gate395inter1));
  and2  gate899(.a(G1060), .b(G9), .O(gate395inter2));
  inv1  gate900(.a(s_50), .O(gate395inter3));
  inv1  gate901(.a(s_51), .O(gate395inter4));
  nand2 gate902(.a(gate395inter4), .b(gate395inter3), .O(gate395inter5));
  nor2  gate903(.a(gate395inter5), .b(gate395inter2), .O(gate395inter6));
  inv1  gate904(.a(G9), .O(gate395inter7));
  inv1  gate905(.a(G1060), .O(gate395inter8));
  nand2 gate906(.a(gate395inter8), .b(gate395inter7), .O(gate395inter9));
  nand2 gate907(.a(s_51), .b(gate395inter3), .O(gate395inter10));
  nor2  gate908(.a(gate395inter10), .b(gate395inter9), .O(gate395inter11));
  nor2  gate909(.a(gate395inter11), .b(gate395inter6), .O(gate395inter12));
  nand2 gate910(.a(gate395inter12), .b(gate395inter1), .O(G1156));
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate1121(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate1122(.a(gate397inter0), .b(s_82), .O(gate397inter1));
  and2  gate1123(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate1124(.a(s_82), .O(gate397inter3));
  inv1  gate1125(.a(s_83), .O(gate397inter4));
  nand2 gate1126(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate1127(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate1128(.a(G11), .O(gate397inter7));
  inv1  gate1129(.a(G1066), .O(gate397inter8));
  nand2 gate1130(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate1131(.a(s_83), .b(gate397inter3), .O(gate397inter10));
  nor2  gate1132(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate1133(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate1134(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate701(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate702(.a(gate400inter0), .b(s_22), .O(gate400inter1));
  and2  gate703(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate704(.a(s_22), .O(gate400inter3));
  inv1  gate705(.a(s_23), .O(gate400inter4));
  nand2 gate706(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate707(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate708(.a(G14), .O(gate400inter7));
  inv1  gate709(.a(G1075), .O(gate400inter8));
  nand2 gate710(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate711(.a(s_23), .b(gate400inter3), .O(gate400inter10));
  nor2  gate712(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate713(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate714(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate1163(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate1164(.a(gate415inter0), .b(s_88), .O(gate415inter1));
  and2  gate1165(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate1166(.a(s_88), .O(gate415inter3));
  inv1  gate1167(.a(s_89), .O(gate415inter4));
  nand2 gate1168(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate1169(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate1170(.a(G29), .O(gate415inter7));
  inv1  gate1171(.a(G1120), .O(gate415inter8));
  nand2 gate1172(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate1173(.a(s_89), .b(gate415inter3), .O(gate415inter10));
  nor2  gate1174(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate1175(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate1176(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate743(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate744(.a(gate420inter0), .b(s_28), .O(gate420inter1));
  and2  gate745(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate746(.a(s_28), .O(gate420inter3));
  inv1  gate747(.a(s_29), .O(gate420inter4));
  nand2 gate748(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate749(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate750(.a(G1036), .O(gate420inter7));
  inv1  gate751(.a(G1132), .O(gate420inter8));
  nand2 gate752(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate753(.a(s_29), .b(gate420inter3), .O(gate420inter10));
  nor2  gate754(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate755(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate756(.a(gate420inter12), .b(gate420inter1), .O(G1229));

  xor2  gate1135(.a(G1135), .b(G2), .O(gate421inter0));
  nand2 gate1136(.a(gate421inter0), .b(s_84), .O(gate421inter1));
  and2  gate1137(.a(G1135), .b(G2), .O(gate421inter2));
  inv1  gate1138(.a(s_84), .O(gate421inter3));
  inv1  gate1139(.a(s_85), .O(gate421inter4));
  nand2 gate1140(.a(gate421inter4), .b(gate421inter3), .O(gate421inter5));
  nor2  gate1141(.a(gate421inter5), .b(gate421inter2), .O(gate421inter6));
  inv1  gate1142(.a(G2), .O(gate421inter7));
  inv1  gate1143(.a(G1135), .O(gate421inter8));
  nand2 gate1144(.a(gate421inter8), .b(gate421inter7), .O(gate421inter9));
  nand2 gate1145(.a(s_85), .b(gate421inter3), .O(gate421inter10));
  nor2  gate1146(.a(gate421inter10), .b(gate421inter9), .O(gate421inter11));
  nor2  gate1147(.a(gate421inter11), .b(gate421inter6), .O(gate421inter12));
  nand2 gate1148(.a(gate421inter12), .b(gate421inter1), .O(G1230));
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );

  xor2  gate785(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate786(.a(gate452inter0), .b(s_34), .O(gate452inter1));
  and2  gate787(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate788(.a(s_34), .O(gate452inter3));
  inv1  gate789(.a(s_35), .O(gate452inter4));
  nand2 gate790(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate791(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate792(.a(G1084), .O(gate452inter7));
  inv1  gate793(.a(G1180), .O(gate452inter8));
  nand2 gate794(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate795(.a(s_35), .b(gate452inter3), .O(gate452inter10));
  nor2  gate796(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate797(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate798(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );

  xor2  gate715(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate716(.a(gate458inter0), .b(s_24), .O(gate458inter1));
  and2  gate717(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate718(.a(s_24), .O(gate458inter3));
  inv1  gate719(.a(s_25), .O(gate458inter4));
  nand2 gate720(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate721(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate722(.a(G1093), .O(gate458inter7));
  inv1  gate723(.a(G1189), .O(gate458inter8));
  nand2 gate724(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate725(.a(s_25), .b(gate458inter3), .O(gate458inter10));
  nor2  gate726(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate727(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate728(.a(gate458inter12), .b(gate458inter1), .O(G1267));
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );

  xor2  gate981(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate982(.a(gate465inter0), .b(s_62), .O(gate465inter1));
  and2  gate983(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate984(.a(s_62), .O(gate465inter3));
  inv1  gate985(.a(s_63), .O(gate465inter4));
  nand2 gate986(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate987(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate988(.a(G24), .O(gate465inter7));
  inv1  gate989(.a(G1201), .O(gate465inter8));
  nand2 gate990(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate991(.a(s_63), .b(gate465inter3), .O(gate465inter10));
  nor2  gate992(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate993(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate994(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate1149(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate1150(.a(gate471inter0), .b(s_86), .O(gate471inter1));
  and2  gate1151(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate1152(.a(s_86), .O(gate471inter3));
  inv1  gate1153(.a(s_87), .O(gate471inter4));
  nand2 gate1154(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate1155(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate1156(.a(G27), .O(gate471inter7));
  inv1  gate1157(.a(G1210), .O(gate471inter8));
  nand2 gate1158(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate1159(.a(s_87), .b(gate471inter3), .O(gate471inter10));
  nor2  gate1160(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate1161(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate1162(.a(gate471inter12), .b(gate471inter1), .O(G1280));
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );

  xor2  gate771(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate772(.a(gate478inter0), .b(s_32), .O(gate478inter1));
  and2  gate773(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate774(.a(s_32), .O(gate478inter3));
  inv1  gate775(.a(s_33), .O(gate478inter4));
  nand2 gate776(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate777(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate778(.a(G1123), .O(gate478inter7));
  inv1  gate779(.a(G1219), .O(gate478inter8));
  nand2 gate780(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate781(.a(s_33), .b(gate478inter3), .O(gate478inter10));
  nor2  gate782(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate783(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate784(.a(gate478inter12), .b(gate478inter1), .O(G1287));
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );

  xor2  gate589(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate590(.a(gate484inter0), .b(s_6), .O(gate484inter1));
  and2  gate591(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate592(.a(s_6), .O(gate484inter3));
  inv1  gate593(.a(s_7), .O(gate484inter4));
  nand2 gate594(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate595(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate596(.a(G1230), .O(gate484inter7));
  inv1  gate597(.a(G1231), .O(gate484inter8));
  nand2 gate598(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate599(.a(s_7), .b(gate484inter3), .O(gate484inter10));
  nor2  gate600(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate601(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate602(.a(gate484inter12), .b(gate484inter1), .O(G1293));
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate925(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate926(.a(gate490inter0), .b(s_54), .O(gate490inter1));
  and2  gate927(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate928(.a(s_54), .O(gate490inter3));
  inv1  gate929(.a(s_55), .O(gate490inter4));
  nand2 gate930(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate931(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate932(.a(G1242), .O(gate490inter7));
  inv1  gate933(.a(G1243), .O(gate490inter8));
  nand2 gate934(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate935(.a(s_55), .b(gate490inter3), .O(gate490inter10));
  nor2  gate936(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate937(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate938(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate1065(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate1066(.a(gate504inter0), .b(s_74), .O(gate504inter1));
  and2  gate1067(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate1068(.a(s_74), .O(gate504inter3));
  inv1  gate1069(.a(s_75), .O(gate504inter4));
  nand2 gate1070(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate1071(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate1072(.a(G1270), .O(gate504inter7));
  inv1  gate1073(.a(G1271), .O(gate504inter8));
  nand2 gate1074(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate1075(.a(s_75), .b(gate504inter3), .O(gate504inter10));
  nor2  gate1076(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate1077(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate1078(.a(gate504inter12), .b(gate504inter1), .O(G1313));

  xor2  gate757(.a(G1273), .b(G1272), .O(gate505inter0));
  nand2 gate758(.a(gate505inter0), .b(s_30), .O(gate505inter1));
  and2  gate759(.a(G1273), .b(G1272), .O(gate505inter2));
  inv1  gate760(.a(s_30), .O(gate505inter3));
  inv1  gate761(.a(s_31), .O(gate505inter4));
  nand2 gate762(.a(gate505inter4), .b(gate505inter3), .O(gate505inter5));
  nor2  gate763(.a(gate505inter5), .b(gate505inter2), .O(gate505inter6));
  inv1  gate764(.a(G1272), .O(gate505inter7));
  inv1  gate765(.a(G1273), .O(gate505inter8));
  nand2 gate766(.a(gate505inter8), .b(gate505inter7), .O(gate505inter9));
  nand2 gate767(.a(s_31), .b(gate505inter3), .O(gate505inter10));
  nor2  gate768(.a(gate505inter10), .b(gate505inter9), .O(gate505inter11));
  nor2  gate769(.a(gate505inter11), .b(gate505inter6), .O(gate505inter12));
  nand2 gate770(.a(gate505inter12), .b(gate505inter1), .O(G1314));

  xor2  gate813(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate814(.a(gate506inter0), .b(s_38), .O(gate506inter1));
  and2  gate815(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate816(.a(s_38), .O(gate506inter3));
  inv1  gate817(.a(s_39), .O(gate506inter4));
  nand2 gate818(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate819(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate820(.a(G1274), .O(gate506inter7));
  inv1  gate821(.a(G1275), .O(gate506inter8));
  nand2 gate822(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate823(.a(s_39), .b(gate506inter3), .O(gate506inter10));
  nor2  gate824(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate825(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate826(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate1037(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate1038(.a(gate510inter0), .b(s_70), .O(gate510inter1));
  and2  gate1039(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate1040(.a(s_70), .O(gate510inter3));
  inv1  gate1041(.a(s_71), .O(gate510inter4));
  nand2 gate1042(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate1043(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate1044(.a(G1282), .O(gate510inter7));
  inv1  gate1045(.a(G1283), .O(gate510inter8));
  nand2 gate1046(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate1047(.a(s_71), .b(gate510inter3), .O(gate510inter10));
  nor2  gate1048(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate1049(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate1050(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule