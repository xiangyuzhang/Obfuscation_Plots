module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251, s_252, s_253, s_254, s_255, s_256, s_257, s_258, s_259, s_260, s_261, s_262, s_263, s_264, s_265, s_266, s_267, s_268, s_269, s_270, s_271, s_272, s_273, s_274, s_275, s_276, s_277, s_278, s_279, s_280, s_281, s_282, s_283, s_284, s_285, s_286, s_287, s_288, s_289, s_290, s_291, s_292, s_293, s_294, s_295, s_296, s_297, s_298, s_299, s_300, s_301, s_302, s_303, s_304, s_305, s_306, s_307, s_308, s_309, s_310, s_311, s_312, s_313, s_314, s_315, s_316, s_317, s_318, s_319, s_320, s_321, s_322, s_323, s_324, s_325, s_326, s_327, s_328, s_329, s_330, s_331, s_332, s_333, s_334, s_335, s_336, s_337, s_338, s_339, s_340, s_341, s_342, s_343, s_344, s_345, s_346, s_347, s_348, s_349, s_350, s_351, s_352, s_353, s_354, s_355, s_356, s_357, s_358, s_359, s_360, s_361;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate74inter0, gate74inter1, gate74inter2, gate74inter3, gate74inter4, gate74inter5, gate74inter6, gate74inter7, gate74inter8, gate74inter9, gate74inter10, gate74inter11, gate74inter12, gate286inter0, gate286inter1, gate286inter2, gate286inter3, gate286inter4, gate286inter5, gate286inter6, gate286inter7, gate286inter8, gate286inter9, gate286inter10, gate286inter11, gate286inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate124inter0, gate124inter1, gate124inter2, gate124inter3, gate124inter4, gate124inter5, gate124inter6, gate124inter7, gate124inter8, gate124inter9, gate124inter10, gate124inter11, gate124inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate141inter0, gate141inter1, gate141inter2, gate141inter3, gate141inter4, gate141inter5, gate141inter6, gate141inter7, gate141inter8, gate141inter9, gate141inter10, gate141inter11, gate141inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate23inter0, gate23inter1, gate23inter2, gate23inter3, gate23inter4, gate23inter5, gate23inter6, gate23inter7, gate23inter8, gate23inter9, gate23inter10, gate23inter11, gate23inter12, gate51inter0, gate51inter1, gate51inter2, gate51inter3, gate51inter4, gate51inter5, gate51inter6, gate51inter7, gate51inter8, gate51inter9, gate51inter10, gate51inter11, gate51inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate228inter0, gate228inter1, gate228inter2, gate228inter3, gate228inter4, gate228inter5, gate228inter6, gate228inter7, gate228inter8, gate228inter9, gate228inter10, gate228inter11, gate228inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate182inter0, gate182inter1, gate182inter2, gate182inter3, gate182inter4, gate182inter5, gate182inter6, gate182inter7, gate182inter8, gate182inter9, gate182inter10, gate182inter11, gate182inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate506inter0, gate506inter1, gate506inter2, gate506inter3, gate506inter4, gate506inter5, gate506inter6, gate506inter7, gate506inter8, gate506inter9, gate506inter10, gate506inter11, gate506inter12, gate498inter0, gate498inter1, gate498inter2, gate498inter3, gate498inter4, gate498inter5, gate498inter6, gate498inter7, gate498inter8, gate498inter9, gate498inter10, gate498inter11, gate498inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate432inter0, gate432inter1, gate432inter2, gate432inter3, gate432inter4, gate432inter5, gate432inter6, gate432inter7, gate432inter8, gate432inter9, gate432inter10, gate432inter11, gate432inter12, gate201inter0, gate201inter1, gate201inter2, gate201inter3, gate201inter4, gate201inter5, gate201inter6, gate201inter7, gate201inter8, gate201inter9, gate201inter10, gate201inter11, gate201inter12, gate39inter0, gate39inter1, gate39inter2, gate39inter3, gate39inter4, gate39inter5, gate39inter6, gate39inter7, gate39inter8, gate39inter9, gate39inter10, gate39inter11, gate39inter12, gate208inter0, gate208inter1, gate208inter2, gate208inter3, gate208inter4, gate208inter5, gate208inter6, gate208inter7, gate208inter8, gate208inter9, gate208inter10, gate208inter11, gate208inter12, gate248inter0, gate248inter1, gate248inter2, gate248inter3, gate248inter4, gate248inter5, gate248inter6, gate248inter7, gate248inter8, gate248inter9, gate248inter10, gate248inter11, gate248inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate223inter0, gate223inter1, gate223inter2, gate223inter3, gate223inter4, gate223inter5, gate223inter6, gate223inter7, gate223inter8, gate223inter9, gate223inter10, gate223inter11, gate223inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate115inter0, gate115inter1, gate115inter2, gate115inter3, gate115inter4, gate115inter5, gate115inter6, gate115inter7, gate115inter8, gate115inter9, gate115inter10, gate115inter11, gate115inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate509inter0, gate509inter1, gate509inter2, gate509inter3, gate509inter4, gate509inter5, gate509inter6, gate509inter7, gate509inter8, gate509inter9, gate509inter10, gate509inter11, gate509inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate187inter0, gate187inter1, gate187inter2, gate187inter3, gate187inter4, gate187inter5, gate187inter6, gate187inter7, gate187inter8, gate187inter9, gate187inter10, gate187inter11, gate187inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate255inter0, gate255inter1, gate255inter2, gate255inter3, gate255inter4, gate255inter5, gate255inter6, gate255inter7, gate255inter8, gate255inter9, gate255inter10, gate255inter11, gate255inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate167inter0, gate167inter1, gate167inter2, gate167inter3, gate167inter4, gate167inter5, gate167inter6, gate167inter7, gate167inter8, gate167inter9, gate167inter10, gate167inter11, gate167inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate100inter0, gate100inter1, gate100inter2, gate100inter3, gate100inter4, gate100inter5, gate100inter6, gate100inter7, gate100inter8, gate100inter9, gate100inter10, gate100inter11, gate100inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate207inter0, gate207inter1, gate207inter2, gate207inter3, gate207inter4, gate207inter5, gate207inter6, gate207inter7, gate207inter8, gate207inter9, gate207inter10, gate207inter11, gate207inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate457inter0, gate457inter1, gate457inter2, gate457inter3, gate457inter4, gate457inter5, gate457inter6, gate457inter7, gate457inter8, gate457inter9, gate457inter10, gate457inter11, gate457inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate102inter0, gate102inter1, gate102inter2, gate102inter3, gate102inter4, gate102inter5, gate102inter6, gate102inter7, gate102inter8, gate102inter9, gate102inter10, gate102inter11, gate102inter12, gate388inter0, gate388inter1, gate388inter2, gate388inter3, gate388inter4, gate388inter5, gate388inter6, gate388inter7, gate388inter8, gate388inter9, gate388inter10, gate388inter11, gate388inter12, gate283inter0, gate283inter1, gate283inter2, gate283inter3, gate283inter4, gate283inter5, gate283inter6, gate283inter7, gate283inter8, gate283inter9, gate283inter10, gate283inter11, gate283inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate143inter0, gate143inter1, gate143inter2, gate143inter3, gate143inter4, gate143inter5, gate143inter6, gate143inter7, gate143inter8, gate143inter9, gate143inter10, gate143inter11, gate143inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate222inter0, gate222inter1, gate222inter2, gate222inter3, gate222inter4, gate222inter5, gate222inter6, gate222inter7, gate222inter8, gate222inter9, gate222inter10, gate222inter11, gate222inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate405inter0, gate405inter1, gate405inter2, gate405inter3, gate405inter4, gate405inter5, gate405inter6, gate405inter7, gate405inter8, gate405inter9, gate405inter10, gate405inter11, gate405inter12, gate55inter0, gate55inter1, gate55inter2, gate55inter3, gate55inter4, gate55inter5, gate55inter6, gate55inter7, gate55inter8, gate55inter9, gate55inter10, gate55inter11, gate55inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate428inter0, gate428inter1, gate428inter2, gate428inter3, gate428inter4, gate428inter5, gate428inter6, gate428inter7, gate428inter8, gate428inter9, gate428inter10, gate428inter11, gate428inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate130inter0, gate130inter1, gate130inter2, gate130inter3, gate130inter4, gate130inter5, gate130inter6, gate130inter7, gate130inter8, gate130inter9, gate130inter10, gate130inter11, gate130inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate271inter0, gate271inter1, gate271inter2, gate271inter3, gate271inter4, gate271inter5, gate271inter6, gate271inter7, gate271inter8, gate271inter9, gate271inter10, gate271inter11, gate271inter12, gate185inter0, gate185inter1, gate185inter2, gate185inter3, gate185inter4, gate185inter5, gate185inter6, gate185inter7, gate185inter8, gate185inter9, gate185inter10, gate185inter11, gate185inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate512inter0, gate512inter1, gate512inter2, gate512inter3, gate512inter4, gate512inter5, gate512inter6, gate512inter7, gate512inter8, gate512inter9, gate512inter10, gate512inter11, gate512inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate394inter0, gate394inter1, gate394inter2, gate394inter3, gate394inter4, gate394inter5, gate394inter6, gate394inter7, gate394inter8, gate394inter9, gate394inter10, gate394inter11, gate394inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate22inter0, gate22inter1, gate22inter2, gate22inter3, gate22inter4, gate22inter5, gate22inter6, gate22inter7, gate22inter8, gate22inter9, gate22inter10, gate22inter11, gate22inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate90inter0, gate90inter1, gate90inter2, gate90inter3, gate90inter4, gate90inter5, gate90inter6, gate90inter7, gate90inter8, gate90inter9, gate90inter10, gate90inter11, gate90inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate52inter0, gate52inter1, gate52inter2, gate52inter3, gate52inter4, gate52inter5, gate52inter6, gate52inter7, gate52inter8, gate52inter9, gate52inter10, gate52inter11, gate52inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate440inter0, gate440inter1, gate440inter2, gate440inter3, gate440inter4, gate440inter5, gate440inter6, gate440inter7, gate440inter8, gate440inter9, gate440inter10, gate440inter11, gate440inter12, gate139inter0, gate139inter1, gate139inter2, gate139inter3, gate139inter4, gate139inter5, gate139inter6, gate139inter7, gate139inter8, gate139inter9, gate139inter10, gate139inter11, gate139inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate397inter0, gate397inter1, gate397inter2, gate397inter3, gate397inter4, gate397inter5, gate397inter6, gate397inter7, gate397inter8, gate397inter9, gate397inter10, gate397inter11, gate397inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate60inter0, gate60inter1, gate60inter2, gate60inter3, gate60inter4, gate60inter5, gate60inter6, gate60inter7, gate60inter8, gate60inter9, gate60inter10, gate60inter11, gate60inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate500inter0, gate500inter1, gate500inter2, gate500inter3, gate500inter4, gate500inter5, gate500inter6, gate500inter7, gate500inter8, gate500inter9, gate500inter10, gate500inter11, gate500inter12, gate233inter0, gate233inter1, gate233inter2, gate233inter3, gate233inter4, gate233inter5, gate233inter6, gate233inter7, gate233inter8, gate233inter9, gate233inter10, gate233inter11, gate233inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate270inter0, gate270inter1, gate270inter2, gate270inter3, gate270inter4, gate270inter5, gate270inter6, gate270inter7, gate270inter8, gate270inter9, gate270inter10, gate270inter11, gate270inter12, gate104inter0, gate104inter1, gate104inter2, gate104inter3, gate104inter4, gate104inter5, gate104inter6, gate104inter7, gate104inter8, gate104inter9, gate104inter10, gate104inter11, gate104inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate50inter0, gate50inter1, gate50inter2, gate50inter3, gate50inter4, gate50inter5, gate50inter6, gate50inter7, gate50inter8, gate50inter9, gate50inter10, gate50inter11, gate50inter12, gate413inter0, gate413inter1, gate413inter2, gate413inter3, gate413inter4, gate413inter5, gate413inter6, gate413inter7, gate413inter8, gate413inter9, gate413inter10, gate413inter11, gate413inter12, gate131inter0, gate131inter1, gate131inter2, gate131inter3, gate131inter4, gate131inter5, gate131inter6, gate131inter7, gate131inter8, gate131inter9, gate131inter10, gate131inter11, gate131inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate114inter0, gate114inter1, gate114inter2, gate114inter3, gate114inter4, gate114inter5, gate114inter6, gate114inter7, gate114inter8, gate114inter9, gate114inter10, gate114inter11, gate114inter12, gate452inter0, gate452inter1, gate452inter2, gate452inter3, gate452inter4, gate452inter5, gate452inter6, gate452inter7, gate452inter8, gate452inter9, gate452inter10, gate452inter11, gate452inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate56inter0, gate56inter1, gate56inter2, gate56inter3, gate56inter4, gate56inter5, gate56inter6, gate56inter7, gate56inter8, gate56inter9, gate56inter10, gate56inter11, gate56inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate158inter0, gate158inter1, gate158inter2, gate158inter3, gate158inter4, gate158inter5, gate158inter6, gate158inter7, gate158inter8, gate158inter9, gate158inter10, gate158inter11, gate158inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate215inter0, gate215inter1, gate215inter2, gate215inter3, gate215inter4, gate215inter5, gate215inter6, gate215inter7, gate215inter8, gate215inter9, gate215inter10, gate215inter11, gate215inter12, gate157inter0, gate157inter1, gate157inter2, gate157inter3, gate157inter4, gate157inter5, gate157inter6, gate157inter7, gate157inter8, gate157inter9, gate157inter10, gate157inter11, gate157inter12, gate256inter0, gate256inter1, gate256inter2, gate256inter3, gate256inter4, gate256inter5, gate256inter6, gate256inter7, gate256inter8, gate256inter9, gate256inter10, gate256inter11, gate256inter12, gate170inter0, gate170inter1, gate170inter2, gate170inter3, gate170inter4, gate170inter5, gate170inter6, gate170inter7, gate170inter8, gate170inter9, gate170inter10, gate170inter11, gate170inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate230inter0, gate230inter1, gate230inter2, gate230inter3, gate230inter4, gate230inter5, gate230inter6, gate230inter7, gate230inter8, gate230inter9, gate230inter10, gate230inter11, gate230inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate152inter0, gate152inter1, gate152inter2, gate152inter3, gate152inter4, gate152inter5, gate152inter6, gate152inter7, gate152inter8, gate152inter9, gate152inter10, gate152inter11, gate152inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate1387(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate1388(.a(gate9inter0), .b(s_120), .O(gate9inter1));
  and2  gate1389(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate1390(.a(s_120), .O(gate9inter3));
  inv1  gate1391(.a(s_121), .O(gate9inter4));
  nand2 gate1392(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate1393(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate1394(.a(G1), .O(gate9inter7));
  inv1  gate1395(.a(G2), .O(gate9inter8));
  nand2 gate1396(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate1397(.a(s_121), .b(gate9inter3), .O(gate9inter10));
  nor2  gate1398(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate1399(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate1400(.a(gate9inter12), .b(gate9inter1), .O(G266));

  xor2  gate1205(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate1206(.a(gate10inter0), .b(s_94), .O(gate10inter1));
  and2  gate1207(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate1208(.a(s_94), .O(gate10inter3));
  inv1  gate1209(.a(s_95), .O(gate10inter4));
  nand2 gate1210(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate1211(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate1212(.a(G3), .O(gate10inter7));
  inv1  gate1213(.a(G4), .O(gate10inter8));
  nand2 gate1214(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate1215(.a(s_95), .b(gate10inter3), .O(gate10inter10));
  nor2  gate1216(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate1217(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate1218(.a(gate10inter12), .b(gate10inter1), .O(G269));
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate2549(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate2550(.a(gate12inter0), .b(s_286), .O(gate12inter1));
  and2  gate2551(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate2552(.a(s_286), .O(gate12inter3));
  inv1  gate2553(.a(s_287), .O(gate12inter4));
  nand2 gate2554(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate2555(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate2556(.a(G7), .O(gate12inter7));
  inv1  gate2557(.a(G8), .O(gate12inter8));
  nand2 gate2558(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate2559(.a(s_287), .b(gate12inter3), .O(gate12inter10));
  nor2  gate2560(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate2561(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate2562(.a(gate12inter12), .b(gate12inter1), .O(G275));
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate2325(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate2326(.a(gate15inter0), .b(s_254), .O(gate15inter1));
  and2  gate2327(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate2328(.a(s_254), .O(gate15inter3));
  inv1  gate2329(.a(s_255), .O(gate15inter4));
  nand2 gate2330(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate2331(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate2332(.a(G13), .O(gate15inter7));
  inv1  gate2333(.a(G14), .O(gate15inter8));
  nand2 gate2334(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate2335(.a(s_255), .b(gate15inter3), .O(gate15inter10));
  nor2  gate2336(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate2337(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate2338(.a(gate15inter12), .b(gate15inter1), .O(G284));

  xor2  gate1947(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate1948(.a(gate16inter0), .b(s_200), .O(gate16inter1));
  and2  gate1949(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate1950(.a(s_200), .O(gate16inter3));
  inv1  gate1951(.a(s_201), .O(gate16inter4));
  nand2 gate1952(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate1953(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate1954(.a(G15), .O(gate16inter7));
  inv1  gate1955(.a(G16), .O(gate16inter8));
  nand2 gate1956(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate1957(.a(s_201), .b(gate16inter3), .O(gate16inter10));
  nor2  gate1958(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate1959(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate1960(.a(gate16inter12), .b(gate16inter1), .O(G287));
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate631(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate632(.a(gate20inter0), .b(s_12), .O(gate20inter1));
  and2  gate633(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate634(.a(s_12), .O(gate20inter3));
  inv1  gate635(.a(s_13), .O(gate20inter4));
  nand2 gate636(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate637(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate638(.a(G23), .O(gate20inter7));
  inv1  gate639(.a(G24), .O(gate20inter8));
  nand2 gate640(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate641(.a(s_13), .b(gate20inter3), .O(gate20inter10));
  nor2  gate642(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate643(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate644(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );

  xor2  gate2213(.a(G28), .b(G27), .O(gate22inter0));
  nand2 gate2214(.a(gate22inter0), .b(s_238), .O(gate22inter1));
  and2  gate2215(.a(G28), .b(G27), .O(gate22inter2));
  inv1  gate2216(.a(s_238), .O(gate22inter3));
  inv1  gate2217(.a(s_239), .O(gate22inter4));
  nand2 gate2218(.a(gate22inter4), .b(gate22inter3), .O(gate22inter5));
  nor2  gate2219(.a(gate22inter5), .b(gate22inter2), .O(gate22inter6));
  inv1  gate2220(.a(G27), .O(gate22inter7));
  inv1  gate2221(.a(G28), .O(gate22inter8));
  nand2 gate2222(.a(gate22inter8), .b(gate22inter7), .O(gate22inter9));
  nand2 gate2223(.a(s_239), .b(gate22inter3), .O(gate22inter10));
  nor2  gate2224(.a(gate22inter10), .b(gate22inter9), .O(gate22inter11));
  nor2  gate2225(.a(gate22inter11), .b(gate22inter6), .O(gate22inter12));
  nand2 gate2226(.a(gate22inter12), .b(gate22inter1), .O(G305));

  xor2  gate715(.a(G30), .b(G29), .O(gate23inter0));
  nand2 gate716(.a(gate23inter0), .b(s_24), .O(gate23inter1));
  and2  gate717(.a(G30), .b(G29), .O(gate23inter2));
  inv1  gate718(.a(s_24), .O(gate23inter3));
  inv1  gate719(.a(s_25), .O(gate23inter4));
  nand2 gate720(.a(gate23inter4), .b(gate23inter3), .O(gate23inter5));
  nor2  gate721(.a(gate23inter5), .b(gate23inter2), .O(gate23inter6));
  inv1  gate722(.a(G29), .O(gate23inter7));
  inv1  gate723(.a(G30), .O(gate23inter8));
  nand2 gate724(.a(gate23inter8), .b(gate23inter7), .O(gate23inter9));
  nand2 gate725(.a(s_25), .b(gate23inter3), .O(gate23inter10));
  nor2  gate726(.a(gate23inter10), .b(gate23inter9), .O(gate23inter11));
  nor2  gate727(.a(gate23inter11), .b(gate23inter6), .O(gate23inter12));
  nand2 gate728(.a(gate23inter12), .b(gate23inter1), .O(G308));
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate2255(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate2256(.a(gate26inter0), .b(s_244), .O(gate26inter1));
  and2  gate2257(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate2258(.a(s_244), .O(gate26inter3));
  inv1  gate2259(.a(s_245), .O(gate26inter4));
  nand2 gate2260(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate2261(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate2262(.a(G9), .O(gate26inter7));
  inv1  gate2263(.a(G13), .O(gate26inter8));
  nand2 gate2264(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate2265(.a(s_245), .b(gate26inter3), .O(gate26inter10));
  nor2  gate2266(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate2267(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate2268(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate897(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate898(.a(gate29inter0), .b(s_50), .O(gate29inter1));
  and2  gate899(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate900(.a(s_50), .O(gate29inter3));
  inv1  gate901(.a(s_51), .O(gate29inter4));
  nand2 gate902(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate903(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate904(.a(G3), .O(gate29inter7));
  inv1  gate905(.a(G7), .O(gate29inter8));
  nand2 gate906(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate907(.a(s_51), .b(gate29inter3), .O(gate29inter10));
  nor2  gate908(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate909(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate910(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate1443(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate1444(.a(gate37inter0), .b(s_128), .O(gate37inter1));
  and2  gate1445(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate1446(.a(s_128), .O(gate37inter3));
  inv1  gate1447(.a(s_129), .O(gate37inter4));
  nand2 gate1448(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate1449(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate1450(.a(G19), .O(gate37inter7));
  inv1  gate1451(.a(G23), .O(gate37inter8));
  nand2 gate1452(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate1453(.a(s_129), .b(gate37inter3), .O(gate37inter10));
  nor2  gate1454(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate1455(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate1456(.a(gate37inter12), .b(gate37inter1), .O(G350));
nand2 gate38( .a(G27), .b(G31), .O(G353) );

  xor2  gate939(.a(G24), .b(G20), .O(gate39inter0));
  nand2 gate940(.a(gate39inter0), .b(s_56), .O(gate39inter1));
  and2  gate941(.a(G24), .b(G20), .O(gate39inter2));
  inv1  gate942(.a(s_56), .O(gate39inter3));
  inv1  gate943(.a(s_57), .O(gate39inter4));
  nand2 gate944(.a(gate39inter4), .b(gate39inter3), .O(gate39inter5));
  nor2  gate945(.a(gate39inter5), .b(gate39inter2), .O(gate39inter6));
  inv1  gate946(.a(G20), .O(gate39inter7));
  inv1  gate947(.a(G24), .O(gate39inter8));
  nand2 gate948(.a(gate39inter8), .b(gate39inter7), .O(gate39inter9));
  nand2 gate949(.a(s_57), .b(gate39inter3), .O(gate39inter10));
  nor2  gate950(.a(gate39inter10), .b(gate39inter9), .O(gate39inter11));
  nor2  gate951(.a(gate39inter11), .b(gate39inter6), .O(gate39inter12));
  nand2 gate952(.a(gate39inter12), .b(gate39inter1), .O(G356));

  xor2  gate743(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate744(.a(gate40inter0), .b(s_28), .O(gate40inter1));
  and2  gate745(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate746(.a(s_28), .O(gate40inter3));
  inv1  gate747(.a(s_29), .O(gate40inter4));
  nand2 gate748(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate749(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate750(.a(G28), .O(gate40inter7));
  inv1  gate751(.a(G32), .O(gate40inter8));
  nand2 gate752(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate753(.a(s_29), .b(gate40inter3), .O(gate40inter10));
  nor2  gate754(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate755(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate756(.a(gate40inter12), .b(gate40inter1), .O(G359));

  xor2  gate1807(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate1808(.a(gate41inter0), .b(s_180), .O(gate41inter1));
  and2  gate1809(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate1810(.a(s_180), .O(gate41inter3));
  inv1  gate1811(.a(s_181), .O(gate41inter4));
  nand2 gate1812(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate1813(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate1814(.a(G1), .O(gate41inter7));
  inv1  gate1815(.a(G266), .O(gate41inter8));
  nand2 gate1816(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate1817(.a(s_181), .b(gate41inter3), .O(gate41inter10));
  nor2  gate1818(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate1819(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate1820(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate2955(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate2956(.a(gate46inter0), .b(s_344), .O(gate46inter1));
  and2  gate2957(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate2958(.a(s_344), .O(gate46inter3));
  inv1  gate2959(.a(s_345), .O(gate46inter4));
  nand2 gate2960(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate2961(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate2962(.a(G6), .O(gate46inter7));
  inv1  gate2963(.a(G272), .O(gate46inter8));
  nand2 gate2964(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate2965(.a(s_345), .b(gate46inter3), .O(gate46inter10));
  nor2  gate2966(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate2967(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate2968(.a(gate46inter12), .b(gate46inter1), .O(G367));

  xor2  gate841(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate842(.a(gate47inter0), .b(s_42), .O(gate47inter1));
  and2  gate843(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate844(.a(s_42), .O(gate47inter3));
  inv1  gate845(.a(s_43), .O(gate47inter4));
  nand2 gate846(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate847(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate848(.a(G7), .O(gate47inter7));
  inv1  gate849(.a(G275), .O(gate47inter8));
  nand2 gate850(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate851(.a(s_43), .b(gate47inter3), .O(gate47inter10));
  nor2  gate852(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate853(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate854(.a(gate47inter12), .b(gate47inter1), .O(G368));

  xor2  gate1933(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate1934(.a(gate48inter0), .b(s_198), .O(gate48inter1));
  and2  gate1935(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate1936(.a(s_198), .O(gate48inter3));
  inv1  gate1937(.a(s_199), .O(gate48inter4));
  nand2 gate1938(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate1939(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate1940(.a(G8), .O(gate48inter7));
  inv1  gate1941(.a(G275), .O(gate48inter8));
  nand2 gate1942(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate1943(.a(s_199), .b(gate48inter3), .O(gate48inter10));
  nor2  gate1944(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate1945(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate1946(.a(gate48inter12), .b(gate48inter1), .O(G369));
nand2 gate49( .a(G9), .b(G278), .O(G370) );

  xor2  gate2591(.a(G278), .b(G10), .O(gate50inter0));
  nand2 gate2592(.a(gate50inter0), .b(s_292), .O(gate50inter1));
  and2  gate2593(.a(G278), .b(G10), .O(gate50inter2));
  inv1  gate2594(.a(s_292), .O(gate50inter3));
  inv1  gate2595(.a(s_293), .O(gate50inter4));
  nand2 gate2596(.a(gate50inter4), .b(gate50inter3), .O(gate50inter5));
  nor2  gate2597(.a(gate50inter5), .b(gate50inter2), .O(gate50inter6));
  inv1  gate2598(.a(G10), .O(gate50inter7));
  inv1  gate2599(.a(G278), .O(gate50inter8));
  nand2 gate2600(.a(gate50inter8), .b(gate50inter7), .O(gate50inter9));
  nand2 gate2601(.a(s_293), .b(gate50inter3), .O(gate50inter10));
  nor2  gate2602(.a(gate50inter10), .b(gate50inter9), .O(gate50inter11));
  nor2  gate2603(.a(gate50inter11), .b(gate50inter6), .O(gate50inter12));
  nand2 gate2604(.a(gate50inter12), .b(gate50inter1), .O(G371));

  xor2  gate729(.a(G281), .b(G11), .O(gate51inter0));
  nand2 gate730(.a(gate51inter0), .b(s_26), .O(gate51inter1));
  and2  gate731(.a(G281), .b(G11), .O(gate51inter2));
  inv1  gate732(.a(s_26), .O(gate51inter3));
  inv1  gate733(.a(s_27), .O(gate51inter4));
  nand2 gate734(.a(gate51inter4), .b(gate51inter3), .O(gate51inter5));
  nor2  gate735(.a(gate51inter5), .b(gate51inter2), .O(gate51inter6));
  inv1  gate736(.a(G11), .O(gate51inter7));
  inv1  gate737(.a(G281), .O(gate51inter8));
  nand2 gate738(.a(gate51inter8), .b(gate51inter7), .O(gate51inter9));
  nand2 gate739(.a(s_27), .b(gate51inter3), .O(gate51inter10));
  nor2  gate740(.a(gate51inter10), .b(gate51inter9), .O(gate51inter11));
  nor2  gate741(.a(gate51inter11), .b(gate51inter6), .O(gate51inter12));
  nand2 gate742(.a(gate51inter12), .b(gate51inter1), .O(G372));

  xor2  gate2311(.a(G281), .b(G12), .O(gate52inter0));
  nand2 gate2312(.a(gate52inter0), .b(s_252), .O(gate52inter1));
  and2  gate2313(.a(G281), .b(G12), .O(gate52inter2));
  inv1  gate2314(.a(s_252), .O(gate52inter3));
  inv1  gate2315(.a(s_253), .O(gate52inter4));
  nand2 gate2316(.a(gate52inter4), .b(gate52inter3), .O(gate52inter5));
  nor2  gate2317(.a(gate52inter5), .b(gate52inter2), .O(gate52inter6));
  inv1  gate2318(.a(G12), .O(gate52inter7));
  inv1  gate2319(.a(G281), .O(gate52inter8));
  nand2 gate2320(.a(gate52inter8), .b(gate52inter7), .O(gate52inter9));
  nand2 gate2321(.a(s_253), .b(gate52inter3), .O(gate52inter10));
  nor2  gate2322(.a(gate52inter10), .b(gate52inter9), .O(gate52inter11));
  nor2  gate2323(.a(gate52inter11), .b(gate52inter6), .O(gate52inter12));
  nand2 gate2324(.a(gate52inter12), .b(gate52inter1), .O(G373));

  xor2  gate1541(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate1542(.a(gate53inter0), .b(s_142), .O(gate53inter1));
  and2  gate1543(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate1544(.a(s_142), .O(gate53inter3));
  inv1  gate1545(.a(s_143), .O(gate53inter4));
  nand2 gate1546(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate1547(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate1548(.a(G13), .O(gate53inter7));
  inv1  gate1549(.a(G284), .O(gate53inter8));
  nand2 gate1550(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate1551(.a(s_143), .b(gate53inter3), .O(gate53inter10));
  nor2  gate1552(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate1553(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate1554(.a(gate53inter12), .b(gate53inter1), .O(G374));

  xor2  gate2465(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate2466(.a(gate54inter0), .b(s_274), .O(gate54inter1));
  and2  gate2467(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate2468(.a(s_274), .O(gate54inter3));
  inv1  gate2469(.a(s_275), .O(gate54inter4));
  nand2 gate2470(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate2471(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate2472(.a(G14), .O(gate54inter7));
  inv1  gate2473(.a(G284), .O(gate54inter8));
  nand2 gate2474(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate2475(.a(s_275), .b(gate54inter3), .O(gate54inter10));
  nor2  gate2476(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate2477(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate2478(.a(gate54inter12), .b(gate54inter1), .O(G375));

  xor2  gate1863(.a(G287), .b(G15), .O(gate55inter0));
  nand2 gate1864(.a(gate55inter0), .b(s_188), .O(gate55inter1));
  and2  gate1865(.a(G287), .b(G15), .O(gate55inter2));
  inv1  gate1866(.a(s_188), .O(gate55inter3));
  inv1  gate1867(.a(s_189), .O(gate55inter4));
  nand2 gate1868(.a(gate55inter4), .b(gate55inter3), .O(gate55inter5));
  nor2  gate1869(.a(gate55inter5), .b(gate55inter2), .O(gate55inter6));
  inv1  gate1870(.a(G15), .O(gate55inter7));
  inv1  gate1871(.a(G287), .O(gate55inter8));
  nand2 gate1872(.a(gate55inter8), .b(gate55inter7), .O(gate55inter9));
  nand2 gate1873(.a(s_189), .b(gate55inter3), .O(gate55inter10));
  nor2  gate1874(.a(gate55inter10), .b(gate55inter9), .O(gate55inter11));
  nor2  gate1875(.a(gate55inter11), .b(gate55inter6), .O(gate55inter12));
  nand2 gate1876(.a(gate55inter12), .b(gate55inter1), .O(G376));

  xor2  gate2773(.a(G287), .b(G16), .O(gate56inter0));
  nand2 gate2774(.a(gate56inter0), .b(s_318), .O(gate56inter1));
  and2  gate2775(.a(G287), .b(G16), .O(gate56inter2));
  inv1  gate2776(.a(s_318), .O(gate56inter3));
  inv1  gate2777(.a(s_319), .O(gate56inter4));
  nand2 gate2778(.a(gate56inter4), .b(gate56inter3), .O(gate56inter5));
  nor2  gate2779(.a(gate56inter5), .b(gate56inter2), .O(gate56inter6));
  inv1  gate2780(.a(G16), .O(gate56inter7));
  inv1  gate2781(.a(G287), .O(gate56inter8));
  nand2 gate2782(.a(gate56inter8), .b(gate56inter7), .O(gate56inter9));
  nand2 gate2783(.a(s_319), .b(gate56inter3), .O(gate56inter10));
  nor2  gate2784(.a(gate56inter10), .b(gate56inter9), .O(gate56inter11));
  nor2  gate2785(.a(gate56inter11), .b(gate56inter6), .O(gate56inter12));
  nand2 gate2786(.a(gate56inter12), .b(gate56inter1), .O(G377));
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );

  xor2  gate2969(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate2970(.a(gate59inter0), .b(s_346), .O(gate59inter1));
  and2  gate2971(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate2972(.a(s_346), .O(gate59inter3));
  inv1  gate2973(.a(s_347), .O(gate59inter4));
  nand2 gate2974(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate2975(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate2976(.a(G19), .O(gate59inter7));
  inv1  gate2977(.a(G293), .O(gate59inter8));
  nand2 gate2978(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate2979(.a(s_347), .b(gate59inter3), .O(gate59inter10));
  nor2  gate2980(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate2981(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate2982(.a(gate59inter12), .b(gate59inter1), .O(G380));

  xor2  gate2451(.a(G293), .b(G20), .O(gate60inter0));
  nand2 gate2452(.a(gate60inter0), .b(s_272), .O(gate60inter1));
  and2  gate2453(.a(G293), .b(G20), .O(gate60inter2));
  inv1  gate2454(.a(s_272), .O(gate60inter3));
  inv1  gate2455(.a(s_273), .O(gate60inter4));
  nand2 gate2456(.a(gate60inter4), .b(gate60inter3), .O(gate60inter5));
  nor2  gate2457(.a(gate60inter5), .b(gate60inter2), .O(gate60inter6));
  inv1  gate2458(.a(G20), .O(gate60inter7));
  inv1  gate2459(.a(G293), .O(gate60inter8));
  nand2 gate2460(.a(gate60inter8), .b(gate60inter7), .O(gate60inter9));
  nand2 gate2461(.a(s_273), .b(gate60inter3), .O(gate60inter10));
  nor2  gate2462(.a(gate60inter10), .b(gate60inter9), .O(gate60inter11));
  nor2  gate2463(.a(gate60inter11), .b(gate60inter6), .O(gate60inter12));
  nand2 gate2464(.a(gate60inter12), .b(gate60inter1), .O(G381));

  xor2  gate1877(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate1878(.a(gate61inter0), .b(s_190), .O(gate61inter1));
  and2  gate1879(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate1880(.a(s_190), .O(gate61inter3));
  inv1  gate1881(.a(s_191), .O(gate61inter4));
  nand2 gate1882(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate1883(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate1884(.a(G21), .O(gate61inter7));
  inv1  gate1885(.a(G296), .O(gate61inter8));
  nand2 gate1886(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate1887(.a(s_191), .b(gate61inter3), .O(gate61inter10));
  nor2  gate1888(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate1889(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate1890(.a(gate61inter12), .b(gate61inter1), .O(G382));
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate2199(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate2200(.a(gate63inter0), .b(s_236), .O(gate63inter1));
  and2  gate2201(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate2202(.a(s_236), .O(gate63inter3));
  inv1  gate2203(.a(s_237), .O(gate63inter4));
  nand2 gate2204(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate2205(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate2206(.a(G23), .O(gate63inter7));
  inv1  gate2207(.a(G299), .O(gate63inter8));
  nand2 gate2208(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate2209(.a(s_237), .b(gate63inter3), .O(gate63inter10));
  nor2  gate2210(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate2211(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate2212(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );

  xor2  gate2661(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate2662(.a(gate68inter0), .b(s_302), .O(gate68inter1));
  and2  gate2663(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate2664(.a(s_302), .O(gate68inter3));
  inv1  gate2665(.a(s_303), .O(gate68inter4));
  nand2 gate2666(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate2667(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate2668(.a(G28), .O(gate68inter7));
  inv1  gate2669(.a(G305), .O(gate68inter8));
  nand2 gate2670(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate2671(.a(s_303), .b(gate68inter3), .O(gate68inter10));
  nor2  gate2672(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate2673(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate2674(.a(gate68inter12), .b(gate68inter1), .O(G389));

  xor2  gate645(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate646(.a(gate69inter0), .b(s_14), .O(gate69inter1));
  and2  gate647(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate648(.a(s_14), .O(gate69inter3));
  inv1  gate649(.a(s_15), .O(gate69inter4));
  nand2 gate650(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate651(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate652(.a(G29), .O(gate69inter7));
  inv1  gate653(.a(G308), .O(gate69inter8));
  nand2 gate654(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate655(.a(s_15), .b(gate69inter3), .O(gate69inter10));
  nor2  gate656(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate657(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate658(.a(gate69inter12), .b(gate69inter1), .O(G390));

  xor2  gate2031(.a(G308), .b(G30), .O(gate70inter0));
  nand2 gate2032(.a(gate70inter0), .b(s_212), .O(gate70inter1));
  and2  gate2033(.a(G308), .b(G30), .O(gate70inter2));
  inv1  gate2034(.a(s_212), .O(gate70inter3));
  inv1  gate2035(.a(s_213), .O(gate70inter4));
  nand2 gate2036(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate2037(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate2038(.a(G30), .O(gate70inter7));
  inv1  gate2039(.a(G308), .O(gate70inter8));
  nand2 gate2040(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate2041(.a(s_213), .b(gate70inter3), .O(gate70inter10));
  nor2  gate2042(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate2043(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate2044(.a(gate70inter12), .b(gate70inter1), .O(G391));
nand2 gate71( .a(G31), .b(G311), .O(G392) );

  xor2  gate2171(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate2172(.a(gate72inter0), .b(s_232), .O(gate72inter1));
  and2  gate2173(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate2174(.a(s_232), .O(gate72inter3));
  inv1  gate2175(.a(s_233), .O(gate72inter4));
  nand2 gate2176(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate2177(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate2178(.a(G32), .O(gate72inter7));
  inv1  gate2179(.a(G311), .O(gate72inter8));
  nand2 gate2180(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate2181(.a(s_233), .b(gate72inter3), .O(gate72inter10));
  nor2  gate2182(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate2183(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate2184(.a(gate72inter12), .b(gate72inter1), .O(G393));
nand2 gate73( .a(G1), .b(G314), .O(G394) );

  xor2  gate561(.a(G314), .b(G5), .O(gate74inter0));
  nand2 gate562(.a(gate74inter0), .b(s_2), .O(gate74inter1));
  and2  gate563(.a(G314), .b(G5), .O(gate74inter2));
  inv1  gate564(.a(s_2), .O(gate74inter3));
  inv1  gate565(.a(s_3), .O(gate74inter4));
  nand2 gate566(.a(gate74inter4), .b(gate74inter3), .O(gate74inter5));
  nor2  gate567(.a(gate74inter5), .b(gate74inter2), .O(gate74inter6));
  inv1  gate568(.a(G5), .O(gate74inter7));
  inv1  gate569(.a(G314), .O(gate74inter8));
  nand2 gate570(.a(gate74inter8), .b(gate74inter7), .O(gate74inter9));
  nand2 gate571(.a(s_3), .b(gate74inter3), .O(gate74inter10));
  nor2  gate572(.a(gate74inter10), .b(gate74inter9), .O(gate74inter11));
  nor2  gate573(.a(gate74inter11), .b(gate74inter6), .O(gate74inter12));
  nand2 gate574(.a(gate74inter12), .b(gate74inter1), .O(G395));

  xor2  gate1401(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate1402(.a(gate75inter0), .b(s_122), .O(gate75inter1));
  and2  gate1403(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate1404(.a(s_122), .O(gate75inter3));
  inv1  gate1405(.a(s_123), .O(gate75inter4));
  nand2 gate1406(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate1407(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate1408(.a(G9), .O(gate75inter7));
  inv1  gate1409(.a(G317), .O(gate75inter8));
  nand2 gate1410(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate1411(.a(s_123), .b(gate75inter3), .O(gate75inter10));
  nor2  gate1412(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate1413(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate1414(.a(gate75inter12), .b(gate75inter1), .O(G396));

  xor2  gate2143(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate2144(.a(gate76inter0), .b(s_228), .O(gate76inter1));
  and2  gate2145(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate2146(.a(s_228), .O(gate76inter3));
  inv1  gate2147(.a(s_229), .O(gate76inter4));
  nand2 gate2148(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate2149(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate2150(.a(G13), .O(gate76inter7));
  inv1  gate2151(.a(G317), .O(gate76inter8));
  nand2 gate2152(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate2153(.a(s_229), .b(gate76inter3), .O(gate76inter10));
  nor2  gate2154(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate2155(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate2156(.a(gate76inter12), .b(gate76inter1), .O(G397));

  xor2  gate589(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate590(.a(gate77inter0), .b(s_6), .O(gate77inter1));
  and2  gate591(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate592(.a(s_6), .O(gate77inter3));
  inv1  gate593(.a(s_7), .O(gate77inter4));
  nand2 gate594(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate595(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate596(.a(G2), .O(gate77inter7));
  inv1  gate597(.a(G320), .O(gate77inter8));
  nand2 gate598(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate599(.a(s_7), .b(gate77inter3), .O(gate77inter10));
  nor2  gate600(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate601(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate602(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate883(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate884(.a(gate80inter0), .b(s_48), .O(gate80inter1));
  and2  gate885(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate886(.a(s_48), .O(gate80inter3));
  inv1  gate887(.a(s_49), .O(gate80inter4));
  nand2 gate888(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate889(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate890(.a(G14), .O(gate80inter7));
  inv1  gate891(.a(G323), .O(gate80inter8));
  nand2 gate892(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate893(.a(s_49), .b(gate80inter3), .O(gate80inter10));
  nor2  gate894(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate895(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate896(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );

  xor2  gate771(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate772(.a(gate83inter0), .b(s_32), .O(gate83inter1));
  and2  gate773(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate774(.a(s_32), .O(gate83inter3));
  inv1  gate775(.a(s_33), .O(gate83inter4));
  nand2 gate776(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate777(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate778(.a(G11), .O(gate83inter7));
  inv1  gate779(.a(G329), .O(gate83inter8));
  nand2 gate780(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate781(.a(s_33), .b(gate83inter3), .O(gate83inter10));
  nor2  gate782(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate783(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate784(.a(gate83inter12), .b(gate83inter1), .O(G404));

  xor2  gate2185(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate2186(.a(gate84inter0), .b(s_234), .O(gate84inter1));
  and2  gate2187(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate2188(.a(s_234), .O(gate84inter3));
  inv1  gate2189(.a(s_235), .O(gate84inter4));
  nand2 gate2190(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate2191(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate2192(.a(G15), .O(gate84inter7));
  inv1  gate2193(.a(G329), .O(gate84inter8));
  nand2 gate2194(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate2195(.a(s_235), .b(gate84inter3), .O(gate84inter10));
  nor2  gate2196(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate2197(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate2198(.a(gate84inter12), .b(gate84inter1), .O(G405));

  xor2  gate2633(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate2634(.a(gate85inter0), .b(s_298), .O(gate85inter1));
  and2  gate2635(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate2636(.a(s_298), .O(gate85inter3));
  inv1  gate2637(.a(s_299), .O(gate85inter4));
  nand2 gate2638(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate2639(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate2640(.a(G4), .O(gate85inter7));
  inv1  gate2641(.a(G332), .O(gate85inter8));
  nand2 gate2642(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate2643(.a(s_299), .b(gate85inter3), .O(gate85inter10));
  nor2  gate2644(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate2645(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate2646(.a(gate85inter12), .b(gate85inter1), .O(G406));

  xor2  gate1247(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate1248(.a(gate86inter0), .b(s_100), .O(gate86inter1));
  and2  gate1249(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate1250(.a(s_100), .O(gate86inter3));
  inv1  gate1251(.a(s_101), .O(gate86inter4));
  nand2 gate1252(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate1253(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate1254(.a(G8), .O(gate86inter7));
  inv1  gate1255(.a(G332), .O(gate86inter8));
  nand2 gate1256(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate1257(.a(s_101), .b(gate86inter3), .O(gate86inter10));
  nor2  gate1258(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate1259(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate1260(.a(gate86inter12), .b(gate86inter1), .O(G407));
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate2563(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate2564(.a(gate88inter0), .b(s_288), .O(gate88inter1));
  and2  gate2565(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate2566(.a(s_288), .O(gate88inter3));
  inv1  gate2567(.a(s_289), .O(gate88inter4));
  nand2 gate2568(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate2569(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate2570(.a(G16), .O(gate88inter7));
  inv1  gate2571(.a(G335), .O(gate88inter8));
  nand2 gate2572(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate2573(.a(s_289), .b(gate88inter3), .O(gate88inter10));
  nor2  gate2574(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate2575(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate2576(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );

  xor2  gate2269(.a(G338), .b(G21), .O(gate90inter0));
  nand2 gate2270(.a(gate90inter0), .b(s_246), .O(gate90inter1));
  and2  gate2271(.a(G338), .b(G21), .O(gate90inter2));
  inv1  gate2272(.a(s_246), .O(gate90inter3));
  inv1  gate2273(.a(s_247), .O(gate90inter4));
  nand2 gate2274(.a(gate90inter4), .b(gate90inter3), .O(gate90inter5));
  nor2  gate2275(.a(gate90inter5), .b(gate90inter2), .O(gate90inter6));
  inv1  gate2276(.a(G21), .O(gate90inter7));
  inv1  gate2277(.a(G338), .O(gate90inter8));
  nand2 gate2278(.a(gate90inter8), .b(gate90inter7), .O(gate90inter9));
  nand2 gate2279(.a(s_247), .b(gate90inter3), .O(gate90inter10));
  nor2  gate2280(.a(gate90inter10), .b(gate90inter9), .O(gate90inter11));
  nor2  gate2281(.a(gate90inter11), .b(gate90inter6), .O(gate90inter12));
  nand2 gate2282(.a(gate90inter12), .b(gate90inter1), .O(G411));
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );

  xor2  gate2101(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate2102(.a(gate95inter0), .b(s_222), .O(gate95inter1));
  and2  gate2103(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate2104(.a(s_222), .O(gate95inter3));
  inv1  gate2105(.a(s_223), .O(gate95inter4));
  nand2 gate2106(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate2107(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate2108(.a(G26), .O(gate95inter7));
  inv1  gate2109(.a(G347), .O(gate95inter8));
  nand2 gate2110(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate2111(.a(s_223), .b(gate95inter3), .O(gate95inter10));
  nor2  gate2112(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate2113(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate2114(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate1513(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate1514(.a(gate99inter0), .b(s_138), .O(gate99inter1));
  and2  gate1515(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate1516(.a(s_138), .O(gate99inter3));
  inv1  gate1517(.a(s_139), .O(gate99inter4));
  nand2 gate1518(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate1519(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate1520(.a(G27), .O(gate99inter7));
  inv1  gate1521(.a(G353), .O(gate99inter8));
  nand2 gate1522(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate1523(.a(s_139), .b(gate99inter3), .O(gate99inter10));
  nor2  gate1524(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate1525(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate1526(.a(gate99inter12), .b(gate99inter1), .O(G420));

  xor2  gate1345(.a(G353), .b(G31), .O(gate100inter0));
  nand2 gate1346(.a(gate100inter0), .b(s_114), .O(gate100inter1));
  and2  gate1347(.a(G353), .b(G31), .O(gate100inter2));
  inv1  gate1348(.a(s_114), .O(gate100inter3));
  inv1  gate1349(.a(s_115), .O(gate100inter4));
  nand2 gate1350(.a(gate100inter4), .b(gate100inter3), .O(gate100inter5));
  nor2  gate1351(.a(gate100inter5), .b(gate100inter2), .O(gate100inter6));
  inv1  gate1352(.a(G31), .O(gate100inter7));
  inv1  gate1353(.a(G353), .O(gate100inter8));
  nand2 gate1354(.a(gate100inter8), .b(gate100inter7), .O(gate100inter9));
  nand2 gate1355(.a(s_115), .b(gate100inter3), .O(gate100inter10));
  nor2  gate1356(.a(gate100inter10), .b(gate100inter9), .O(gate100inter11));
  nor2  gate1357(.a(gate100inter11), .b(gate100inter6), .O(gate100inter12));
  nand2 gate1358(.a(gate100inter12), .b(gate100inter1), .O(G421));
nand2 gate101( .a(G20), .b(G356), .O(G422) );

  xor2  gate1597(.a(G356), .b(G24), .O(gate102inter0));
  nand2 gate1598(.a(gate102inter0), .b(s_150), .O(gate102inter1));
  and2  gate1599(.a(G356), .b(G24), .O(gate102inter2));
  inv1  gate1600(.a(s_150), .O(gate102inter3));
  inv1  gate1601(.a(s_151), .O(gate102inter4));
  nand2 gate1602(.a(gate102inter4), .b(gate102inter3), .O(gate102inter5));
  nor2  gate1603(.a(gate102inter5), .b(gate102inter2), .O(gate102inter6));
  inv1  gate1604(.a(G24), .O(gate102inter7));
  inv1  gate1605(.a(G356), .O(gate102inter8));
  nand2 gate1606(.a(gate102inter8), .b(gate102inter7), .O(gate102inter9));
  nand2 gate1607(.a(s_151), .b(gate102inter3), .O(gate102inter10));
  nor2  gate1608(.a(gate102inter10), .b(gate102inter9), .O(gate102inter11));
  nor2  gate1609(.a(gate102inter11), .b(gate102inter6), .O(gate102inter12));
  nand2 gate1610(.a(gate102inter12), .b(gate102inter1), .O(G423));
nand2 gate103( .a(G28), .b(G359), .O(G424) );

  xor2  gate2535(.a(G359), .b(G32), .O(gate104inter0));
  nand2 gate2536(.a(gate104inter0), .b(s_284), .O(gate104inter1));
  and2  gate2537(.a(G359), .b(G32), .O(gate104inter2));
  inv1  gate2538(.a(s_284), .O(gate104inter3));
  inv1  gate2539(.a(s_285), .O(gate104inter4));
  nand2 gate2540(.a(gate104inter4), .b(gate104inter3), .O(gate104inter5));
  nor2  gate2541(.a(gate104inter5), .b(gate104inter2), .O(gate104inter6));
  inv1  gate2542(.a(G32), .O(gate104inter7));
  inv1  gate2543(.a(G359), .O(gate104inter8));
  nand2 gate2544(.a(gate104inter8), .b(gate104inter7), .O(gate104inter9));
  nand2 gate2545(.a(s_285), .b(gate104inter3), .O(gate104inter10));
  nor2  gate2546(.a(gate104inter10), .b(gate104inter9), .O(gate104inter11));
  nor2  gate2547(.a(gate104inter11), .b(gate104inter6), .O(gate104inter12));
  nand2 gate2548(.a(gate104inter12), .b(gate104inter1), .O(G425));

  xor2  gate2801(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate2802(.a(gate105inter0), .b(s_322), .O(gate105inter1));
  and2  gate2803(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate2804(.a(s_322), .O(gate105inter3));
  inv1  gate2805(.a(s_323), .O(gate105inter4));
  nand2 gate2806(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate2807(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate2808(.a(G362), .O(gate105inter7));
  inv1  gate2809(.a(G363), .O(gate105inter8));
  nand2 gate2810(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate2811(.a(s_323), .b(gate105inter3), .O(gate105inter10));
  nor2  gate2812(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate2813(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate2814(.a(gate105inter12), .b(gate105inter1), .O(G426));
nand2 gate106( .a(G364), .b(G365), .O(G429) );

  xor2  gate1821(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate1822(.a(gate107inter0), .b(s_182), .O(gate107inter1));
  and2  gate1823(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate1824(.a(s_182), .O(gate107inter3));
  inv1  gate1825(.a(s_183), .O(gate107inter4));
  nand2 gate1826(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate1827(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate1828(.a(G366), .O(gate107inter7));
  inv1  gate1829(.a(G367), .O(gate107inter8));
  nand2 gate1830(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate1831(.a(s_183), .b(gate107inter3), .O(gate107inter10));
  nor2  gate1832(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate1833(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate1834(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );

  xor2  gate2703(.a(G381), .b(G380), .O(gate114inter0));
  nand2 gate2704(.a(gate114inter0), .b(s_308), .O(gate114inter1));
  and2  gate2705(.a(G381), .b(G380), .O(gate114inter2));
  inv1  gate2706(.a(s_308), .O(gate114inter3));
  inv1  gate2707(.a(s_309), .O(gate114inter4));
  nand2 gate2708(.a(gate114inter4), .b(gate114inter3), .O(gate114inter5));
  nor2  gate2709(.a(gate114inter5), .b(gate114inter2), .O(gate114inter6));
  inv1  gate2710(.a(G380), .O(gate114inter7));
  inv1  gate2711(.a(G381), .O(gate114inter8));
  nand2 gate2712(.a(gate114inter8), .b(gate114inter7), .O(gate114inter9));
  nand2 gate2713(.a(s_309), .b(gate114inter3), .O(gate114inter10));
  nor2  gate2714(.a(gate114inter10), .b(gate114inter9), .O(gate114inter11));
  nor2  gate2715(.a(gate114inter11), .b(gate114inter6), .O(gate114inter12));
  nand2 gate2716(.a(gate114inter12), .b(gate114inter1), .O(G453));

  xor2  gate1051(.a(G383), .b(G382), .O(gate115inter0));
  nand2 gate1052(.a(gate115inter0), .b(s_72), .O(gate115inter1));
  and2  gate1053(.a(G383), .b(G382), .O(gate115inter2));
  inv1  gate1054(.a(s_72), .O(gate115inter3));
  inv1  gate1055(.a(s_73), .O(gate115inter4));
  nand2 gate1056(.a(gate115inter4), .b(gate115inter3), .O(gate115inter5));
  nor2  gate1057(.a(gate115inter5), .b(gate115inter2), .O(gate115inter6));
  inv1  gate1058(.a(G382), .O(gate115inter7));
  inv1  gate1059(.a(G383), .O(gate115inter8));
  nand2 gate1060(.a(gate115inter8), .b(gate115inter7), .O(gate115inter9));
  nand2 gate1061(.a(s_73), .b(gate115inter3), .O(gate115inter10));
  nor2  gate1062(.a(gate115inter10), .b(gate115inter9), .O(gate115inter11));
  nor2  gate1063(.a(gate115inter11), .b(gate115inter6), .O(gate115inter12));
  nand2 gate1064(.a(gate115inter12), .b(gate115inter1), .O(G456));

  xor2  gate2577(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate2578(.a(gate116inter0), .b(s_290), .O(gate116inter1));
  and2  gate2579(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate2580(.a(s_290), .O(gate116inter3));
  inv1  gate2581(.a(s_291), .O(gate116inter4));
  nand2 gate2582(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate2583(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate2584(.a(G384), .O(gate116inter7));
  inv1  gate2585(.a(G385), .O(gate116inter8));
  nand2 gate2586(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate2587(.a(s_291), .b(gate116inter3), .O(gate116inter10));
  nor2  gate2588(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate2589(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate2590(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );

  xor2  gate617(.a(G401), .b(G400), .O(gate124inter0));
  nand2 gate618(.a(gate124inter0), .b(s_10), .O(gate124inter1));
  and2  gate619(.a(G401), .b(G400), .O(gate124inter2));
  inv1  gate620(.a(s_10), .O(gate124inter3));
  inv1  gate621(.a(s_11), .O(gate124inter4));
  nand2 gate622(.a(gate124inter4), .b(gate124inter3), .O(gate124inter5));
  nor2  gate623(.a(gate124inter5), .b(gate124inter2), .O(gate124inter6));
  inv1  gate624(.a(G400), .O(gate124inter7));
  inv1  gate625(.a(G401), .O(gate124inter8));
  nand2 gate626(.a(gate124inter8), .b(gate124inter7), .O(gate124inter9));
  nand2 gate627(.a(s_11), .b(gate124inter3), .O(gate124inter10));
  nor2  gate628(.a(gate124inter10), .b(gate124inter9), .O(gate124inter11));
  nor2  gate629(.a(gate124inter11), .b(gate124inter6), .O(gate124inter12));
  nand2 gate630(.a(gate124inter12), .b(gate124inter1), .O(G483));

  xor2  gate1289(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate1290(.a(gate125inter0), .b(s_106), .O(gate125inter1));
  and2  gate1291(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate1292(.a(s_106), .O(gate125inter3));
  inv1  gate1293(.a(s_107), .O(gate125inter4));
  nand2 gate1294(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate1295(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate1296(.a(G402), .O(gate125inter7));
  inv1  gate1297(.a(G403), .O(gate125inter8));
  nand2 gate1298(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate1299(.a(s_107), .b(gate125inter3), .O(gate125inter10));
  nor2  gate1300(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate1301(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate1302(.a(gate125inter12), .b(gate125inter1), .O(G486));

  xor2  gate1429(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate1430(.a(gate126inter0), .b(s_126), .O(gate126inter1));
  and2  gate1431(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate1432(.a(s_126), .O(gate126inter3));
  inv1  gate1433(.a(s_127), .O(gate126inter4));
  nand2 gate1434(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate1435(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate1436(.a(G404), .O(gate126inter7));
  inv1  gate1437(.a(G405), .O(gate126inter8));
  nand2 gate1438(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate1439(.a(s_127), .b(gate126inter3), .O(gate126inter10));
  nor2  gate1440(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate1441(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate1442(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );

  xor2  gate3039(.a(G409), .b(G408), .O(gate128inter0));
  nand2 gate3040(.a(gate128inter0), .b(s_356), .O(gate128inter1));
  and2  gate3041(.a(G409), .b(G408), .O(gate128inter2));
  inv1  gate3042(.a(s_356), .O(gate128inter3));
  inv1  gate3043(.a(s_357), .O(gate128inter4));
  nand2 gate3044(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate3045(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate3046(.a(G408), .O(gate128inter7));
  inv1  gate3047(.a(G409), .O(gate128inter8));
  nand2 gate3048(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate3049(.a(s_357), .b(gate128inter3), .O(gate128inter10));
  nor2  gate3050(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate3051(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate3052(.a(gate128inter12), .b(gate128inter1), .O(G495));

  xor2  gate3025(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate3026(.a(gate129inter0), .b(s_354), .O(gate129inter1));
  and2  gate3027(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate3028(.a(s_354), .O(gate129inter3));
  inv1  gate3029(.a(s_355), .O(gate129inter4));
  nand2 gate3030(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate3031(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate3032(.a(G410), .O(gate129inter7));
  inv1  gate3033(.a(G411), .O(gate129inter8));
  nand2 gate3034(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate3035(.a(s_355), .b(gate129inter3), .O(gate129inter10));
  nor2  gate3036(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate3037(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate3038(.a(gate129inter12), .b(gate129inter1), .O(G498));

  xor2  gate1989(.a(G413), .b(G412), .O(gate130inter0));
  nand2 gate1990(.a(gate130inter0), .b(s_206), .O(gate130inter1));
  and2  gate1991(.a(G413), .b(G412), .O(gate130inter2));
  inv1  gate1992(.a(s_206), .O(gate130inter3));
  inv1  gate1993(.a(s_207), .O(gate130inter4));
  nand2 gate1994(.a(gate130inter4), .b(gate130inter3), .O(gate130inter5));
  nor2  gate1995(.a(gate130inter5), .b(gate130inter2), .O(gate130inter6));
  inv1  gate1996(.a(G412), .O(gate130inter7));
  inv1  gate1997(.a(G413), .O(gate130inter8));
  nand2 gate1998(.a(gate130inter8), .b(gate130inter7), .O(gate130inter9));
  nand2 gate1999(.a(s_207), .b(gate130inter3), .O(gate130inter10));
  nor2  gate2000(.a(gate130inter10), .b(gate130inter9), .O(gate130inter11));
  nor2  gate2001(.a(gate130inter11), .b(gate130inter6), .O(gate130inter12));
  nand2 gate2002(.a(gate130inter12), .b(gate130inter1), .O(G501));

  xor2  gate2619(.a(G415), .b(G414), .O(gate131inter0));
  nand2 gate2620(.a(gate131inter0), .b(s_296), .O(gate131inter1));
  and2  gate2621(.a(G415), .b(G414), .O(gate131inter2));
  inv1  gate2622(.a(s_296), .O(gate131inter3));
  inv1  gate2623(.a(s_297), .O(gate131inter4));
  nand2 gate2624(.a(gate131inter4), .b(gate131inter3), .O(gate131inter5));
  nor2  gate2625(.a(gate131inter5), .b(gate131inter2), .O(gate131inter6));
  inv1  gate2626(.a(G414), .O(gate131inter7));
  inv1  gate2627(.a(G415), .O(gate131inter8));
  nand2 gate2628(.a(gate131inter8), .b(gate131inter7), .O(gate131inter9));
  nand2 gate2629(.a(s_297), .b(gate131inter3), .O(gate131inter10));
  nor2  gate2630(.a(gate131inter10), .b(gate131inter9), .O(gate131inter11));
  nor2  gate2631(.a(gate131inter11), .b(gate131inter6), .O(gate131inter12));
  nand2 gate2632(.a(gate131inter12), .b(gate131inter1), .O(G504));
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate1835(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate1836(.a(gate136inter0), .b(s_184), .O(gate136inter1));
  and2  gate1837(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate1838(.a(s_184), .O(gate136inter3));
  inv1  gate1839(.a(s_185), .O(gate136inter4));
  nand2 gate1840(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate1841(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate1842(.a(G424), .O(gate136inter7));
  inv1  gate1843(.a(G425), .O(gate136inter8));
  nand2 gate1844(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate1845(.a(s_185), .b(gate136inter3), .O(gate136inter10));
  nor2  gate1846(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate1847(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate1848(.a(gate136inter12), .b(gate136inter1), .O(G519));

  xor2  gate1191(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate1192(.a(gate137inter0), .b(s_92), .O(gate137inter1));
  and2  gate1193(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate1194(.a(s_92), .O(gate137inter3));
  inv1  gate1195(.a(s_93), .O(gate137inter4));
  nand2 gate1196(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate1197(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate1198(.a(G426), .O(gate137inter7));
  inv1  gate1199(.a(G429), .O(gate137inter8));
  nand2 gate1200(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate1201(.a(s_93), .b(gate137inter3), .O(gate137inter10));
  nor2  gate1202(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate1203(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate1204(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );

  xor2  gate2367(.a(G441), .b(G438), .O(gate139inter0));
  nand2 gate2368(.a(gate139inter0), .b(s_260), .O(gate139inter1));
  and2  gate2369(.a(G441), .b(G438), .O(gate139inter2));
  inv1  gate2370(.a(s_260), .O(gate139inter3));
  inv1  gate2371(.a(s_261), .O(gate139inter4));
  nand2 gate2372(.a(gate139inter4), .b(gate139inter3), .O(gate139inter5));
  nor2  gate2373(.a(gate139inter5), .b(gate139inter2), .O(gate139inter6));
  inv1  gate2374(.a(G438), .O(gate139inter7));
  inv1  gate2375(.a(G441), .O(gate139inter8));
  nand2 gate2376(.a(gate139inter8), .b(gate139inter7), .O(gate139inter9));
  nand2 gate2377(.a(s_261), .b(gate139inter3), .O(gate139inter10));
  nor2  gate2378(.a(gate139inter10), .b(gate139inter9), .O(gate139inter11));
  nor2  gate2379(.a(gate139inter11), .b(gate139inter6), .O(gate139inter12));
  nand2 gate2380(.a(gate139inter12), .b(gate139inter1), .O(G528));

  xor2  gate1555(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate1556(.a(gate140inter0), .b(s_144), .O(gate140inter1));
  and2  gate1557(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate1558(.a(s_144), .O(gate140inter3));
  inv1  gate1559(.a(s_145), .O(gate140inter4));
  nand2 gate1560(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate1561(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate1562(.a(G444), .O(gate140inter7));
  inv1  gate1563(.a(G447), .O(gate140inter8));
  nand2 gate1564(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate1565(.a(s_145), .b(gate140inter3), .O(gate140inter10));
  nor2  gate1566(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate1567(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate1568(.a(gate140inter12), .b(gate140inter1), .O(G531));

  xor2  gate659(.a(G453), .b(G450), .O(gate141inter0));
  nand2 gate660(.a(gate141inter0), .b(s_16), .O(gate141inter1));
  and2  gate661(.a(G453), .b(G450), .O(gate141inter2));
  inv1  gate662(.a(s_16), .O(gate141inter3));
  inv1  gate663(.a(s_17), .O(gate141inter4));
  nand2 gate664(.a(gate141inter4), .b(gate141inter3), .O(gate141inter5));
  nor2  gate665(.a(gate141inter5), .b(gate141inter2), .O(gate141inter6));
  inv1  gate666(.a(G450), .O(gate141inter7));
  inv1  gate667(.a(G453), .O(gate141inter8));
  nand2 gate668(.a(gate141inter8), .b(gate141inter7), .O(gate141inter9));
  nand2 gate669(.a(s_17), .b(gate141inter3), .O(gate141inter10));
  nor2  gate670(.a(gate141inter10), .b(gate141inter9), .O(gate141inter11));
  nor2  gate671(.a(gate141inter11), .b(gate141inter6), .O(gate141inter12));
  nand2 gate672(.a(gate141inter12), .b(gate141inter1), .O(G534));

  xor2  gate981(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate982(.a(gate142inter0), .b(s_62), .O(gate142inter1));
  and2  gate983(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate984(.a(s_62), .O(gate142inter3));
  inv1  gate985(.a(s_63), .O(gate142inter4));
  nand2 gate986(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate987(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate988(.a(G456), .O(gate142inter7));
  inv1  gate989(.a(G459), .O(gate142inter8));
  nand2 gate990(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate991(.a(s_63), .b(gate142inter3), .O(gate142inter10));
  nor2  gate992(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate993(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate994(.a(gate142inter12), .b(gate142inter1), .O(G537));

  xor2  gate1737(.a(G465), .b(G462), .O(gate143inter0));
  nand2 gate1738(.a(gate143inter0), .b(s_170), .O(gate143inter1));
  and2  gate1739(.a(G465), .b(G462), .O(gate143inter2));
  inv1  gate1740(.a(s_170), .O(gate143inter3));
  inv1  gate1741(.a(s_171), .O(gate143inter4));
  nand2 gate1742(.a(gate143inter4), .b(gate143inter3), .O(gate143inter5));
  nor2  gate1743(.a(gate143inter5), .b(gate143inter2), .O(gate143inter6));
  inv1  gate1744(.a(G462), .O(gate143inter7));
  inv1  gate1745(.a(G465), .O(gate143inter8));
  nand2 gate1746(.a(gate143inter8), .b(gate143inter7), .O(gate143inter9));
  nand2 gate1747(.a(s_171), .b(gate143inter3), .O(gate143inter10));
  nor2  gate1748(.a(gate143inter10), .b(gate143inter9), .O(gate143inter11));
  nor2  gate1749(.a(gate143inter11), .b(gate143inter6), .O(gate143inter12));
  nand2 gate1750(.a(gate143inter12), .b(gate143inter1), .O(G540));
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );

  xor2  gate2283(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate2284(.a(gate146inter0), .b(s_248), .O(gate146inter1));
  and2  gate2285(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate2286(.a(s_248), .O(gate146inter3));
  inv1  gate2287(.a(s_249), .O(gate146inter4));
  nand2 gate2288(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate2289(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate2290(.a(G480), .O(gate146inter7));
  inv1  gate2291(.a(G483), .O(gate146inter8));
  nand2 gate2292(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate2293(.a(s_249), .b(gate146inter3), .O(gate146inter10));
  nor2  gate2294(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate2295(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate2296(.a(gate146inter12), .b(gate146inter1), .O(G549));
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate2129(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate2130(.a(gate148inter0), .b(s_226), .O(gate148inter1));
  and2  gate2131(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate2132(.a(s_226), .O(gate148inter3));
  inv1  gate2133(.a(s_227), .O(gate148inter4));
  nand2 gate2134(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate2135(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate2136(.a(G492), .O(gate148inter7));
  inv1  gate2137(.a(G495), .O(gate148inter8));
  nand2 gate2138(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate2139(.a(s_227), .b(gate148inter3), .O(gate148inter10));
  nor2  gate2140(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate2141(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate2142(.a(gate148inter12), .b(gate148inter1), .O(G555));

  xor2  gate1667(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate1668(.a(gate149inter0), .b(s_160), .O(gate149inter1));
  and2  gate1669(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate1670(.a(s_160), .O(gate149inter3));
  inv1  gate1671(.a(s_161), .O(gate149inter4));
  nand2 gate1672(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate1673(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate1674(.a(G498), .O(gate149inter7));
  inv1  gate1675(.a(G501), .O(gate149inter8));
  nand2 gate1676(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate1677(.a(s_161), .b(gate149inter3), .O(gate149inter10));
  nor2  gate1678(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate1679(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate1680(.a(gate149inter12), .b(gate149inter1), .O(G558));

  xor2  gate1233(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate1234(.a(gate150inter0), .b(s_98), .O(gate150inter1));
  and2  gate1235(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate1236(.a(s_98), .O(gate150inter3));
  inv1  gate1237(.a(s_99), .O(gate150inter4));
  nand2 gate1238(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate1239(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate1240(.a(G504), .O(gate150inter7));
  inv1  gate1241(.a(G507), .O(gate150inter8));
  nand2 gate1242(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate1243(.a(s_99), .b(gate150inter3), .O(gate150inter10));
  nor2  gate1244(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate1245(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate1246(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );

  xor2  gate3011(.a(G519), .b(G516), .O(gate152inter0));
  nand2 gate3012(.a(gate152inter0), .b(s_352), .O(gate152inter1));
  and2  gate3013(.a(G519), .b(G516), .O(gate152inter2));
  inv1  gate3014(.a(s_352), .O(gate152inter3));
  inv1  gate3015(.a(s_353), .O(gate152inter4));
  nand2 gate3016(.a(gate152inter4), .b(gate152inter3), .O(gate152inter5));
  nor2  gate3017(.a(gate152inter5), .b(gate152inter2), .O(gate152inter6));
  inv1  gate3018(.a(G516), .O(gate152inter7));
  inv1  gate3019(.a(G519), .O(gate152inter8));
  nand2 gate3020(.a(gate152inter8), .b(gate152inter7), .O(gate152inter9));
  nand2 gate3021(.a(s_353), .b(gate152inter3), .O(gate152inter10));
  nor2  gate3022(.a(gate152inter10), .b(gate152inter9), .O(gate152inter11));
  nor2  gate3023(.a(gate152inter11), .b(gate152inter6), .O(gate152inter12));
  nand2 gate3024(.a(gate152inter12), .b(gate152inter1), .O(G567));

  xor2  gate673(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate674(.a(gate153inter0), .b(s_18), .O(gate153inter1));
  and2  gate675(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate676(.a(s_18), .O(gate153inter3));
  inv1  gate677(.a(s_19), .O(gate153inter4));
  nand2 gate678(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate679(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate680(.a(G426), .O(gate153inter7));
  inv1  gate681(.a(G522), .O(gate153inter8));
  nand2 gate682(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate683(.a(s_19), .b(gate153inter3), .O(gate153inter10));
  nor2  gate684(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate685(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate686(.a(gate153inter12), .b(gate153inter1), .O(G570));

  xor2  gate799(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate800(.a(gate154inter0), .b(s_36), .O(gate154inter1));
  and2  gate801(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate802(.a(s_36), .O(gate154inter3));
  inv1  gate803(.a(s_37), .O(gate154inter4));
  nand2 gate804(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate805(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate806(.a(G429), .O(gate154inter7));
  inv1  gate807(.a(G522), .O(gate154inter8));
  nand2 gate808(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate809(.a(s_37), .b(gate154inter3), .O(gate154inter10));
  nor2  gate810(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate811(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate812(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );

  xor2  gate2913(.a(G528), .b(G438), .O(gate157inter0));
  nand2 gate2914(.a(gate157inter0), .b(s_338), .O(gate157inter1));
  and2  gate2915(.a(G528), .b(G438), .O(gate157inter2));
  inv1  gate2916(.a(s_338), .O(gate157inter3));
  inv1  gate2917(.a(s_339), .O(gate157inter4));
  nand2 gate2918(.a(gate157inter4), .b(gate157inter3), .O(gate157inter5));
  nor2  gate2919(.a(gate157inter5), .b(gate157inter2), .O(gate157inter6));
  inv1  gate2920(.a(G438), .O(gate157inter7));
  inv1  gate2921(.a(G528), .O(gate157inter8));
  nand2 gate2922(.a(gate157inter8), .b(gate157inter7), .O(gate157inter9));
  nand2 gate2923(.a(s_339), .b(gate157inter3), .O(gate157inter10));
  nor2  gate2924(.a(gate157inter10), .b(gate157inter9), .O(gate157inter11));
  nor2  gate2925(.a(gate157inter11), .b(gate157inter6), .O(gate157inter12));
  nand2 gate2926(.a(gate157inter12), .b(gate157inter1), .O(G574));

  xor2  gate2857(.a(G528), .b(G441), .O(gate158inter0));
  nand2 gate2858(.a(gate158inter0), .b(s_330), .O(gate158inter1));
  and2  gate2859(.a(G528), .b(G441), .O(gate158inter2));
  inv1  gate2860(.a(s_330), .O(gate158inter3));
  inv1  gate2861(.a(s_331), .O(gate158inter4));
  nand2 gate2862(.a(gate158inter4), .b(gate158inter3), .O(gate158inter5));
  nor2  gate2863(.a(gate158inter5), .b(gate158inter2), .O(gate158inter6));
  inv1  gate2864(.a(G441), .O(gate158inter7));
  inv1  gate2865(.a(G528), .O(gate158inter8));
  nand2 gate2866(.a(gate158inter8), .b(gate158inter7), .O(gate158inter9));
  nand2 gate2867(.a(s_331), .b(gate158inter3), .O(gate158inter10));
  nor2  gate2868(.a(gate158inter10), .b(gate158inter9), .O(gate158inter11));
  nor2  gate2869(.a(gate158inter11), .b(gate158inter6), .O(gate158inter12));
  nand2 gate2870(.a(gate158inter12), .b(gate158inter1), .O(G575));

  xor2  gate2227(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate2228(.a(gate159inter0), .b(s_240), .O(gate159inter1));
  and2  gate2229(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate2230(.a(s_240), .O(gate159inter3));
  inv1  gate2231(.a(s_241), .O(gate159inter4));
  nand2 gate2232(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate2233(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate2234(.a(G444), .O(gate159inter7));
  inv1  gate2235(.a(G531), .O(gate159inter8));
  nand2 gate2236(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate2237(.a(s_241), .b(gate159inter3), .O(gate159inter10));
  nor2  gate2238(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate2239(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate2240(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate1695(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate1696(.a(gate162inter0), .b(s_164), .O(gate162inter1));
  and2  gate1697(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate1698(.a(s_164), .O(gate162inter3));
  inv1  gate1699(.a(s_165), .O(gate162inter4));
  nand2 gate1700(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate1701(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate1702(.a(G453), .O(gate162inter7));
  inv1  gate1703(.a(G534), .O(gate162inter8));
  nand2 gate1704(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate1705(.a(s_165), .b(gate162inter3), .O(gate162inter10));
  nor2  gate1706(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate1707(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate1708(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate1373(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate1374(.a(gate165inter0), .b(s_118), .O(gate165inter1));
  and2  gate1375(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate1376(.a(s_118), .O(gate165inter3));
  inv1  gate1377(.a(s_119), .O(gate165inter4));
  nand2 gate1378(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate1379(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate1380(.a(G462), .O(gate165inter7));
  inv1  gate1381(.a(G540), .O(gate165inter8));
  nand2 gate1382(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate1383(.a(s_119), .b(gate165inter3), .O(gate165inter10));
  nor2  gate1384(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate1385(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate1386(.a(gate165inter12), .b(gate165inter1), .O(G582));
nand2 gate166( .a(G465), .b(G540), .O(G583) );

  xor2  gate1303(.a(G543), .b(G468), .O(gate167inter0));
  nand2 gate1304(.a(gate167inter0), .b(s_108), .O(gate167inter1));
  and2  gate1305(.a(G543), .b(G468), .O(gate167inter2));
  inv1  gate1306(.a(s_108), .O(gate167inter3));
  inv1  gate1307(.a(s_109), .O(gate167inter4));
  nand2 gate1308(.a(gate167inter4), .b(gate167inter3), .O(gate167inter5));
  nor2  gate1309(.a(gate167inter5), .b(gate167inter2), .O(gate167inter6));
  inv1  gate1310(.a(G468), .O(gate167inter7));
  inv1  gate1311(.a(G543), .O(gate167inter8));
  nand2 gate1312(.a(gate167inter8), .b(gate167inter7), .O(gate167inter9));
  nand2 gate1313(.a(s_109), .b(gate167inter3), .O(gate167inter10));
  nor2  gate1314(.a(gate167inter10), .b(gate167inter9), .O(gate167inter11));
  nor2  gate1315(.a(gate167inter11), .b(gate167inter6), .O(gate167inter12));
  nand2 gate1316(.a(gate167inter12), .b(gate167inter1), .O(G584));
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );

  xor2  gate2941(.a(G546), .b(G477), .O(gate170inter0));
  nand2 gate2942(.a(gate170inter0), .b(s_342), .O(gate170inter1));
  and2  gate2943(.a(G546), .b(G477), .O(gate170inter2));
  inv1  gate2944(.a(s_342), .O(gate170inter3));
  inv1  gate2945(.a(s_343), .O(gate170inter4));
  nand2 gate2946(.a(gate170inter4), .b(gate170inter3), .O(gate170inter5));
  nor2  gate2947(.a(gate170inter5), .b(gate170inter2), .O(gate170inter6));
  inv1  gate2948(.a(G477), .O(gate170inter7));
  inv1  gate2949(.a(G546), .O(gate170inter8));
  nand2 gate2950(.a(gate170inter8), .b(gate170inter7), .O(gate170inter9));
  nand2 gate2951(.a(s_343), .b(gate170inter3), .O(gate170inter10));
  nor2  gate2952(.a(gate170inter10), .b(gate170inter9), .O(gate170inter11));
  nor2  gate2953(.a(gate170inter11), .b(gate170inter6), .O(gate170inter12));
  nand2 gate2954(.a(gate170inter12), .b(gate170inter1), .O(G587));
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate2759(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate2760(.a(gate173inter0), .b(s_316), .O(gate173inter1));
  and2  gate2761(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate2762(.a(s_316), .O(gate173inter3));
  inv1  gate2763(.a(s_317), .O(gate173inter4));
  nand2 gate2764(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate2765(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate2766(.a(G486), .O(gate173inter7));
  inv1  gate2767(.a(G552), .O(gate173inter8));
  nand2 gate2768(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate2769(.a(s_317), .b(gate173inter3), .O(gate173inter10));
  nor2  gate2770(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate2771(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate2772(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate1639(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate1640(.a(gate178inter0), .b(s_156), .O(gate178inter1));
  and2  gate1641(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate1642(.a(s_156), .O(gate178inter3));
  inv1  gate1643(.a(s_157), .O(gate178inter4));
  nand2 gate1644(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate1645(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate1646(.a(G501), .O(gate178inter7));
  inv1  gate1647(.a(G558), .O(gate178inter8));
  nand2 gate1648(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate1649(.a(s_157), .b(gate178inter3), .O(gate178inter10));
  nor2  gate1650(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate1651(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate1652(.a(gate178inter12), .b(gate178inter1), .O(G595));

  xor2  gate2997(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate2998(.a(gate179inter0), .b(s_350), .O(gate179inter1));
  and2  gate2999(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate3000(.a(s_350), .O(gate179inter3));
  inv1  gate3001(.a(s_351), .O(gate179inter4));
  nand2 gate3002(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate3003(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate3004(.a(G504), .O(gate179inter7));
  inv1  gate3005(.a(G561), .O(gate179inter8));
  nand2 gate3006(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate3007(.a(s_351), .b(gate179inter3), .O(gate179inter10));
  nor2  gate3008(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate3009(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate3010(.a(gate179inter12), .b(gate179inter1), .O(G596));
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );

  xor2  gate827(.a(G564), .b(G513), .O(gate182inter0));
  nand2 gate828(.a(gate182inter0), .b(s_40), .O(gate182inter1));
  and2  gate829(.a(G564), .b(G513), .O(gate182inter2));
  inv1  gate830(.a(s_40), .O(gate182inter3));
  inv1  gate831(.a(s_41), .O(gate182inter4));
  nand2 gate832(.a(gate182inter4), .b(gate182inter3), .O(gate182inter5));
  nor2  gate833(.a(gate182inter5), .b(gate182inter2), .O(gate182inter6));
  inv1  gate834(.a(G513), .O(gate182inter7));
  inv1  gate835(.a(G564), .O(gate182inter8));
  nand2 gate836(.a(gate182inter8), .b(gate182inter7), .O(gate182inter9));
  nand2 gate837(.a(s_41), .b(gate182inter3), .O(gate182inter10));
  nor2  gate838(.a(gate182inter10), .b(gate182inter9), .O(gate182inter11));
  nor2  gate839(.a(gate182inter11), .b(gate182inter6), .O(gate182inter12));
  nand2 gate840(.a(gate182inter12), .b(gate182inter1), .O(G599));
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );

  xor2  gate2087(.a(G571), .b(G570), .O(gate185inter0));
  nand2 gate2088(.a(gate185inter0), .b(s_220), .O(gate185inter1));
  and2  gate2089(.a(G571), .b(G570), .O(gate185inter2));
  inv1  gate2090(.a(s_220), .O(gate185inter3));
  inv1  gate2091(.a(s_221), .O(gate185inter4));
  nand2 gate2092(.a(gate185inter4), .b(gate185inter3), .O(gate185inter5));
  nor2  gate2093(.a(gate185inter5), .b(gate185inter2), .O(gate185inter6));
  inv1  gate2094(.a(G570), .O(gate185inter7));
  inv1  gate2095(.a(G571), .O(gate185inter8));
  nand2 gate2096(.a(gate185inter8), .b(gate185inter7), .O(gate185inter9));
  nand2 gate2097(.a(s_221), .b(gate185inter3), .O(gate185inter10));
  nor2  gate2098(.a(gate185inter10), .b(gate185inter9), .O(gate185inter11));
  nor2  gate2099(.a(gate185inter11), .b(gate185inter6), .O(gate185inter12));
  nand2 gate2100(.a(gate185inter12), .b(gate185inter1), .O(G602));
nand2 gate186( .a(G572), .b(G573), .O(G607) );

  xor2  gate1219(.a(G575), .b(G574), .O(gate187inter0));
  nand2 gate1220(.a(gate187inter0), .b(s_96), .O(gate187inter1));
  and2  gate1221(.a(G575), .b(G574), .O(gate187inter2));
  inv1  gate1222(.a(s_96), .O(gate187inter3));
  inv1  gate1223(.a(s_97), .O(gate187inter4));
  nand2 gate1224(.a(gate187inter4), .b(gate187inter3), .O(gate187inter5));
  nor2  gate1225(.a(gate187inter5), .b(gate187inter2), .O(gate187inter6));
  inv1  gate1226(.a(G574), .O(gate187inter7));
  inv1  gate1227(.a(G575), .O(gate187inter8));
  nand2 gate1228(.a(gate187inter8), .b(gate187inter7), .O(gate187inter9));
  nand2 gate1229(.a(s_97), .b(gate187inter3), .O(gate187inter10));
  nor2  gate1230(.a(gate187inter10), .b(gate187inter9), .O(gate187inter11));
  nor2  gate1231(.a(gate187inter11), .b(gate187inter6), .O(gate187inter12));
  nand2 gate1232(.a(gate187inter12), .b(gate187inter1), .O(G612));

  xor2  gate1569(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate1570(.a(gate188inter0), .b(s_146), .O(gate188inter1));
  and2  gate1571(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate1572(.a(s_146), .O(gate188inter3));
  inv1  gate1573(.a(s_147), .O(gate188inter4));
  nand2 gate1574(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate1575(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate1576(.a(G576), .O(gate188inter7));
  inv1  gate1577(.a(G577), .O(gate188inter8));
  nand2 gate1578(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate1579(.a(s_147), .b(gate188inter3), .O(gate188inter10));
  nor2  gate1580(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate1581(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate1582(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );

  xor2  gate1583(.a(G583), .b(G582), .O(gate191inter0));
  nand2 gate1584(.a(gate191inter0), .b(s_148), .O(gate191inter1));
  and2  gate1585(.a(G583), .b(G582), .O(gate191inter2));
  inv1  gate1586(.a(s_148), .O(gate191inter3));
  inv1  gate1587(.a(s_149), .O(gate191inter4));
  nand2 gate1588(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate1589(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate1590(.a(G582), .O(gate191inter7));
  inv1  gate1591(.a(G583), .O(gate191inter8));
  nand2 gate1592(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate1593(.a(s_149), .b(gate191inter3), .O(gate191inter10));
  nor2  gate1594(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate1595(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate1596(.a(gate191inter12), .b(gate191inter1), .O(G632));
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate1163(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate1164(.a(gate193inter0), .b(s_88), .O(gate193inter1));
  and2  gate1165(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate1166(.a(s_88), .O(gate193inter3));
  inv1  gate1167(.a(s_89), .O(gate193inter4));
  nand2 gate1168(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate1169(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate1170(.a(G586), .O(gate193inter7));
  inv1  gate1171(.a(G587), .O(gate193inter8));
  nand2 gate1172(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate1173(.a(s_89), .b(gate193inter3), .O(gate193inter10));
  nor2  gate1174(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate1175(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate1176(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate1135(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate1136(.a(gate195inter0), .b(s_84), .O(gate195inter1));
  and2  gate1137(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate1138(.a(s_84), .O(gate195inter3));
  inv1  gate1139(.a(s_85), .O(gate195inter4));
  nand2 gate1140(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate1141(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate1142(.a(G590), .O(gate195inter7));
  inv1  gate1143(.a(G591), .O(gate195inter8));
  nand2 gate1144(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate1145(.a(s_85), .b(gate195inter3), .O(gate195inter10));
  nor2  gate1146(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate1147(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate1148(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate2647(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate2648(.a(gate197inter0), .b(s_300), .O(gate197inter1));
  and2  gate2649(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate2650(.a(s_300), .O(gate197inter3));
  inv1  gate2651(.a(s_301), .O(gate197inter4));
  nand2 gate2652(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate2653(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate2654(.a(G594), .O(gate197inter7));
  inv1  gate2655(.a(G595), .O(gate197inter8));
  nand2 gate2656(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate2657(.a(s_301), .b(gate197inter3), .O(gate197inter10));
  nor2  gate2658(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate2659(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate2660(.a(gate197inter12), .b(gate197inter1), .O(G654));

  xor2  gate1751(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate1752(.a(gate198inter0), .b(s_172), .O(gate198inter1));
  and2  gate1753(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate1754(.a(s_172), .O(gate198inter3));
  inv1  gate1755(.a(s_173), .O(gate198inter4));
  nand2 gate1756(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate1757(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate1758(.a(G596), .O(gate198inter7));
  inv1  gate1759(.a(G597), .O(gate198inter8));
  nand2 gate1760(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate1761(.a(s_173), .b(gate198inter3), .O(gate198inter10));
  nor2  gate1762(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate1763(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate1764(.a(gate198inter12), .b(gate198inter1), .O(G657));

  xor2  gate1149(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate1150(.a(gate199inter0), .b(s_86), .O(gate199inter1));
  and2  gate1151(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate1152(.a(s_86), .O(gate199inter3));
  inv1  gate1153(.a(s_87), .O(gate199inter4));
  nand2 gate1154(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate1155(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate1156(.a(G598), .O(gate199inter7));
  inv1  gate1157(.a(G599), .O(gate199inter8));
  nand2 gate1158(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate1159(.a(s_87), .b(gate199inter3), .O(gate199inter10));
  nor2  gate1160(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate1161(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate1162(.a(gate199inter12), .b(gate199inter1), .O(G660));

  xor2  gate1485(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate1486(.a(gate200inter0), .b(s_134), .O(gate200inter1));
  and2  gate1487(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate1488(.a(s_134), .O(gate200inter3));
  inv1  gate1489(.a(s_135), .O(gate200inter4));
  nand2 gate1490(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate1491(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate1492(.a(G600), .O(gate200inter7));
  inv1  gate1493(.a(G601), .O(gate200inter8));
  nand2 gate1494(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate1495(.a(s_135), .b(gate200inter3), .O(gate200inter10));
  nor2  gate1496(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate1497(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate1498(.a(gate200inter12), .b(gate200inter1), .O(G663));

  xor2  gate925(.a(G607), .b(G602), .O(gate201inter0));
  nand2 gate926(.a(gate201inter0), .b(s_54), .O(gate201inter1));
  and2  gate927(.a(G607), .b(G602), .O(gate201inter2));
  inv1  gate928(.a(s_54), .O(gate201inter3));
  inv1  gate929(.a(s_55), .O(gate201inter4));
  nand2 gate930(.a(gate201inter4), .b(gate201inter3), .O(gate201inter5));
  nor2  gate931(.a(gate201inter5), .b(gate201inter2), .O(gate201inter6));
  inv1  gate932(.a(G602), .O(gate201inter7));
  inv1  gate933(.a(G607), .O(gate201inter8));
  nand2 gate934(.a(gate201inter8), .b(gate201inter7), .O(gate201inter9));
  nand2 gate935(.a(s_55), .b(gate201inter3), .O(gate201inter10));
  nor2  gate936(.a(gate201inter10), .b(gate201inter9), .O(gate201inter11));
  nor2  gate937(.a(gate201inter11), .b(gate201inter6), .O(gate201inter12));
  nand2 gate938(.a(gate201inter12), .b(gate201inter1), .O(G666));

  xor2  gate1457(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate1458(.a(gate202inter0), .b(s_130), .O(gate202inter1));
  and2  gate1459(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate1460(.a(s_130), .O(gate202inter3));
  inv1  gate1461(.a(s_131), .O(gate202inter4));
  nand2 gate1462(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate1463(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate1464(.a(G612), .O(gate202inter7));
  inv1  gate1465(.a(G617), .O(gate202inter8));
  nand2 gate1466(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate1467(.a(s_131), .b(gate202inter3), .O(gate202inter10));
  nor2  gate1468(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate1469(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate1470(.a(gate202inter12), .b(gate202inter1), .O(G669));

  xor2  gate687(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate688(.a(gate203inter0), .b(s_20), .O(gate203inter1));
  and2  gate689(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate690(.a(s_20), .O(gate203inter3));
  inv1  gate691(.a(s_21), .O(gate203inter4));
  nand2 gate692(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate693(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate694(.a(G602), .O(gate203inter7));
  inv1  gate695(.a(G612), .O(gate203inter8));
  nand2 gate696(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate697(.a(s_21), .b(gate203inter3), .O(gate203inter10));
  nor2  gate698(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate699(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate700(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );

  xor2  gate2423(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate2424(.a(gate206inter0), .b(s_268), .O(gate206inter1));
  and2  gate2425(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate2426(.a(s_268), .O(gate206inter3));
  inv1  gate2427(.a(s_269), .O(gate206inter4));
  nand2 gate2428(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate2429(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate2430(.a(G632), .O(gate206inter7));
  inv1  gate2431(.a(G637), .O(gate206inter8));
  nand2 gate2432(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate2433(.a(s_269), .b(gate206inter3), .O(gate206inter10));
  nor2  gate2434(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate2435(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate2436(.a(gate206inter12), .b(gate206inter1), .O(G681));

  xor2  gate1471(.a(G632), .b(G622), .O(gate207inter0));
  nand2 gate1472(.a(gate207inter0), .b(s_132), .O(gate207inter1));
  and2  gate1473(.a(G632), .b(G622), .O(gate207inter2));
  inv1  gate1474(.a(s_132), .O(gate207inter3));
  inv1  gate1475(.a(s_133), .O(gate207inter4));
  nand2 gate1476(.a(gate207inter4), .b(gate207inter3), .O(gate207inter5));
  nor2  gate1477(.a(gate207inter5), .b(gate207inter2), .O(gate207inter6));
  inv1  gate1478(.a(G622), .O(gate207inter7));
  inv1  gate1479(.a(G632), .O(gate207inter8));
  nand2 gate1480(.a(gate207inter8), .b(gate207inter7), .O(gate207inter9));
  nand2 gate1481(.a(s_133), .b(gate207inter3), .O(gate207inter10));
  nor2  gate1482(.a(gate207inter10), .b(gate207inter9), .O(gate207inter11));
  nor2  gate1483(.a(gate207inter11), .b(gate207inter6), .O(gate207inter12));
  nand2 gate1484(.a(gate207inter12), .b(gate207inter1), .O(G684));

  xor2  gate953(.a(G637), .b(G627), .O(gate208inter0));
  nand2 gate954(.a(gate208inter0), .b(s_58), .O(gate208inter1));
  and2  gate955(.a(G637), .b(G627), .O(gate208inter2));
  inv1  gate956(.a(s_58), .O(gate208inter3));
  inv1  gate957(.a(s_59), .O(gate208inter4));
  nand2 gate958(.a(gate208inter4), .b(gate208inter3), .O(gate208inter5));
  nor2  gate959(.a(gate208inter5), .b(gate208inter2), .O(gate208inter6));
  inv1  gate960(.a(G627), .O(gate208inter7));
  inv1  gate961(.a(G637), .O(gate208inter8));
  nand2 gate962(.a(gate208inter8), .b(gate208inter7), .O(gate208inter9));
  nand2 gate963(.a(s_59), .b(gate208inter3), .O(gate208inter10));
  nor2  gate964(.a(gate208inter10), .b(gate208inter9), .O(gate208inter11));
  nor2  gate965(.a(gate208inter11), .b(gate208inter6), .O(gate208inter12));
  nand2 gate966(.a(gate208inter12), .b(gate208inter1), .O(G687));
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );

  xor2  gate2899(.a(G675), .b(G607), .O(gate215inter0));
  nand2 gate2900(.a(gate215inter0), .b(s_336), .O(gate215inter1));
  and2  gate2901(.a(G675), .b(G607), .O(gate215inter2));
  inv1  gate2902(.a(s_336), .O(gate215inter3));
  inv1  gate2903(.a(s_337), .O(gate215inter4));
  nand2 gate2904(.a(gate215inter4), .b(gate215inter3), .O(gate215inter5));
  nor2  gate2905(.a(gate215inter5), .b(gate215inter2), .O(gate215inter6));
  inv1  gate2906(.a(G607), .O(gate215inter7));
  inv1  gate2907(.a(G675), .O(gate215inter8));
  nand2 gate2908(.a(gate215inter8), .b(gate215inter7), .O(gate215inter9));
  nand2 gate2909(.a(s_337), .b(gate215inter3), .O(gate215inter10));
  nor2  gate2910(.a(gate215inter10), .b(gate215inter9), .O(gate215inter11));
  nor2  gate2911(.a(gate215inter11), .b(gate215inter6), .O(gate215inter12));
  nand2 gate2912(.a(gate215inter12), .b(gate215inter1), .O(G696));

  xor2  gate1079(.a(G675), .b(G617), .O(gate216inter0));
  nand2 gate1080(.a(gate216inter0), .b(s_76), .O(gate216inter1));
  and2  gate1081(.a(G675), .b(G617), .O(gate216inter2));
  inv1  gate1082(.a(s_76), .O(gate216inter3));
  inv1  gate1083(.a(s_77), .O(gate216inter4));
  nand2 gate1084(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate1085(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate1086(.a(G617), .O(gate216inter7));
  inv1  gate1087(.a(G675), .O(gate216inter8));
  nand2 gate1088(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate1089(.a(s_77), .b(gate216inter3), .O(gate216inter10));
  nor2  gate1090(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate1091(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate1092(.a(gate216inter12), .b(gate216inter1), .O(G697));
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );

  xor2  gate1779(.a(G684), .b(G632), .O(gate222inter0));
  nand2 gate1780(.a(gate222inter0), .b(s_176), .O(gate222inter1));
  and2  gate1781(.a(G684), .b(G632), .O(gate222inter2));
  inv1  gate1782(.a(s_176), .O(gate222inter3));
  inv1  gate1783(.a(s_177), .O(gate222inter4));
  nand2 gate1784(.a(gate222inter4), .b(gate222inter3), .O(gate222inter5));
  nor2  gate1785(.a(gate222inter5), .b(gate222inter2), .O(gate222inter6));
  inv1  gate1786(.a(G632), .O(gate222inter7));
  inv1  gate1787(.a(G684), .O(gate222inter8));
  nand2 gate1788(.a(gate222inter8), .b(gate222inter7), .O(gate222inter9));
  nand2 gate1789(.a(s_177), .b(gate222inter3), .O(gate222inter10));
  nor2  gate1790(.a(gate222inter10), .b(gate222inter9), .O(gate222inter11));
  nor2  gate1791(.a(gate222inter11), .b(gate222inter6), .O(gate222inter12));
  nand2 gate1792(.a(gate222inter12), .b(gate222inter1), .O(G703));

  xor2  gate1023(.a(G687), .b(G627), .O(gate223inter0));
  nand2 gate1024(.a(gate223inter0), .b(s_68), .O(gate223inter1));
  and2  gate1025(.a(G687), .b(G627), .O(gate223inter2));
  inv1  gate1026(.a(s_68), .O(gate223inter3));
  inv1  gate1027(.a(s_69), .O(gate223inter4));
  nand2 gate1028(.a(gate223inter4), .b(gate223inter3), .O(gate223inter5));
  nor2  gate1029(.a(gate223inter5), .b(gate223inter2), .O(gate223inter6));
  inv1  gate1030(.a(G627), .O(gate223inter7));
  inv1  gate1031(.a(G687), .O(gate223inter8));
  nand2 gate1032(.a(gate223inter8), .b(gate223inter7), .O(gate223inter9));
  nand2 gate1033(.a(s_69), .b(gate223inter3), .O(gate223inter10));
  nor2  gate1034(.a(gate223inter10), .b(gate223inter9), .O(gate223inter11));
  nor2  gate1035(.a(gate223inter11), .b(gate223inter6), .O(gate223inter12));
  nand2 gate1036(.a(gate223inter12), .b(gate223inter1), .O(G704));
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );

  xor2  gate785(.a(G697), .b(G696), .O(gate228inter0));
  nand2 gate786(.a(gate228inter0), .b(s_34), .O(gate228inter1));
  and2  gate787(.a(G697), .b(G696), .O(gate228inter2));
  inv1  gate788(.a(s_34), .O(gate228inter3));
  inv1  gate789(.a(s_35), .O(gate228inter4));
  nand2 gate790(.a(gate228inter4), .b(gate228inter3), .O(gate228inter5));
  nor2  gate791(.a(gate228inter5), .b(gate228inter2), .O(gate228inter6));
  inv1  gate792(.a(G696), .O(gate228inter7));
  inv1  gate793(.a(G697), .O(gate228inter8));
  nand2 gate794(.a(gate228inter8), .b(gate228inter7), .O(gate228inter9));
  nand2 gate795(.a(s_35), .b(gate228inter3), .O(gate228inter10));
  nor2  gate796(.a(gate228inter10), .b(gate228inter9), .O(gate228inter11));
  nor2  gate797(.a(gate228inter11), .b(gate228inter6), .O(gate228inter12));
  nand2 gate798(.a(gate228inter12), .b(gate228inter1), .O(G715));
nand2 gate229( .a(G698), .b(G699), .O(G718) );

  xor2  gate2983(.a(G701), .b(G700), .O(gate230inter0));
  nand2 gate2984(.a(gate230inter0), .b(s_348), .O(gate230inter1));
  and2  gate2985(.a(G701), .b(G700), .O(gate230inter2));
  inv1  gate2986(.a(s_348), .O(gate230inter3));
  inv1  gate2987(.a(s_349), .O(gate230inter4));
  nand2 gate2988(.a(gate230inter4), .b(gate230inter3), .O(gate230inter5));
  nor2  gate2989(.a(gate230inter5), .b(gate230inter2), .O(gate230inter6));
  inv1  gate2990(.a(G700), .O(gate230inter7));
  inv1  gate2991(.a(G701), .O(gate230inter8));
  nand2 gate2992(.a(gate230inter8), .b(gate230inter7), .O(gate230inter9));
  nand2 gate2993(.a(s_349), .b(gate230inter3), .O(gate230inter10));
  nor2  gate2994(.a(gate230inter10), .b(gate230inter9), .O(gate230inter11));
  nor2  gate2995(.a(gate230inter11), .b(gate230inter6), .O(gate230inter12));
  nand2 gate2996(.a(gate230inter12), .b(gate230inter1), .O(G721));
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );

  xor2  gate2493(.a(G718), .b(G242), .O(gate233inter0));
  nand2 gate2494(.a(gate233inter0), .b(s_278), .O(gate233inter1));
  and2  gate2495(.a(G718), .b(G242), .O(gate233inter2));
  inv1  gate2496(.a(s_278), .O(gate233inter3));
  inv1  gate2497(.a(s_279), .O(gate233inter4));
  nand2 gate2498(.a(gate233inter4), .b(gate233inter3), .O(gate233inter5));
  nor2  gate2499(.a(gate233inter5), .b(gate233inter2), .O(gate233inter6));
  inv1  gate2500(.a(G242), .O(gate233inter7));
  inv1  gate2501(.a(G718), .O(gate233inter8));
  nand2 gate2502(.a(gate233inter8), .b(gate233inter7), .O(gate233inter9));
  nand2 gate2503(.a(s_279), .b(gate233inter3), .O(gate233inter10));
  nor2  gate2504(.a(gate233inter10), .b(gate233inter9), .O(gate233inter11));
  nor2  gate2505(.a(gate233inter11), .b(gate233inter6), .O(gate233inter12));
  nand2 gate2506(.a(gate233inter12), .b(gate233inter1), .O(G730));
nand2 gate234( .a(G245), .b(G721), .O(G733) );

  xor2  gate1317(.a(G724), .b(G248), .O(gate235inter0));
  nand2 gate1318(.a(gate235inter0), .b(s_110), .O(gate235inter1));
  and2  gate1319(.a(G724), .b(G248), .O(gate235inter2));
  inv1  gate1320(.a(s_110), .O(gate235inter3));
  inv1  gate1321(.a(s_111), .O(gate235inter4));
  nand2 gate1322(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate1323(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate1324(.a(G248), .O(gate235inter7));
  inv1  gate1325(.a(G724), .O(gate235inter8));
  nand2 gate1326(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate1327(.a(s_111), .b(gate235inter3), .O(gate235inter10));
  nor2  gate1328(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate1329(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate1330(.a(gate235inter12), .b(gate235inter1), .O(G736));

  xor2  gate2395(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate2396(.a(gate236inter0), .b(s_264), .O(gate236inter1));
  and2  gate2397(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate2398(.a(s_264), .O(gate236inter3));
  inv1  gate2399(.a(s_265), .O(gate236inter4));
  nand2 gate2400(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate2401(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate2402(.a(G251), .O(gate236inter7));
  inv1  gate2403(.a(G727), .O(gate236inter8));
  nand2 gate2404(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate2405(.a(s_265), .b(gate236inter3), .O(gate236inter10));
  nor2  gate2406(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate2407(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate2408(.a(gate236inter12), .b(gate236inter1), .O(G739));

  xor2  gate1905(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate1906(.a(gate237inter0), .b(s_194), .O(gate237inter1));
  and2  gate1907(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate1908(.a(s_194), .O(gate237inter3));
  inv1  gate1909(.a(s_195), .O(gate237inter4));
  nand2 gate1910(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate1911(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate1912(.a(G254), .O(gate237inter7));
  inv1  gate1913(.a(G706), .O(gate237inter8));
  nand2 gate1914(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate1915(.a(s_195), .b(gate237inter3), .O(gate237inter10));
  nor2  gate1916(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate1917(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate1918(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate2885(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate2886(.a(gate240inter0), .b(s_334), .O(gate240inter1));
  and2  gate2887(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate2888(.a(s_334), .O(gate240inter3));
  inv1  gate2889(.a(s_335), .O(gate240inter4));
  nand2 gate2890(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate2891(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate2892(.a(G263), .O(gate240inter7));
  inv1  gate2893(.a(G715), .O(gate240inter8));
  nand2 gate2894(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate2895(.a(s_335), .b(gate240inter3), .O(gate240inter10));
  nor2  gate2896(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate2897(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate2898(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );

  xor2  gate1765(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate1766(.a(gate242inter0), .b(s_174), .O(gate242inter1));
  and2  gate1767(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate1768(.a(s_174), .O(gate242inter3));
  inv1  gate1769(.a(s_175), .O(gate242inter4));
  nand2 gate1770(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate1771(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate1772(.a(G718), .O(gate242inter7));
  inv1  gate1773(.a(G730), .O(gate242inter8));
  nand2 gate1774(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate1775(.a(s_175), .b(gate242inter3), .O(gate242inter10));
  nor2  gate1776(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate1777(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate1778(.a(gate242inter12), .b(gate242inter1), .O(G755));

  xor2  gate813(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate814(.a(gate243inter0), .b(s_38), .O(gate243inter1));
  and2  gate815(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate816(.a(s_38), .O(gate243inter3));
  inv1  gate817(.a(s_39), .O(gate243inter4));
  nand2 gate818(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate819(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate820(.a(G245), .O(gate243inter7));
  inv1  gate821(.a(G733), .O(gate243inter8));
  nand2 gate822(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate823(.a(s_39), .b(gate243inter3), .O(gate243inter10));
  nor2  gate824(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate825(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate826(.a(gate243inter12), .b(gate243inter1), .O(G756));

  xor2  gate2017(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate2018(.a(gate244inter0), .b(s_210), .O(gate244inter1));
  and2  gate2019(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate2020(.a(s_210), .O(gate244inter3));
  inv1  gate2021(.a(s_211), .O(gate244inter4));
  nand2 gate2022(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate2023(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate2024(.a(G721), .O(gate244inter7));
  inv1  gate2025(.a(G733), .O(gate244inter8));
  nand2 gate2026(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate2027(.a(s_211), .b(gate244inter3), .O(gate244inter10));
  nor2  gate2028(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate2029(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate2030(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );

  xor2  gate1919(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate1920(.a(gate247inter0), .b(s_196), .O(gate247inter1));
  and2  gate1921(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate1922(.a(s_196), .O(gate247inter3));
  inv1  gate1923(.a(s_197), .O(gate247inter4));
  nand2 gate1924(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate1925(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate1926(.a(G251), .O(gate247inter7));
  inv1  gate1927(.a(G739), .O(gate247inter8));
  nand2 gate1928(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate1929(.a(s_197), .b(gate247inter3), .O(gate247inter10));
  nor2  gate1930(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate1931(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate1932(.a(gate247inter12), .b(gate247inter1), .O(G760));

  xor2  gate967(.a(G739), .b(G727), .O(gate248inter0));
  nand2 gate968(.a(gate248inter0), .b(s_60), .O(gate248inter1));
  and2  gate969(.a(G739), .b(G727), .O(gate248inter2));
  inv1  gate970(.a(s_60), .O(gate248inter3));
  inv1  gate971(.a(s_61), .O(gate248inter4));
  nand2 gate972(.a(gate248inter4), .b(gate248inter3), .O(gate248inter5));
  nor2  gate973(.a(gate248inter5), .b(gate248inter2), .O(gate248inter6));
  inv1  gate974(.a(G727), .O(gate248inter7));
  inv1  gate975(.a(G739), .O(gate248inter8));
  nand2 gate976(.a(gate248inter8), .b(gate248inter7), .O(gate248inter9));
  nand2 gate977(.a(s_61), .b(gate248inter3), .O(gate248inter10));
  nor2  gate978(.a(gate248inter10), .b(gate248inter9), .O(gate248inter11));
  nor2  gate979(.a(gate248inter11), .b(gate248inter6), .O(gate248inter12));
  nand2 gate980(.a(gate248inter12), .b(gate248inter1), .O(G761));
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );

  xor2  gate1093(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate1094(.a(gate251inter0), .b(s_78), .O(gate251inter1));
  and2  gate1095(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate1096(.a(s_78), .O(gate251inter3));
  inv1  gate1097(.a(s_79), .O(gate251inter4));
  nand2 gate1098(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate1099(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate1100(.a(G257), .O(gate251inter7));
  inv1  gate1101(.a(G745), .O(gate251inter8));
  nand2 gate1102(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate1103(.a(s_79), .b(gate251inter3), .O(gate251inter10));
  nor2  gate1104(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate1105(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate1106(.a(gate251inter12), .b(gate251inter1), .O(G764));

  xor2  gate1009(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate1010(.a(gate252inter0), .b(s_66), .O(gate252inter1));
  and2  gate1011(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate1012(.a(s_66), .O(gate252inter3));
  inv1  gate1013(.a(s_67), .O(gate252inter4));
  nand2 gate1014(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate1015(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate1016(.a(G709), .O(gate252inter7));
  inv1  gate1017(.a(G745), .O(gate252inter8));
  nand2 gate1018(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate1019(.a(s_67), .b(gate252inter3), .O(gate252inter10));
  nor2  gate1020(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate1021(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate1022(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );

  xor2  gate3053(.a(G748), .b(G712), .O(gate254inter0));
  nand2 gate3054(.a(gate254inter0), .b(s_358), .O(gate254inter1));
  and2  gate3055(.a(G748), .b(G712), .O(gate254inter2));
  inv1  gate3056(.a(s_358), .O(gate254inter3));
  inv1  gate3057(.a(s_359), .O(gate254inter4));
  nand2 gate3058(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate3059(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate3060(.a(G712), .O(gate254inter7));
  inv1  gate3061(.a(G748), .O(gate254inter8));
  nand2 gate3062(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate3063(.a(s_359), .b(gate254inter3), .O(gate254inter10));
  nor2  gate3064(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate3065(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate3066(.a(gate254inter12), .b(gate254inter1), .O(G767));

  xor2  gate1261(.a(G751), .b(G263), .O(gate255inter0));
  nand2 gate1262(.a(gate255inter0), .b(s_102), .O(gate255inter1));
  and2  gate1263(.a(G751), .b(G263), .O(gate255inter2));
  inv1  gate1264(.a(s_102), .O(gate255inter3));
  inv1  gate1265(.a(s_103), .O(gate255inter4));
  nand2 gate1266(.a(gate255inter4), .b(gate255inter3), .O(gate255inter5));
  nor2  gate1267(.a(gate255inter5), .b(gate255inter2), .O(gate255inter6));
  inv1  gate1268(.a(G263), .O(gate255inter7));
  inv1  gate1269(.a(G751), .O(gate255inter8));
  nand2 gate1270(.a(gate255inter8), .b(gate255inter7), .O(gate255inter9));
  nand2 gate1271(.a(s_103), .b(gate255inter3), .O(gate255inter10));
  nor2  gate1272(.a(gate255inter10), .b(gate255inter9), .O(gate255inter11));
  nor2  gate1273(.a(gate255inter11), .b(gate255inter6), .O(gate255inter12));
  nand2 gate1274(.a(gate255inter12), .b(gate255inter1), .O(G768));

  xor2  gate2927(.a(G751), .b(G715), .O(gate256inter0));
  nand2 gate2928(.a(gate256inter0), .b(s_340), .O(gate256inter1));
  and2  gate2929(.a(G751), .b(G715), .O(gate256inter2));
  inv1  gate2930(.a(s_340), .O(gate256inter3));
  inv1  gate2931(.a(s_341), .O(gate256inter4));
  nand2 gate2932(.a(gate256inter4), .b(gate256inter3), .O(gate256inter5));
  nor2  gate2933(.a(gate256inter5), .b(gate256inter2), .O(gate256inter6));
  inv1  gate2934(.a(G715), .O(gate256inter7));
  inv1  gate2935(.a(G751), .O(gate256inter8));
  nand2 gate2936(.a(gate256inter8), .b(gate256inter7), .O(gate256inter9));
  nand2 gate2937(.a(s_341), .b(gate256inter3), .O(gate256inter10));
  nor2  gate2938(.a(gate256inter10), .b(gate256inter9), .O(gate256inter11));
  nor2  gate2939(.a(gate256inter11), .b(gate256inter6), .O(gate256inter12));
  nand2 gate2940(.a(gate256inter12), .b(gate256inter1), .O(G769));

  xor2  gate995(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate996(.a(gate257inter0), .b(s_64), .O(gate257inter1));
  and2  gate997(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate998(.a(s_64), .O(gate257inter3));
  inv1  gate999(.a(s_65), .O(gate257inter4));
  nand2 gate1000(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate1001(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate1002(.a(G754), .O(gate257inter7));
  inv1  gate1003(.a(G755), .O(gate257inter8));
  nand2 gate1004(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate1005(.a(s_65), .b(gate257inter3), .O(gate257inter10));
  nor2  gate1006(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate1007(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate1008(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );

  xor2  gate1723(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate1724(.a(gate260inter0), .b(s_168), .O(gate260inter1));
  and2  gate1725(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate1726(.a(s_168), .O(gate260inter3));
  inv1  gate1727(.a(s_169), .O(gate260inter4));
  nand2 gate1728(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate1729(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate1730(.a(G760), .O(gate260inter7));
  inv1  gate1731(.a(G761), .O(gate260inter8));
  nand2 gate1732(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate1733(.a(s_169), .b(gate260inter3), .O(gate260inter10));
  nor2  gate1734(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate1735(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate1736(.a(gate260inter12), .b(gate260inter1), .O(G779));

  xor2  gate2437(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate2438(.a(gate261inter0), .b(s_270), .O(gate261inter1));
  and2  gate2439(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate2440(.a(s_270), .O(gate261inter3));
  inv1  gate2441(.a(s_271), .O(gate261inter4));
  nand2 gate2442(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate2443(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate2444(.a(G762), .O(gate261inter7));
  inv1  gate2445(.a(G763), .O(gate261inter8));
  nand2 gate2446(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate2447(.a(s_271), .b(gate261inter3), .O(gate261inter10));
  nor2  gate2448(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate2449(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate2450(.a(gate261inter12), .b(gate261inter1), .O(G782));
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate2241(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate2242(.a(gate268inter0), .b(s_242), .O(gate268inter1));
  and2  gate2243(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate2244(.a(s_242), .O(gate268inter3));
  inv1  gate2245(.a(s_243), .O(gate268inter4));
  nand2 gate2246(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate2247(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate2248(.a(G651), .O(gate268inter7));
  inv1  gate2249(.a(G779), .O(gate268inter8));
  nand2 gate2250(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate2251(.a(s_243), .b(gate268inter3), .O(gate268inter10));
  nor2  gate2252(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate2253(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate2254(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );

  xor2  gate2521(.a(G785), .b(G657), .O(gate270inter0));
  nand2 gate2522(.a(gate270inter0), .b(s_282), .O(gate270inter1));
  and2  gate2523(.a(G785), .b(G657), .O(gate270inter2));
  inv1  gate2524(.a(s_282), .O(gate270inter3));
  inv1  gate2525(.a(s_283), .O(gate270inter4));
  nand2 gate2526(.a(gate270inter4), .b(gate270inter3), .O(gate270inter5));
  nor2  gate2527(.a(gate270inter5), .b(gate270inter2), .O(gate270inter6));
  inv1  gate2528(.a(G657), .O(gate270inter7));
  inv1  gate2529(.a(G785), .O(gate270inter8));
  nand2 gate2530(.a(gate270inter8), .b(gate270inter7), .O(gate270inter9));
  nand2 gate2531(.a(s_283), .b(gate270inter3), .O(gate270inter10));
  nor2  gate2532(.a(gate270inter10), .b(gate270inter9), .O(gate270inter11));
  nor2  gate2533(.a(gate270inter11), .b(gate270inter6), .O(gate270inter12));
  nand2 gate2534(.a(gate270inter12), .b(gate270inter1), .O(G809));

  xor2  gate2073(.a(G788), .b(G660), .O(gate271inter0));
  nand2 gate2074(.a(gate271inter0), .b(s_218), .O(gate271inter1));
  and2  gate2075(.a(G788), .b(G660), .O(gate271inter2));
  inv1  gate2076(.a(s_218), .O(gate271inter3));
  inv1  gate2077(.a(s_219), .O(gate271inter4));
  nand2 gate2078(.a(gate271inter4), .b(gate271inter3), .O(gate271inter5));
  nor2  gate2079(.a(gate271inter5), .b(gate271inter2), .O(gate271inter6));
  inv1  gate2080(.a(G660), .O(gate271inter7));
  inv1  gate2081(.a(G788), .O(gate271inter8));
  nand2 gate2082(.a(gate271inter8), .b(gate271inter7), .O(gate271inter9));
  nand2 gate2083(.a(s_219), .b(gate271inter3), .O(gate271inter10));
  nor2  gate2084(.a(gate271inter10), .b(gate271inter9), .O(gate271inter11));
  nor2  gate2085(.a(gate271inter11), .b(gate271inter6), .O(gate271inter12));
  nand2 gate2086(.a(gate271inter12), .b(gate271inter1), .O(G812));
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );

  xor2  gate1975(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate1976(.a(gate274inter0), .b(s_204), .O(gate274inter1));
  and2  gate1977(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate1978(.a(s_204), .O(gate274inter3));
  inv1  gate1979(.a(s_205), .O(gate274inter4));
  nand2 gate1980(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate1981(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate1982(.a(G770), .O(gate274inter7));
  inv1  gate1983(.a(G794), .O(gate274inter8));
  nand2 gate1984(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate1985(.a(s_205), .b(gate274inter3), .O(gate274inter10));
  nor2  gate1986(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate1987(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate1988(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );

  xor2  gate757(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate758(.a(gate280inter0), .b(s_30), .O(gate280inter1));
  and2  gate759(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate760(.a(s_30), .O(gate280inter3));
  inv1  gate761(.a(s_31), .O(gate280inter4));
  nand2 gate762(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate763(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate764(.a(G779), .O(gate280inter7));
  inv1  gate765(.a(G803), .O(gate280inter8));
  nand2 gate766(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate767(.a(s_31), .b(gate280inter3), .O(gate280inter10));
  nor2  gate768(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate769(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate770(.a(gate280inter12), .b(gate280inter1), .O(G825));
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );

  xor2  gate1625(.a(G809), .b(G657), .O(gate283inter0));
  nand2 gate1626(.a(gate283inter0), .b(s_154), .O(gate283inter1));
  and2  gate1627(.a(G809), .b(G657), .O(gate283inter2));
  inv1  gate1628(.a(s_154), .O(gate283inter3));
  inv1  gate1629(.a(s_155), .O(gate283inter4));
  nand2 gate1630(.a(gate283inter4), .b(gate283inter3), .O(gate283inter5));
  nor2  gate1631(.a(gate283inter5), .b(gate283inter2), .O(gate283inter6));
  inv1  gate1632(.a(G657), .O(gate283inter7));
  inv1  gate1633(.a(G809), .O(gate283inter8));
  nand2 gate1634(.a(gate283inter8), .b(gate283inter7), .O(gate283inter9));
  nand2 gate1635(.a(s_155), .b(gate283inter3), .O(gate283inter10));
  nor2  gate1636(.a(gate283inter10), .b(gate283inter9), .O(gate283inter11));
  nor2  gate1637(.a(gate283inter11), .b(gate283inter6), .O(gate283inter12));
  nand2 gate1638(.a(gate283inter12), .b(gate283inter1), .O(G828));
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate1793(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate1794(.a(gate285inter0), .b(s_178), .O(gate285inter1));
  and2  gate1795(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate1796(.a(s_178), .O(gate285inter3));
  inv1  gate1797(.a(s_179), .O(gate285inter4));
  nand2 gate1798(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate1799(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate1800(.a(G660), .O(gate285inter7));
  inv1  gate1801(.a(G812), .O(gate285inter8));
  nand2 gate1802(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate1803(.a(s_179), .b(gate285inter3), .O(gate285inter10));
  nor2  gate1804(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate1805(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate1806(.a(gate285inter12), .b(gate285inter1), .O(G830));

  xor2  gate575(.a(G812), .b(G788), .O(gate286inter0));
  nand2 gate576(.a(gate286inter0), .b(s_4), .O(gate286inter1));
  and2  gate577(.a(G812), .b(G788), .O(gate286inter2));
  inv1  gate578(.a(s_4), .O(gate286inter3));
  inv1  gate579(.a(s_5), .O(gate286inter4));
  nand2 gate580(.a(gate286inter4), .b(gate286inter3), .O(gate286inter5));
  nor2  gate581(.a(gate286inter5), .b(gate286inter2), .O(gate286inter6));
  inv1  gate582(.a(G788), .O(gate286inter7));
  inv1  gate583(.a(G812), .O(gate286inter8));
  nand2 gate584(.a(gate286inter8), .b(gate286inter7), .O(gate286inter9));
  nand2 gate585(.a(s_5), .b(gate286inter3), .O(gate286inter10));
  nor2  gate586(.a(gate286inter10), .b(gate286inter9), .O(gate286inter11));
  nor2  gate587(.a(gate286inter11), .b(gate286inter6), .O(gate286inter12));
  nand2 gate588(.a(gate286inter12), .b(gate286inter1), .O(G831));

  xor2  gate1121(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate1122(.a(gate287inter0), .b(s_82), .O(gate287inter1));
  and2  gate1123(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate1124(.a(s_82), .O(gate287inter3));
  inv1  gate1125(.a(s_83), .O(gate287inter4));
  nand2 gate1126(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate1127(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate1128(.a(G663), .O(gate287inter7));
  inv1  gate1129(.a(G815), .O(gate287inter8));
  nand2 gate1130(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate1131(.a(s_83), .b(gate287inter3), .O(gate287inter10));
  nor2  gate1132(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate1133(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate1134(.a(gate287inter12), .b(gate287inter1), .O(G832));
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate2507(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate2508(.a(gate291inter0), .b(s_280), .O(gate291inter1));
  and2  gate2509(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate2510(.a(s_280), .O(gate291inter3));
  inv1  gate2511(.a(s_281), .O(gate291inter4));
  nand2 gate2512(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate2513(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate2514(.a(G822), .O(gate291inter7));
  inv1  gate2515(.a(G823), .O(gate291inter8));
  nand2 gate2516(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate2517(.a(s_281), .b(gate291inter3), .O(gate291inter10));
  nor2  gate2518(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate2519(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate2520(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );

  xor2  gate2871(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate2872(.a(gate293inter0), .b(s_332), .O(gate293inter1));
  and2  gate2873(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate2874(.a(s_332), .O(gate293inter3));
  inv1  gate2875(.a(s_333), .O(gate293inter4));
  nand2 gate2876(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate2877(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate2878(.a(G828), .O(gate293inter7));
  inv1  gate2879(.a(G829), .O(gate293inter8));
  nand2 gate2880(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate2881(.a(s_333), .b(gate293inter3), .O(gate293inter10));
  nor2  gate2882(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate2883(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate2884(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate1065(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate1066(.a(gate295inter0), .b(s_74), .O(gate295inter1));
  and2  gate1067(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate1068(.a(s_74), .O(gate295inter3));
  inv1  gate1069(.a(s_75), .O(gate295inter4));
  nand2 gate1070(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate1071(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate1072(.a(G830), .O(gate295inter7));
  inv1  gate1073(.a(G831), .O(gate295inter8));
  nand2 gate1074(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate1075(.a(s_75), .b(gate295inter3), .O(gate295inter10));
  nor2  gate1076(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate1077(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate1078(.a(gate295inter12), .b(gate295inter1), .O(G912));
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );

  xor2  gate1611(.a(G1039), .b(G2), .O(gate388inter0));
  nand2 gate1612(.a(gate388inter0), .b(s_152), .O(gate388inter1));
  and2  gate1613(.a(G1039), .b(G2), .O(gate388inter2));
  inv1  gate1614(.a(s_152), .O(gate388inter3));
  inv1  gate1615(.a(s_153), .O(gate388inter4));
  nand2 gate1616(.a(gate388inter4), .b(gate388inter3), .O(gate388inter5));
  nor2  gate1617(.a(gate388inter5), .b(gate388inter2), .O(gate388inter6));
  inv1  gate1618(.a(G2), .O(gate388inter7));
  inv1  gate1619(.a(G1039), .O(gate388inter8));
  nand2 gate1620(.a(gate388inter8), .b(gate388inter7), .O(gate388inter9));
  nand2 gate1621(.a(s_153), .b(gate388inter3), .O(gate388inter10));
  nor2  gate1622(.a(gate388inter10), .b(gate388inter9), .O(gate388inter11));
  nor2  gate1623(.a(gate388inter11), .b(gate388inter6), .O(gate388inter12));
  nand2 gate1624(.a(gate388inter12), .b(gate388inter1), .O(G1135));
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate2297(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate2298(.a(gate390inter0), .b(s_250), .O(gate390inter1));
  and2  gate2299(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate2300(.a(s_250), .O(gate390inter3));
  inv1  gate2301(.a(s_251), .O(gate390inter4));
  nand2 gate2302(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate2303(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate2304(.a(G4), .O(gate390inter7));
  inv1  gate2305(.a(G1045), .O(gate390inter8));
  nand2 gate2306(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate2307(.a(s_251), .b(gate390inter3), .O(gate390inter10));
  nor2  gate2308(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate2309(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate2310(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );

  xor2  gate2157(.a(G1057), .b(G8), .O(gate394inter0));
  nand2 gate2158(.a(gate394inter0), .b(s_230), .O(gate394inter1));
  and2  gate2159(.a(G1057), .b(G8), .O(gate394inter2));
  inv1  gate2160(.a(s_230), .O(gate394inter3));
  inv1  gate2161(.a(s_231), .O(gate394inter4));
  nand2 gate2162(.a(gate394inter4), .b(gate394inter3), .O(gate394inter5));
  nor2  gate2163(.a(gate394inter5), .b(gate394inter2), .O(gate394inter6));
  inv1  gate2164(.a(G8), .O(gate394inter7));
  inv1  gate2165(.a(G1057), .O(gate394inter8));
  nand2 gate2166(.a(gate394inter8), .b(gate394inter7), .O(gate394inter9));
  nand2 gate2167(.a(s_231), .b(gate394inter3), .O(gate394inter10));
  nor2  gate2168(.a(gate394inter10), .b(gate394inter9), .O(gate394inter11));
  nor2  gate2169(.a(gate394inter11), .b(gate394inter6), .O(gate394inter12));
  nand2 gate2170(.a(gate394inter12), .b(gate394inter1), .O(G1153));
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );

  xor2  gate2409(.a(G1066), .b(G11), .O(gate397inter0));
  nand2 gate2410(.a(gate397inter0), .b(s_266), .O(gate397inter1));
  and2  gate2411(.a(G1066), .b(G11), .O(gate397inter2));
  inv1  gate2412(.a(s_266), .O(gate397inter3));
  inv1  gate2413(.a(s_267), .O(gate397inter4));
  nand2 gate2414(.a(gate397inter4), .b(gate397inter3), .O(gate397inter5));
  nor2  gate2415(.a(gate397inter5), .b(gate397inter2), .O(gate397inter6));
  inv1  gate2416(.a(G11), .O(gate397inter7));
  inv1  gate2417(.a(G1066), .O(gate397inter8));
  nand2 gate2418(.a(gate397inter8), .b(gate397inter7), .O(gate397inter9));
  nand2 gate2419(.a(s_267), .b(gate397inter3), .O(gate397inter10));
  nor2  gate2420(.a(gate397inter10), .b(gate397inter9), .O(gate397inter11));
  nor2  gate2421(.a(gate397inter11), .b(gate397inter6), .O(gate397inter12));
  nand2 gate2422(.a(gate397inter12), .b(gate397inter1), .O(G1162));
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate2045(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate2046(.a(gate403inter0), .b(s_214), .O(gate403inter1));
  and2  gate2047(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate2048(.a(s_214), .O(gate403inter3));
  inv1  gate2049(.a(s_215), .O(gate403inter4));
  nand2 gate2050(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate2051(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate2052(.a(G17), .O(gate403inter7));
  inv1  gate2053(.a(G1084), .O(gate403inter8));
  nand2 gate2054(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate2055(.a(s_215), .b(gate403inter3), .O(gate403inter10));
  nor2  gate2056(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate2057(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate2058(.a(gate403inter12), .b(gate403inter1), .O(G1180));
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );

  xor2  gate1849(.a(G1090), .b(G19), .O(gate405inter0));
  nand2 gate1850(.a(gate405inter0), .b(s_186), .O(gate405inter1));
  and2  gate1851(.a(G1090), .b(G19), .O(gate405inter2));
  inv1  gate1852(.a(s_186), .O(gate405inter3));
  inv1  gate1853(.a(s_187), .O(gate405inter4));
  nand2 gate1854(.a(gate405inter4), .b(gate405inter3), .O(gate405inter5));
  nor2  gate1855(.a(gate405inter5), .b(gate405inter2), .O(gate405inter6));
  inv1  gate1856(.a(G19), .O(gate405inter7));
  inv1  gate1857(.a(G1090), .O(gate405inter8));
  nand2 gate1858(.a(gate405inter8), .b(gate405inter7), .O(gate405inter9));
  nand2 gate1859(.a(s_187), .b(gate405inter3), .O(gate405inter10));
  nor2  gate1860(.a(gate405inter10), .b(gate405inter9), .O(gate405inter11));
  nor2  gate1861(.a(gate405inter11), .b(gate405inter6), .O(gate405inter12));
  nand2 gate1862(.a(gate405inter12), .b(gate405inter1), .O(G1186));
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );

  xor2  gate2731(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate2732(.a(gate408inter0), .b(s_312), .O(gate408inter1));
  and2  gate2733(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate2734(.a(s_312), .O(gate408inter3));
  inv1  gate2735(.a(s_313), .O(gate408inter4));
  nand2 gate2736(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate2737(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate2738(.a(G22), .O(gate408inter7));
  inv1  gate2739(.a(G1099), .O(gate408inter8));
  nand2 gate2740(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate2741(.a(s_313), .b(gate408inter3), .O(gate408inter10));
  nor2  gate2742(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate2743(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate2744(.a(gate408inter12), .b(gate408inter1), .O(G1195));
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate2059(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate2060(.a(gate411inter0), .b(s_216), .O(gate411inter1));
  and2  gate2061(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate2062(.a(s_216), .O(gate411inter3));
  inv1  gate2063(.a(s_217), .O(gate411inter4));
  nand2 gate2064(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate2065(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate2066(.a(G25), .O(gate411inter7));
  inv1  gate2067(.a(G1108), .O(gate411inter8));
  nand2 gate2068(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate2069(.a(s_217), .b(gate411inter3), .O(gate411inter10));
  nor2  gate2070(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate2071(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate2072(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );

  xor2  gate2605(.a(G1114), .b(G27), .O(gate413inter0));
  nand2 gate2606(.a(gate413inter0), .b(s_294), .O(gate413inter1));
  and2  gate2607(.a(G1114), .b(G27), .O(gate413inter2));
  inv1  gate2608(.a(s_294), .O(gate413inter3));
  inv1  gate2609(.a(s_295), .O(gate413inter4));
  nand2 gate2610(.a(gate413inter4), .b(gate413inter3), .O(gate413inter5));
  nor2  gate2611(.a(gate413inter5), .b(gate413inter2), .O(gate413inter6));
  inv1  gate2612(.a(G27), .O(gate413inter7));
  inv1  gate2613(.a(G1114), .O(gate413inter8));
  nand2 gate2614(.a(gate413inter8), .b(gate413inter7), .O(gate413inter9));
  nand2 gate2615(.a(s_295), .b(gate413inter3), .O(gate413inter10));
  nor2  gate2616(.a(gate413inter10), .b(gate413inter9), .O(gate413inter11));
  nor2  gate2617(.a(gate413inter11), .b(gate413inter6), .O(gate413inter12));
  nand2 gate2618(.a(gate413inter12), .b(gate413inter1), .O(G1210));
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate2689(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate2690(.a(gate420inter0), .b(s_306), .O(gate420inter1));
  and2  gate2691(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate2692(.a(s_306), .O(gate420inter3));
  inv1  gate2693(.a(s_307), .O(gate420inter4));
  nand2 gate2694(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate2695(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate2696(.a(G1036), .O(gate420inter7));
  inv1  gate2697(.a(G1132), .O(gate420inter8));
  nand2 gate2698(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate2699(.a(s_307), .b(gate420inter3), .O(gate420inter10));
  nor2  gate2700(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate2701(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate2702(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate1331(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate1332(.a(gate422inter0), .b(s_112), .O(gate422inter1));
  and2  gate1333(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate1334(.a(s_112), .O(gate422inter3));
  inv1  gate1335(.a(s_113), .O(gate422inter4));
  nand2 gate1336(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate1337(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate1338(.a(G1039), .O(gate422inter7));
  inv1  gate1339(.a(G1135), .O(gate422inter8));
  nand2 gate1340(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate1341(.a(s_113), .b(gate422inter3), .O(gate422inter10));
  nor2  gate1342(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate1343(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate1344(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );

  xor2  gate2003(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate2004(.a(gate424inter0), .b(s_208), .O(gate424inter1));
  and2  gate2005(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate2006(.a(s_208), .O(gate424inter3));
  inv1  gate2007(.a(s_209), .O(gate424inter4));
  nand2 gate2008(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate2009(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate2010(.a(G1042), .O(gate424inter7));
  inv1  gate2011(.a(G1138), .O(gate424inter8));
  nand2 gate2012(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate2013(.a(s_209), .b(gate424inter3), .O(gate424inter10));
  nor2  gate2014(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate2015(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate2016(.a(gate424inter12), .b(gate424inter1), .O(G1233));

  xor2  gate603(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate604(.a(gate425inter0), .b(s_8), .O(gate425inter1));
  and2  gate605(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate606(.a(s_8), .O(gate425inter3));
  inv1  gate607(.a(s_9), .O(gate425inter4));
  nand2 gate608(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate609(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate610(.a(G4), .O(gate425inter7));
  inv1  gate611(.a(G1141), .O(gate425inter8));
  nand2 gate612(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate613(.a(s_9), .b(gate425inter3), .O(gate425inter10));
  nor2  gate614(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate615(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate616(.a(gate425inter12), .b(gate425inter1), .O(G1234));
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );

  xor2  gate1359(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate1360(.a(gate427inter0), .b(s_116), .O(gate427inter1));
  and2  gate1361(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate1362(.a(s_116), .O(gate427inter3));
  inv1  gate1363(.a(s_117), .O(gate427inter4));
  nand2 gate1364(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate1365(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate1366(.a(G5), .O(gate427inter7));
  inv1  gate1367(.a(G1144), .O(gate427inter8));
  nand2 gate1368(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate1369(.a(s_117), .b(gate427inter3), .O(gate427inter10));
  nor2  gate1370(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate1371(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate1372(.a(gate427inter12), .b(gate427inter1), .O(G1236));

  xor2  gate1961(.a(G1144), .b(G1048), .O(gate428inter0));
  nand2 gate1962(.a(gate428inter0), .b(s_202), .O(gate428inter1));
  and2  gate1963(.a(G1144), .b(G1048), .O(gate428inter2));
  inv1  gate1964(.a(s_202), .O(gate428inter3));
  inv1  gate1965(.a(s_203), .O(gate428inter4));
  nand2 gate1966(.a(gate428inter4), .b(gate428inter3), .O(gate428inter5));
  nor2  gate1967(.a(gate428inter5), .b(gate428inter2), .O(gate428inter6));
  inv1  gate1968(.a(G1048), .O(gate428inter7));
  inv1  gate1969(.a(G1144), .O(gate428inter8));
  nand2 gate1970(.a(gate428inter8), .b(gate428inter7), .O(gate428inter9));
  nand2 gate1971(.a(s_203), .b(gate428inter3), .O(gate428inter10));
  nor2  gate1972(.a(gate428inter10), .b(gate428inter9), .O(gate428inter11));
  nor2  gate1973(.a(gate428inter11), .b(gate428inter6), .O(gate428inter12));
  nand2 gate1974(.a(gate428inter12), .b(gate428inter1), .O(G1237));
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate2745(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate2746(.a(gate430inter0), .b(s_314), .O(gate430inter1));
  and2  gate2747(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate2748(.a(s_314), .O(gate430inter3));
  inv1  gate2749(.a(s_315), .O(gate430inter4));
  nand2 gate2750(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate2751(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate2752(.a(G1051), .O(gate430inter7));
  inv1  gate2753(.a(G1147), .O(gate430inter8));
  nand2 gate2754(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate2755(.a(s_315), .b(gate430inter3), .O(gate430inter10));
  nor2  gate2756(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate2757(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate2758(.a(gate430inter12), .b(gate430inter1), .O(G1239));

  xor2  gate1275(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate1276(.a(gate431inter0), .b(s_104), .O(gate431inter1));
  and2  gate1277(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate1278(.a(s_104), .O(gate431inter3));
  inv1  gate1279(.a(s_105), .O(gate431inter4));
  nand2 gate1280(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate1281(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate1282(.a(G7), .O(gate431inter7));
  inv1  gate1283(.a(G1150), .O(gate431inter8));
  nand2 gate1284(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate1285(.a(s_105), .b(gate431inter3), .O(gate431inter10));
  nor2  gate1286(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate1287(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate1288(.a(gate431inter12), .b(gate431inter1), .O(G1240));

  xor2  gate911(.a(G1150), .b(G1054), .O(gate432inter0));
  nand2 gate912(.a(gate432inter0), .b(s_52), .O(gate432inter1));
  and2  gate913(.a(G1150), .b(G1054), .O(gate432inter2));
  inv1  gate914(.a(s_52), .O(gate432inter3));
  inv1  gate915(.a(s_53), .O(gate432inter4));
  nand2 gate916(.a(gate432inter4), .b(gate432inter3), .O(gate432inter5));
  nor2  gate917(.a(gate432inter5), .b(gate432inter2), .O(gate432inter6));
  inv1  gate918(.a(G1054), .O(gate432inter7));
  inv1  gate919(.a(G1150), .O(gate432inter8));
  nand2 gate920(.a(gate432inter8), .b(gate432inter7), .O(gate432inter9));
  nand2 gate921(.a(s_53), .b(gate432inter3), .O(gate432inter10));
  nor2  gate922(.a(gate432inter10), .b(gate432inter9), .O(gate432inter11));
  nor2  gate923(.a(gate432inter11), .b(gate432inter6), .O(gate432inter12));
  nand2 gate924(.a(gate432inter12), .b(gate432inter1), .O(G1241));

  xor2  gate1653(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate1654(.a(gate433inter0), .b(s_158), .O(gate433inter1));
  and2  gate1655(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate1656(.a(s_158), .O(gate433inter3));
  inv1  gate1657(.a(s_159), .O(gate433inter4));
  nand2 gate1658(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate1659(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate1660(.a(G8), .O(gate433inter7));
  inv1  gate1661(.a(G1153), .O(gate433inter8));
  nand2 gate1662(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate1663(.a(s_159), .b(gate433inter3), .O(gate433inter10));
  nor2  gate1664(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate1665(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate1666(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate1681(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate1682(.a(gate439inter0), .b(s_162), .O(gate439inter1));
  and2  gate1683(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate1684(.a(s_162), .O(gate439inter3));
  inv1  gate1685(.a(s_163), .O(gate439inter4));
  nand2 gate1686(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate1687(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate1688(.a(G11), .O(gate439inter7));
  inv1  gate1689(.a(G1162), .O(gate439inter8));
  nand2 gate1690(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate1691(.a(s_163), .b(gate439inter3), .O(gate439inter10));
  nor2  gate1692(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate1693(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate1694(.a(gate439inter12), .b(gate439inter1), .O(G1248));

  xor2  gate2353(.a(G1162), .b(G1066), .O(gate440inter0));
  nand2 gate2354(.a(gate440inter0), .b(s_258), .O(gate440inter1));
  and2  gate2355(.a(G1162), .b(G1066), .O(gate440inter2));
  inv1  gate2356(.a(s_258), .O(gate440inter3));
  inv1  gate2357(.a(s_259), .O(gate440inter4));
  nand2 gate2358(.a(gate440inter4), .b(gate440inter3), .O(gate440inter5));
  nor2  gate2359(.a(gate440inter5), .b(gate440inter2), .O(gate440inter6));
  inv1  gate2360(.a(G1066), .O(gate440inter7));
  inv1  gate2361(.a(G1162), .O(gate440inter8));
  nand2 gate2362(.a(gate440inter8), .b(gate440inter7), .O(gate440inter9));
  nand2 gate2363(.a(s_259), .b(gate440inter3), .O(gate440inter10));
  nor2  gate2364(.a(gate440inter10), .b(gate440inter9), .O(gate440inter11));
  nor2  gate2365(.a(gate440inter11), .b(gate440inter6), .O(gate440inter12));
  nand2 gate2366(.a(gate440inter12), .b(gate440inter1), .O(G1249));
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate1891(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate1892(.a(gate442inter0), .b(s_192), .O(gate442inter1));
  and2  gate1893(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate1894(.a(s_192), .O(gate442inter3));
  inv1  gate1895(.a(s_193), .O(gate442inter4));
  nand2 gate1896(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate1897(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate1898(.a(G1069), .O(gate442inter7));
  inv1  gate1899(.a(G1165), .O(gate442inter8));
  nand2 gate1900(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate1901(.a(s_193), .b(gate442inter3), .O(gate442inter10));
  nor2  gate1902(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate1903(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate1904(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );

  xor2  gate3067(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate3068(.a(gate446inter0), .b(s_360), .O(gate446inter1));
  and2  gate3069(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate3070(.a(s_360), .O(gate446inter3));
  inv1  gate3071(.a(s_361), .O(gate446inter4));
  nand2 gate3072(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate3073(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate3074(.a(G1075), .O(gate446inter7));
  inv1  gate3075(.a(G1171), .O(gate446inter8));
  nand2 gate3076(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate3077(.a(s_361), .b(gate446inter3), .O(gate446inter10));
  nor2  gate3078(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate3079(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate3080(.a(gate446inter12), .b(gate446inter1), .O(G1255));
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );

  xor2  gate2717(.a(G1180), .b(G1084), .O(gate452inter0));
  nand2 gate2718(.a(gate452inter0), .b(s_310), .O(gate452inter1));
  and2  gate2719(.a(G1180), .b(G1084), .O(gate452inter2));
  inv1  gate2720(.a(s_310), .O(gate452inter3));
  inv1  gate2721(.a(s_311), .O(gate452inter4));
  nand2 gate2722(.a(gate452inter4), .b(gate452inter3), .O(gate452inter5));
  nor2  gate2723(.a(gate452inter5), .b(gate452inter2), .O(gate452inter6));
  inv1  gate2724(.a(G1084), .O(gate452inter7));
  inv1  gate2725(.a(G1180), .O(gate452inter8));
  nand2 gate2726(.a(gate452inter8), .b(gate452inter7), .O(gate452inter9));
  nand2 gate2727(.a(s_311), .b(gate452inter3), .O(gate452inter10));
  nor2  gate2728(.a(gate452inter10), .b(gate452inter9), .O(gate452inter11));
  nor2  gate2729(.a(gate452inter11), .b(gate452inter6), .O(gate452inter12));
  nand2 gate2730(.a(gate452inter12), .b(gate452inter1), .O(G1261));
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );

  xor2  gate1499(.a(G1189), .b(G20), .O(gate457inter0));
  nand2 gate1500(.a(gate457inter0), .b(s_136), .O(gate457inter1));
  and2  gate1501(.a(G1189), .b(G20), .O(gate457inter2));
  inv1  gate1502(.a(s_136), .O(gate457inter3));
  inv1  gate1503(.a(s_137), .O(gate457inter4));
  nand2 gate1504(.a(gate457inter4), .b(gate457inter3), .O(gate457inter5));
  nor2  gate1505(.a(gate457inter5), .b(gate457inter2), .O(gate457inter6));
  inv1  gate1506(.a(G20), .O(gate457inter7));
  inv1  gate1507(.a(G1189), .O(gate457inter8));
  nand2 gate1508(.a(gate457inter8), .b(gate457inter7), .O(gate457inter9));
  nand2 gate1509(.a(s_137), .b(gate457inter3), .O(gate457inter10));
  nor2  gate1510(.a(gate457inter10), .b(gate457inter9), .O(gate457inter11));
  nor2  gate1511(.a(gate457inter11), .b(gate457inter6), .O(gate457inter12));
  nand2 gate1512(.a(gate457inter12), .b(gate457inter1), .O(G1266));
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate2787(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate2788(.a(gate460inter0), .b(s_320), .O(gate460inter1));
  and2  gate2789(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate2790(.a(s_320), .O(gate460inter3));
  inv1  gate2791(.a(s_321), .O(gate460inter4));
  nand2 gate2792(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate2793(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate2794(.a(G1096), .O(gate460inter7));
  inv1  gate2795(.a(G1192), .O(gate460inter8));
  nand2 gate2796(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate2797(.a(s_321), .b(gate460inter3), .O(gate460inter10));
  nor2  gate2798(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate2799(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate2800(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );

  xor2  gate1107(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate1108(.a(gate462inter0), .b(s_80), .O(gate462inter1));
  and2  gate1109(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate1110(.a(s_80), .O(gate462inter3));
  inv1  gate1111(.a(s_81), .O(gate462inter4));
  nand2 gate1112(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate1113(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate1114(.a(G1099), .O(gate462inter7));
  inv1  gate1115(.a(G1195), .O(gate462inter8));
  nand2 gate1116(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate1117(.a(s_81), .b(gate462inter3), .O(gate462inter10));
  nor2  gate1118(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate1119(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate1120(.a(gate462inter12), .b(gate462inter1), .O(G1271));

  xor2  gate2675(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate2676(.a(gate463inter0), .b(s_304), .O(gate463inter1));
  and2  gate2677(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate2678(.a(s_304), .O(gate463inter3));
  inv1  gate2679(.a(s_305), .O(gate463inter4));
  nand2 gate2680(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate2681(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate2682(.a(G23), .O(gate463inter7));
  inv1  gate2683(.a(G1198), .O(gate463inter8));
  nand2 gate2684(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate2685(.a(s_305), .b(gate463inter3), .O(gate463inter10));
  nor2  gate2686(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate2687(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate2688(.a(gate463inter12), .b(gate463inter1), .O(G1272));

  xor2  gate2843(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate2844(.a(gate464inter0), .b(s_328), .O(gate464inter1));
  and2  gate2845(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate2846(.a(s_328), .O(gate464inter3));
  inv1  gate2847(.a(s_329), .O(gate464inter4));
  nand2 gate2848(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate2849(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate2850(.a(G1102), .O(gate464inter7));
  inv1  gate2851(.a(G1198), .O(gate464inter8));
  nand2 gate2852(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate2853(.a(s_329), .b(gate464inter3), .O(gate464inter10));
  nor2  gate2854(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate2855(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate2856(.a(gate464inter12), .b(gate464inter1), .O(G1273));

  xor2  gate2339(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate2340(.a(gate465inter0), .b(s_256), .O(gate465inter1));
  and2  gate2341(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate2342(.a(s_256), .O(gate465inter3));
  inv1  gate2343(.a(s_257), .O(gate465inter4));
  nand2 gate2344(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate2345(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate2346(.a(G24), .O(gate465inter7));
  inv1  gate2347(.a(G1201), .O(gate465inter8));
  nand2 gate2348(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate2349(.a(s_257), .b(gate465inter3), .O(gate465inter10));
  nor2  gate2350(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate2351(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate2352(.a(gate465inter12), .b(gate465inter1), .O(G1274));

  xor2  gate2815(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate2816(.a(gate466inter0), .b(s_324), .O(gate466inter1));
  and2  gate2817(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate2818(.a(s_324), .O(gate466inter3));
  inv1  gate2819(.a(s_325), .O(gate466inter4));
  nand2 gate2820(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate2821(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate2822(.a(G1105), .O(gate466inter7));
  inv1  gate2823(.a(G1201), .O(gate466inter8));
  nand2 gate2824(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate2825(.a(s_325), .b(gate466inter3), .O(gate466inter10));
  nor2  gate2826(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate2827(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate2828(.a(gate466inter12), .b(gate466inter1), .O(G1275));

  xor2  gate2829(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate2830(.a(gate467inter0), .b(s_326), .O(gate467inter1));
  and2  gate2831(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate2832(.a(s_326), .O(gate467inter3));
  inv1  gate2833(.a(s_327), .O(gate467inter4));
  nand2 gate2834(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate2835(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate2836(.a(G25), .O(gate467inter7));
  inv1  gate2837(.a(G1204), .O(gate467inter8));
  nand2 gate2838(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate2839(.a(s_327), .b(gate467inter3), .O(gate467inter10));
  nor2  gate2840(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate2841(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate2842(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate1415(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate1416(.a(gate472inter0), .b(s_124), .O(gate472inter1));
  and2  gate1417(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate1418(.a(s_124), .O(gate472inter3));
  inv1  gate1419(.a(s_125), .O(gate472inter4));
  nand2 gate1420(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate1421(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate1422(.a(G1114), .O(gate472inter7));
  inv1  gate1423(.a(G1210), .O(gate472inter8));
  nand2 gate1424(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate1425(.a(s_125), .b(gate472inter3), .O(gate472inter10));
  nor2  gate1426(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate1427(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate1428(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate2381(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate2382(.a(gate480inter0), .b(s_262), .O(gate480inter1));
  and2  gate2383(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate2384(.a(s_262), .O(gate480inter3));
  inv1  gate2385(.a(s_263), .O(gate480inter4));
  nand2 gate2386(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate2387(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate2388(.a(G1126), .O(gate480inter7));
  inv1  gate2389(.a(G1222), .O(gate480inter8));
  nand2 gate2390(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate2391(.a(s_263), .b(gate480inter3), .O(gate480inter10));
  nor2  gate2392(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate2393(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate2394(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate1037(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate1038(.a(gate485inter0), .b(s_70), .O(gate485inter1));
  and2  gate1039(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate1040(.a(s_70), .O(gate485inter3));
  inv1  gate1041(.a(s_71), .O(gate485inter4));
  nand2 gate1042(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate1043(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate1044(.a(G1232), .O(gate485inter7));
  inv1  gate1045(.a(G1233), .O(gate485inter8));
  nand2 gate1046(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate1047(.a(s_71), .b(gate485inter3), .O(gate485inter10));
  nor2  gate1048(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate1049(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate1050(.a(gate485inter12), .b(gate485inter1), .O(G1294));
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate1527(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate1528(.a(gate492inter0), .b(s_140), .O(gate492inter1));
  and2  gate1529(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate1530(.a(s_140), .O(gate492inter3));
  inv1  gate1531(.a(s_141), .O(gate492inter4));
  nand2 gate1532(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate1533(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate1534(.a(G1246), .O(gate492inter7));
  inv1  gate1535(.a(G1247), .O(gate492inter8));
  nand2 gate1536(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate1537(.a(s_141), .b(gate492inter3), .O(gate492inter10));
  nor2  gate1538(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate1539(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate1540(.a(gate492inter12), .b(gate492inter1), .O(G1301));
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );

  xor2  gate1709(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate1710(.a(gate495inter0), .b(s_166), .O(gate495inter1));
  and2  gate1711(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate1712(.a(s_166), .O(gate495inter3));
  inv1  gate1713(.a(s_167), .O(gate495inter4));
  nand2 gate1714(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate1715(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate1716(.a(G1252), .O(gate495inter7));
  inv1  gate1717(.a(G1253), .O(gate495inter8));
  nand2 gate1718(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate1719(.a(s_167), .b(gate495inter3), .O(gate495inter10));
  nor2  gate1720(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate1721(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate1722(.a(gate495inter12), .b(gate495inter1), .O(G1304));

  xor2  gate701(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate702(.a(gate496inter0), .b(s_22), .O(gate496inter1));
  and2  gate703(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate704(.a(s_22), .O(gate496inter3));
  inv1  gate705(.a(s_23), .O(gate496inter4));
  nand2 gate706(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate707(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate708(.a(G1254), .O(gate496inter7));
  inv1  gate709(.a(G1255), .O(gate496inter8));
  nand2 gate710(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate711(.a(s_23), .b(gate496inter3), .O(gate496inter10));
  nor2  gate712(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate713(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate714(.a(gate496inter12), .b(gate496inter1), .O(G1305));
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );

  xor2  gate869(.a(G1259), .b(G1258), .O(gate498inter0));
  nand2 gate870(.a(gate498inter0), .b(s_46), .O(gate498inter1));
  and2  gate871(.a(G1259), .b(G1258), .O(gate498inter2));
  inv1  gate872(.a(s_46), .O(gate498inter3));
  inv1  gate873(.a(s_47), .O(gate498inter4));
  nand2 gate874(.a(gate498inter4), .b(gate498inter3), .O(gate498inter5));
  nor2  gate875(.a(gate498inter5), .b(gate498inter2), .O(gate498inter6));
  inv1  gate876(.a(G1258), .O(gate498inter7));
  inv1  gate877(.a(G1259), .O(gate498inter8));
  nand2 gate878(.a(gate498inter8), .b(gate498inter7), .O(gate498inter9));
  nand2 gate879(.a(s_47), .b(gate498inter3), .O(gate498inter10));
  nor2  gate880(.a(gate498inter10), .b(gate498inter9), .O(gate498inter11));
  nor2  gate881(.a(gate498inter11), .b(gate498inter6), .O(gate498inter12));
  nand2 gate882(.a(gate498inter12), .b(gate498inter1), .O(G1307));
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );

  xor2  gate2479(.a(G1263), .b(G1262), .O(gate500inter0));
  nand2 gate2480(.a(gate500inter0), .b(s_276), .O(gate500inter1));
  and2  gate2481(.a(G1263), .b(G1262), .O(gate500inter2));
  inv1  gate2482(.a(s_276), .O(gate500inter3));
  inv1  gate2483(.a(s_277), .O(gate500inter4));
  nand2 gate2484(.a(gate500inter4), .b(gate500inter3), .O(gate500inter5));
  nor2  gate2485(.a(gate500inter5), .b(gate500inter2), .O(gate500inter6));
  inv1  gate2486(.a(G1262), .O(gate500inter7));
  inv1  gate2487(.a(G1263), .O(gate500inter8));
  nand2 gate2488(.a(gate500inter8), .b(gate500inter7), .O(gate500inter9));
  nand2 gate2489(.a(s_277), .b(gate500inter3), .O(gate500inter10));
  nor2  gate2490(.a(gate500inter10), .b(gate500inter9), .O(gate500inter11));
  nor2  gate2491(.a(gate500inter11), .b(gate500inter6), .O(gate500inter12));
  nand2 gate2492(.a(gate500inter12), .b(gate500inter1), .O(G1309));
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate547(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate548(.a(gate504inter0), .b(s_0), .O(gate504inter1));
  and2  gate549(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate550(.a(s_0), .O(gate504inter3));
  inv1  gate551(.a(s_1), .O(gate504inter4));
  nand2 gate552(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate553(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate554(.a(G1270), .O(gate504inter7));
  inv1  gate555(.a(G1271), .O(gate504inter8));
  nand2 gate556(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate557(.a(s_1), .b(gate504inter3), .O(gate504inter10));
  nor2  gate558(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate559(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate560(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );

  xor2  gate855(.a(G1275), .b(G1274), .O(gate506inter0));
  nand2 gate856(.a(gate506inter0), .b(s_44), .O(gate506inter1));
  and2  gate857(.a(G1275), .b(G1274), .O(gate506inter2));
  inv1  gate858(.a(s_44), .O(gate506inter3));
  inv1  gate859(.a(s_45), .O(gate506inter4));
  nand2 gate860(.a(gate506inter4), .b(gate506inter3), .O(gate506inter5));
  nor2  gate861(.a(gate506inter5), .b(gate506inter2), .O(gate506inter6));
  inv1  gate862(.a(G1274), .O(gate506inter7));
  inv1  gate863(.a(G1275), .O(gate506inter8));
  nand2 gate864(.a(gate506inter8), .b(gate506inter7), .O(gate506inter9));
  nand2 gate865(.a(s_45), .b(gate506inter3), .O(gate506inter10));
  nor2  gate866(.a(gate506inter10), .b(gate506inter9), .O(gate506inter11));
  nor2  gate867(.a(gate506inter11), .b(gate506inter6), .O(gate506inter12));
  nand2 gate868(.a(gate506inter12), .b(gate506inter1), .O(G1315));
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );

  xor2  gate1177(.a(G1281), .b(G1280), .O(gate509inter0));
  nand2 gate1178(.a(gate509inter0), .b(s_90), .O(gate509inter1));
  and2  gate1179(.a(G1281), .b(G1280), .O(gate509inter2));
  inv1  gate1180(.a(s_90), .O(gate509inter3));
  inv1  gate1181(.a(s_91), .O(gate509inter4));
  nand2 gate1182(.a(gate509inter4), .b(gate509inter3), .O(gate509inter5));
  nor2  gate1183(.a(gate509inter5), .b(gate509inter2), .O(gate509inter6));
  inv1  gate1184(.a(G1280), .O(gate509inter7));
  inv1  gate1185(.a(G1281), .O(gate509inter8));
  nand2 gate1186(.a(gate509inter8), .b(gate509inter7), .O(gate509inter9));
  nand2 gate1187(.a(s_91), .b(gate509inter3), .O(gate509inter10));
  nor2  gate1188(.a(gate509inter10), .b(gate509inter9), .O(gate509inter11));
  nor2  gate1189(.a(gate509inter11), .b(gate509inter6), .O(gate509inter12));
  nand2 gate1190(.a(gate509inter12), .b(gate509inter1), .O(G1318));
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );

  xor2  gate2115(.a(G1287), .b(G1286), .O(gate512inter0));
  nand2 gate2116(.a(gate512inter0), .b(s_224), .O(gate512inter1));
  and2  gate2117(.a(G1287), .b(G1286), .O(gate512inter2));
  inv1  gate2118(.a(s_224), .O(gate512inter3));
  inv1  gate2119(.a(s_225), .O(gate512inter4));
  nand2 gate2120(.a(gate512inter4), .b(gate512inter3), .O(gate512inter5));
  nor2  gate2121(.a(gate512inter5), .b(gate512inter2), .O(gate512inter6));
  inv1  gate2122(.a(G1286), .O(gate512inter7));
  inv1  gate2123(.a(G1287), .O(gate512inter8));
  nand2 gate2124(.a(gate512inter8), .b(gate512inter7), .O(gate512inter9));
  nand2 gate2125(.a(s_225), .b(gate512inter3), .O(gate512inter10));
  nor2  gate2126(.a(gate512inter10), .b(gate512inter9), .O(gate512inter11));
  nor2  gate2127(.a(gate512inter11), .b(gate512inter6), .O(gate512inter12));
  nand2 gate2128(.a(gate512inter12), .b(gate512inter1), .O(G1321));
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule