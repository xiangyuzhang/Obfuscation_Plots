module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate495inter0, gate495inter1, gate495inter2, gate495inter3, gate495inter4, gate495inter5, gate495inter6, gate495inter7, gate495inter8, gate495inter9, gate495inter10, gate495inter11, gate495inter12, gate249inter0, gate249inter1, gate249inter2, gate249inter3, gate249inter4, gate249inter5, gate249inter6, gate249inter7, gate249inter8, gate249inter9, gate249inter10, gate249inter11, gate249inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate156inter0, gate156inter1, gate156inter2, gate156inter3, gate156inter4, gate156inter5, gate156inter6, gate156inter7, gate156inter8, gate156inter9, gate156inter10, gate156inter11, gate156inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate120inter0, gate120inter1, gate120inter2, gate120inter3, gate120inter4, gate120inter5, gate120inter6, gate120inter7, gate120inter8, gate120inter9, gate120inter10, gate120inter11, gate120inter12, gate438inter0, gate438inter1, gate438inter2, gate438inter3, gate438inter4, gate438inter5, gate438inter6, gate438inter7, gate438inter8, gate438inter9, gate438inter10, gate438inter11, gate438inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate465inter0, gate465inter1, gate465inter2, gate465inter3, gate465inter4, gate465inter5, gate465inter6, gate465inter7, gate465inter8, gate465inter9, gate465inter10, gate465inter11, gate465inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate75inter0, gate75inter1, gate75inter2, gate75inter3, gate75inter4, gate75inter5, gate75inter6, gate75inter7, gate75inter8, gate75inter9, gate75inter10, gate75inter11, gate75inter12, gate146inter0, gate146inter1, gate146inter2, gate146inter3, gate146inter4, gate146inter5, gate146inter6, gate146inter7, gate146inter8, gate146inter9, gate146inter10, gate146inter11, gate146inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate411inter0, gate411inter1, gate411inter2, gate411inter3, gate411inter4, gate411inter5, gate411inter6, gate411inter7, gate411inter8, gate411inter9, gate411inter10, gate411inter11, gate411inter12, gate444inter0, gate444inter1, gate444inter2, gate444inter3, gate444inter4, gate444inter5, gate444inter6, gate444inter7, gate444inter8, gate444inter9, gate444inter10, gate444inter11, gate444inter12, gate110inter0, gate110inter1, gate110inter2, gate110inter3, gate110inter4, gate110inter5, gate110inter6, gate110inter7, gate110inter8, gate110inter9, gate110inter10, gate110inter11, gate110inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate95inter0, gate95inter1, gate95inter2, gate95inter3, gate95inter4, gate95inter5, gate95inter6, gate95inter7, gate95inter8, gate95inter9, gate95inter10, gate95inter11, gate95inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate118inter0, gate118inter1, gate118inter2, gate118inter3, gate118inter4, gate118inter5, gate118inter6, gate118inter7, gate118inter8, gate118inter9, gate118inter10, gate118inter11, gate118inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate211inter0, gate211inter1, gate211inter2, gate211inter3, gate211inter4, gate211inter5, gate211inter6, gate211inter7, gate211inter8, gate211inter9, gate211inter10, gate211inter11, gate211inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate278inter0, gate278inter1, gate278inter2, gate278inter3, gate278inter4, gate278inter5, gate278inter6, gate278inter7, gate278inter8, gate278inter9, gate278inter10, gate278inter11, gate278inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate82inter0, gate82inter1, gate82inter2, gate82inter3, gate82inter4, gate82inter5, gate82inter6, gate82inter7, gate82inter8, gate82inter9, gate82inter10, gate82inter11, gate82inter12, gate430inter0, gate430inter1, gate430inter2, gate430inter3, gate430inter4, gate430inter5, gate430inter6, gate430inter7, gate430inter8, gate430inter9, gate430inter10, gate430inter11, gate430inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate122inter0, gate122inter1, gate122inter2, gate122inter3, gate122inter4, gate122inter5, gate122inter6, gate122inter7, gate122inter8, gate122inter9, gate122inter10, gate122inter11, gate122inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate431inter0, gate431inter1, gate431inter2, gate431inter3, gate431inter4, gate431inter5, gate431inter6, gate431inter7, gate431inter8, gate431inter9, gate431inter10, gate431inter11, gate431inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate68inter0, gate68inter1, gate68inter2, gate68inter3, gate68inter4, gate68inter5, gate68inter6, gate68inter7, gate68inter8, gate68inter9, gate68inter10, gate68inter11, gate68inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate80inter0, gate80inter1, gate80inter2, gate80inter3, gate80inter4, gate80inter5, gate80inter6, gate80inter7, gate80inter8, gate80inter9, gate80inter10, gate80inter11, gate80inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate175inter0, gate175inter1, gate175inter2, gate175inter3, gate175inter4, gate175inter5, gate175inter6, gate175inter7, gate175inter8, gate175inter9, gate175inter10, gate175inter11, gate175inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate54inter0, gate54inter1, gate54inter2, gate54inter3, gate54inter4, gate54inter5, gate54inter6, gate54inter7, gate54inter8, gate54inter9, gate54inter10, gate54inter11, gate54inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate458inter0, gate458inter1, gate458inter2, gate458inter3, gate458inter4, gate458inter5, gate458inter6, gate458inter7, gate458inter8, gate458inter9, gate458inter10, gate458inter11, gate458inter12, gate241inter0, gate241inter1, gate241inter2, gate241inter3, gate241inter4, gate241inter5, gate241inter6, gate241inter7, gate241inter8, gate241inter9, gate241inter10, gate241inter11, gate241inter12, gate264inter0, gate264inter1, gate264inter2, gate264inter3, gate264inter4, gate264inter5, gate264inter6, gate264inter7, gate264inter8, gate264inter9, gate264inter10, gate264inter11, gate264inter12, gate427inter0, gate427inter1, gate427inter2, gate427inter3, gate427inter4, gate427inter5, gate427inter6, gate427inter7, gate427inter8, gate427inter9, gate427inter10, gate427inter11, gate427inter12, gate406inter0, gate406inter1, gate406inter2, gate406inter3, gate406inter4, gate406inter5, gate406inter6, gate406inter7, gate406inter8, gate406inter9, gate406inter10, gate406inter11, gate406inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate129inter0, gate129inter1, gate129inter2, gate129inter3, gate129inter4, gate129inter5, gate129inter6, gate129inter7, gate129inter8, gate129inter9, gate129inter10, gate129inter11, gate129inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate437inter0, gate437inter1, gate437inter2, gate437inter3, gate437inter4, gate437inter5, gate437inter6, gate437inter7, gate437inter8, gate437inter9, gate437inter10, gate437inter11, gate437inter12, gate126inter0, gate126inter1, gate126inter2, gate126inter3, gate126inter4, gate126inter5, gate126inter6, gate126inter7, gate126inter8, gate126inter9, gate126inter10, gate126inter11, gate126inter12, gate34inter0, gate34inter1, gate34inter2, gate34inter3, gate34inter4, gate34inter5, gate34inter6, gate34inter7, gate34inter8, gate34inter9, gate34inter10, gate34inter11, gate34inter12, gate491inter0, gate491inter1, gate491inter2, gate491inter3, gate491inter4, gate491inter5, gate491inter6, gate491inter7, gate491inter8, gate491inter9, gate491inter10, gate491inter11, gate491inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate147inter0, gate147inter1, gate147inter2, gate147inter3, gate147inter4, gate147inter5, gate147inter6, gate147inter7, gate147inter8, gate147inter9, gate147inter10, gate147inter11, gate147inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate111inter0, gate111inter1, gate111inter2, gate111inter3, gate111inter4, gate111inter5, gate111inter6, gate111inter7, gate111inter8, gate111inter9, gate111inter10, gate111inter11, gate111inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );

  xor2  gate1275(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate1276(.a(gate10inter0), .b(s_104), .O(gate10inter1));
  and2  gate1277(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate1278(.a(s_104), .O(gate10inter3));
  inv1  gate1279(.a(s_105), .O(gate10inter4));
  nand2 gate1280(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate1281(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate1282(.a(G3), .O(gate10inter7));
  inv1  gate1283(.a(G4), .O(gate10inter8));
  nand2 gate1284(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate1285(.a(s_105), .b(gate10inter3), .O(gate10inter10));
  nor2  gate1286(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate1287(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate1288(.a(gate10inter12), .b(gate10inter1), .O(G269));
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate617(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate618(.a(gate12inter0), .b(s_10), .O(gate12inter1));
  and2  gate619(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate620(.a(s_10), .O(gate12inter3));
  inv1  gate621(.a(s_11), .O(gate12inter4));
  nand2 gate622(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate623(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate624(.a(G7), .O(gate12inter7));
  inv1  gate625(.a(G8), .O(gate12inter8));
  nand2 gate626(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate627(.a(s_11), .b(gate12inter3), .O(gate12inter10));
  nor2  gate628(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate629(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate630(.a(gate12inter12), .b(gate12inter1), .O(G275));

  xor2  gate813(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate814(.a(gate13inter0), .b(s_38), .O(gate13inter1));
  and2  gate815(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate816(.a(s_38), .O(gate13inter3));
  inv1  gate817(.a(s_39), .O(gate13inter4));
  nand2 gate818(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate819(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate820(.a(G9), .O(gate13inter7));
  inv1  gate821(.a(G10), .O(gate13inter8));
  nand2 gate822(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate823(.a(s_39), .b(gate13inter3), .O(gate13inter10));
  nor2  gate824(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate825(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate826(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate827(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate828(.a(gate20inter0), .b(s_40), .O(gate20inter1));
  and2  gate829(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate830(.a(s_40), .O(gate20inter3));
  inv1  gate831(.a(s_41), .O(gate20inter4));
  nand2 gate832(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate833(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate834(.a(G23), .O(gate20inter7));
  inv1  gate835(.a(G24), .O(gate20inter8));
  nand2 gate836(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate837(.a(s_41), .b(gate20inter3), .O(gate20inter10));
  nor2  gate838(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate839(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate840(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );

  xor2  gate1653(.a(G13), .b(G9), .O(gate26inter0));
  nand2 gate1654(.a(gate26inter0), .b(s_158), .O(gate26inter1));
  and2  gate1655(.a(G13), .b(G9), .O(gate26inter2));
  inv1  gate1656(.a(s_158), .O(gate26inter3));
  inv1  gate1657(.a(s_159), .O(gate26inter4));
  nand2 gate1658(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate1659(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate1660(.a(G9), .O(gate26inter7));
  inv1  gate1661(.a(G13), .O(gate26inter8));
  nand2 gate1662(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate1663(.a(s_159), .b(gate26inter3), .O(gate26inter10));
  nor2  gate1664(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate1665(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate1666(.a(gate26inter12), .b(gate26inter1), .O(G317));
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );
nand2 gate31( .a(G4), .b(G8), .O(G332) );
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );

  xor2  gate1541(.a(G29), .b(G25), .O(gate34inter0));
  nand2 gate1542(.a(gate34inter0), .b(s_142), .O(gate34inter1));
  and2  gate1543(.a(G29), .b(G25), .O(gate34inter2));
  inv1  gate1544(.a(s_142), .O(gate34inter3));
  inv1  gate1545(.a(s_143), .O(gate34inter4));
  nand2 gate1546(.a(gate34inter4), .b(gate34inter3), .O(gate34inter5));
  nor2  gate1547(.a(gate34inter5), .b(gate34inter2), .O(gate34inter6));
  inv1  gate1548(.a(G25), .O(gate34inter7));
  inv1  gate1549(.a(G29), .O(gate34inter8));
  nand2 gate1550(.a(gate34inter8), .b(gate34inter7), .O(gate34inter9));
  nand2 gate1551(.a(s_143), .b(gate34inter3), .O(gate34inter10));
  nor2  gate1552(.a(gate34inter10), .b(gate34inter9), .O(gate34inter11));
  nor2  gate1553(.a(gate34inter11), .b(gate34inter6), .O(gate34inter12));
  nand2 gate1554(.a(gate34inter12), .b(gate34inter1), .O(G341));
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate1219(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate1220(.a(gate41inter0), .b(s_96), .O(gate41inter1));
  and2  gate1221(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate1222(.a(s_96), .O(gate41inter3));
  inv1  gate1223(.a(s_97), .O(gate41inter4));
  nand2 gate1224(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate1225(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate1226(.a(G1), .O(gate41inter7));
  inv1  gate1227(.a(G266), .O(gate41inter8));
  nand2 gate1228(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate1229(.a(s_97), .b(gate41inter3), .O(gate41inter10));
  nor2  gate1230(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate1231(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate1232(.a(gate41inter12), .b(gate41inter1), .O(G362));

  xor2  gate1065(.a(G266), .b(G2), .O(gate42inter0));
  nand2 gate1066(.a(gate42inter0), .b(s_74), .O(gate42inter1));
  and2  gate1067(.a(G266), .b(G2), .O(gate42inter2));
  inv1  gate1068(.a(s_74), .O(gate42inter3));
  inv1  gate1069(.a(s_75), .O(gate42inter4));
  nand2 gate1070(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate1071(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate1072(.a(G2), .O(gate42inter7));
  inv1  gate1073(.a(G266), .O(gate42inter8));
  nand2 gate1074(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate1075(.a(s_75), .b(gate42inter3), .O(gate42inter10));
  nor2  gate1076(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate1077(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate1078(.a(gate42inter12), .b(gate42inter1), .O(G363));

  xor2  gate1303(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate1304(.a(gate43inter0), .b(s_108), .O(gate43inter1));
  and2  gate1305(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate1306(.a(s_108), .O(gate43inter3));
  inv1  gate1307(.a(s_109), .O(gate43inter4));
  nand2 gate1308(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate1309(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate1310(.a(G3), .O(gate43inter7));
  inv1  gate1311(.a(G269), .O(gate43inter8));
  nand2 gate1312(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate1313(.a(s_109), .b(gate43inter3), .O(gate43inter10));
  nor2  gate1314(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate1315(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate1316(.a(gate43inter12), .b(gate43inter1), .O(G364));
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate785(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate786(.a(gate46inter0), .b(s_34), .O(gate46inter1));
  and2  gate787(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate788(.a(s_34), .O(gate46inter3));
  inv1  gate789(.a(s_35), .O(gate46inter4));
  nand2 gate790(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate791(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate792(.a(G6), .O(gate46inter7));
  inv1  gate793(.a(G272), .O(gate46inter8));
  nand2 gate794(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate795(.a(s_35), .b(gate46inter3), .O(gate46inter10));
  nor2  gate796(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate797(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate798(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );

  xor2  gate1289(.a(G284), .b(G14), .O(gate54inter0));
  nand2 gate1290(.a(gate54inter0), .b(s_106), .O(gate54inter1));
  and2  gate1291(.a(G284), .b(G14), .O(gate54inter2));
  inv1  gate1292(.a(s_106), .O(gate54inter3));
  inv1  gate1293(.a(s_107), .O(gate54inter4));
  nand2 gate1294(.a(gate54inter4), .b(gate54inter3), .O(gate54inter5));
  nor2  gate1295(.a(gate54inter5), .b(gate54inter2), .O(gate54inter6));
  inv1  gate1296(.a(G14), .O(gate54inter7));
  inv1  gate1297(.a(G284), .O(gate54inter8));
  nand2 gate1298(.a(gate54inter8), .b(gate54inter7), .O(gate54inter9));
  nand2 gate1299(.a(s_107), .b(gate54inter3), .O(gate54inter10));
  nor2  gate1300(.a(gate54inter10), .b(gate54inter9), .O(gate54inter11));
  nor2  gate1301(.a(gate54inter11), .b(gate54inter6), .O(gate54inter12));
  nand2 gate1302(.a(gate54inter12), .b(gate54inter1), .O(G375));
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate1121(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate1122(.a(gate57inter0), .b(s_82), .O(gate57inter1));
  and2  gate1123(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate1124(.a(s_82), .O(gate57inter3));
  inv1  gate1125(.a(s_83), .O(gate57inter4));
  nand2 gate1126(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate1127(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate1128(.a(G17), .O(gate57inter7));
  inv1  gate1129(.a(G290), .O(gate57inter8));
  nand2 gate1130(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate1131(.a(s_83), .b(gate57inter3), .O(gate57inter10));
  nor2  gate1132(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate1133(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate1134(.a(gate57inter12), .b(gate57inter1), .O(G378));
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );
nand2 gate67( .a(G27), .b(G305), .O(G388) );

  xor2  gate1205(.a(G305), .b(G28), .O(gate68inter0));
  nand2 gate1206(.a(gate68inter0), .b(s_94), .O(gate68inter1));
  and2  gate1207(.a(G305), .b(G28), .O(gate68inter2));
  inv1  gate1208(.a(s_94), .O(gate68inter3));
  inv1  gate1209(.a(s_95), .O(gate68inter4));
  nand2 gate1210(.a(gate68inter4), .b(gate68inter3), .O(gate68inter5));
  nor2  gate1211(.a(gate68inter5), .b(gate68inter2), .O(gate68inter6));
  inv1  gate1212(.a(G28), .O(gate68inter7));
  inv1  gate1213(.a(G305), .O(gate68inter8));
  nand2 gate1214(.a(gate68inter8), .b(gate68inter7), .O(gate68inter9));
  nand2 gate1215(.a(s_95), .b(gate68inter3), .O(gate68inter10));
  nor2  gate1216(.a(gate68inter10), .b(gate68inter9), .O(gate68inter11));
  nor2  gate1217(.a(gate68inter11), .b(gate68inter6), .O(gate68inter12));
  nand2 gate1218(.a(gate68inter12), .b(gate68inter1), .O(G389));
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate1009(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate1010(.a(gate71inter0), .b(s_66), .O(gate71inter1));
  and2  gate1011(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate1012(.a(s_66), .O(gate71inter3));
  inv1  gate1013(.a(s_67), .O(gate71inter4));
  nand2 gate1014(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate1015(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate1016(.a(G31), .O(gate71inter7));
  inv1  gate1017(.a(G311), .O(gate71inter8));
  nand2 gate1018(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate1019(.a(s_67), .b(gate71inter3), .O(gate71inter10));
  nor2  gate1020(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate1021(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate1022(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );

  xor2  gate729(.a(G317), .b(G9), .O(gate75inter0));
  nand2 gate730(.a(gate75inter0), .b(s_26), .O(gate75inter1));
  and2  gate731(.a(G317), .b(G9), .O(gate75inter2));
  inv1  gate732(.a(s_26), .O(gate75inter3));
  inv1  gate733(.a(s_27), .O(gate75inter4));
  nand2 gate734(.a(gate75inter4), .b(gate75inter3), .O(gate75inter5));
  nor2  gate735(.a(gate75inter5), .b(gate75inter2), .O(gate75inter6));
  inv1  gate736(.a(G9), .O(gate75inter7));
  inv1  gate737(.a(G317), .O(gate75inter8));
  nand2 gate738(.a(gate75inter8), .b(gate75inter7), .O(gate75inter9));
  nand2 gate739(.a(s_27), .b(gate75inter3), .O(gate75inter10));
  nor2  gate740(.a(gate75inter10), .b(gate75inter9), .O(gate75inter11));
  nor2  gate741(.a(gate75inter11), .b(gate75inter6), .O(gate75inter12));
  nand2 gate742(.a(gate75inter12), .b(gate75inter1), .O(G396));
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );

  xor2  gate1233(.a(G323), .b(G14), .O(gate80inter0));
  nand2 gate1234(.a(gate80inter0), .b(s_98), .O(gate80inter1));
  and2  gate1235(.a(G323), .b(G14), .O(gate80inter2));
  inv1  gate1236(.a(s_98), .O(gate80inter3));
  inv1  gate1237(.a(s_99), .O(gate80inter4));
  nand2 gate1238(.a(gate80inter4), .b(gate80inter3), .O(gate80inter5));
  nor2  gate1239(.a(gate80inter5), .b(gate80inter2), .O(gate80inter6));
  inv1  gate1240(.a(G14), .O(gate80inter7));
  inv1  gate1241(.a(G323), .O(gate80inter8));
  nand2 gate1242(.a(gate80inter8), .b(gate80inter7), .O(gate80inter9));
  nand2 gate1243(.a(s_99), .b(gate80inter3), .O(gate80inter10));
  nor2  gate1244(.a(gate80inter10), .b(gate80inter9), .O(gate80inter11));
  nor2  gate1245(.a(gate80inter11), .b(gate80inter6), .O(gate80inter12));
  nand2 gate1246(.a(gate80inter12), .b(gate80inter1), .O(G401));
nand2 gate81( .a(G3), .b(G326), .O(G402) );

  xor2  gate1079(.a(G326), .b(G7), .O(gate82inter0));
  nand2 gate1080(.a(gate82inter0), .b(s_76), .O(gate82inter1));
  and2  gate1081(.a(G326), .b(G7), .O(gate82inter2));
  inv1  gate1082(.a(s_76), .O(gate82inter3));
  inv1  gate1083(.a(s_77), .O(gate82inter4));
  nand2 gate1084(.a(gate82inter4), .b(gate82inter3), .O(gate82inter5));
  nor2  gate1085(.a(gate82inter5), .b(gate82inter2), .O(gate82inter6));
  inv1  gate1086(.a(G7), .O(gate82inter7));
  inv1  gate1087(.a(G326), .O(gate82inter8));
  nand2 gate1088(.a(gate82inter8), .b(gate82inter7), .O(gate82inter9));
  nand2 gate1089(.a(s_77), .b(gate82inter3), .O(gate82inter10));
  nor2  gate1090(.a(gate82inter10), .b(gate82inter9), .O(gate82inter11));
  nor2  gate1091(.a(gate82inter11), .b(gate82inter6), .O(gate82inter12));
  nand2 gate1092(.a(gate82inter12), .b(gate82inter1), .O(G403));
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate981(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate982(.a(gate94inter0), .b(s_62), .O(gate94inter1));
  and2  gate983(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate984(.a(s_62), .O(gate94inter3));
  inv1  gate985(.a(s_63), .O(gate94inter4));
  nand2 gate986(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate987(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate988(.a(G22), .O(gate94inter7));
  inv1  gate989(.a(G344), .O(gate94inter8));
  nand2 gate990(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate991(.a(s_63), .b(gate94inter3), .O(gate94inter10));
  nor2  gate992(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate993(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate994(.a(gate94inter12), .b(gate94inter1), .O(G415));

  xor2  gate911(.a(G347), .b(G26), .O(gate95inter0));
  nand2 gate912(.a(gate95inter0), .b(s_52), .O(gate95inter1));
  and2  gate913(.a(G347), .b(G26), .O(gate95inter2));
  inv1  gate914(.a(s_52), .O(gate95inter3));
  inv1  gate915(.a(s_53), .O(gate95inter4));
  nand2 gate916(.a(gate95inter4), .b(gate95inter3), .O(gate95inter5));
  nor2  gate917(.a(gate95inter5), .b(gate95inter2), .O(gate95inter6));
  inv1  gate918(.a(G26), .O(gate95inter7));
  inv1  gate919(.a(G347), .O(gate95inter8));
  nand2 gate920(.a(gate95inter8), .b(gate95inter7), .O(gate95inter9));
  nand2 gate921(.a(s_53), .b(gate95inter3), .O(gate95inter10));
  nor2  gate922(.a(gate95inter10), .b(gate95inter9), .O(gate95inter11));
  nor2  gate923(.a(gate95inter11), .b(gate95inter6), .O(gate95inter12));
  nand2 gate924(.a(gate95inter12), .b(gate95inter1), .O(G416));
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate799(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate800(.a(gate98inter0), .b(s_36), .O(gate98inter1));
  and2  gate801(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate802(.a(s_36), .O(gate98inter3));
  inv1  gate803(.a(s_37), .O(gate98inter4));
  nand2 gate804(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate805(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate806(.a(G23), .O(gate98inter7));
  inv1  gate807(.a(G350), .O(gate98inter8));
  nand2 gate808(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate809(.a(s_37), .b(gate98inter3), .O(gate98inter10));
  nor2  gate810(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate811(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate812(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );

  xor2  gate995(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate996(.a(gate105inter0), .b(s_64), .O(gate105inter1));
  and2  gate997(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate998(.a(s_64), .O(gate105inter3));
  inv1  gate999(.a(s_65), .O(gate105inter4));
  nand2 gate1000(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate1001(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate1002(.a(G362), .O(gate105inter7));
  inv1  gate1003(.a(G363), .O(gate105inter8));
  nand2 gate1004(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate1005(.a(s_65), .b(gate105inter3), .O(gate105inter10));
  nor2  gate1006(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate1007(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate1008(.a(gate105inter12), .b(gate105inter1), .O(G426));

  xor2  gate1583(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate1584(.a(gate106inter0), .b(s_148), .O(gate106inter1));
  and2  gate1585(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate1586(.a(s_148), .O(gate106inter3));
  inv1  gate1587(.a(s_149), .O(gate106inter4));
  nand2 gate1588(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate1589(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate1590(.a(G364), .O(gate106inter7));
  inv1  gate1591(.a(G365), .O(gate106inter8));
  nand2 gate1592(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate1593(.a(s_149), .b(gate106inter3), .O(gate106inter10));
  nor2  gate1594(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate1595(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate1596(.a(gate106inter12), .b(gate106inter1), .O(G429));
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );

  xor2  gate883(.a(G373), .b(G372), .O(gate110inter0));
  nand2 gate884(.a(gate110inter0), .b(s_48), .O(gate110inter1));
  and2  gate885(.a(G373), .b(G372), .O(gate110inter2));
  inv1  gate886(.a(s_48), .O(gate110inter3));
  inv1  gate887(.a(s_49), .O(gate110inter4));
  nand2 gate888(.a(gate110inter4), .b(gate110inter3), .O(gate110inter5));
  nor2  gate889(.a(gate110inter5), .b(gate110inter2), .O(gate110inter6));
  inv1  gate890(.a(G372), .O(gate110inter7));
  inv1  gate891(.a(G373), .O(gate110inter8));
  nand2 gate892(.a(gate110inter8), .b(gate110inter7), .O(gate110inter9));
  nand2 gate893(.a(s_49), .b(gate110inter3), .O(gate110inter10));
  nor2  gate894(.a(gate110inter10), .b(gate110inter9), .O(gate110inter11));
  nor2  gate895(.a(gate110inter11), .b(gate110inter6), .O(gate110inter12));
  nand2 gate896(.a(gate110inter12), .b(gate110inter1), .O(G441));

  xor2  gate1667(.a(G375), .b(G374), .O(gate111inter0));
  nand2 gate1668(.a(gate111inter0), .b(s_160), .O(gate111inter1));
  and2  gate1669(.a(G375), .b(G374), .O(gate111inter2));
  inv1  gate1670(.a(s_160), .O(gate111inter3));
  inv1  gate1671(.a(s_161), .O(gate111inter4));
  nand2 gate1672(.a(gate111inter4), .b(gate111inter3), .O(gate111inter5));
  nor2  gate1673(.a(gate111inter5), .b(gate111inter2), .O(gate111inter6));
  inv1  gate1674(.a(G374), .O(gate111inter7));
  inv1  gate1675(.a(G375), .O(gate111inter8));
  nand2 gate1676(.a(gate111inter8), .b(gate111inter7), .O(gate111inter9));
  nand2 gate1677(.a(s_161), .b(gate111inter3), .O(gate111inter10));
  nor2  gate1678(.a(gate111inter10), .b(gate111inter9), .O(gate111inter11));
  nor2  gate1679(.a(gate111inter11), .b(gate111inter6), .O(gate111inter12));
  nand2 gate1680(.a(gate111inter12), .b(gate111inter1), .O(G444));
nand2 gate112( .a(G376), .b(G377), .O(G447) );

  xor2  gate1569(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate1570(.a(gate113inter0), .b(s_146), .O(gate113inter1));
  and2  gate1571(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate1572(.a(s_146), .O(gate113inter3));
  inv1  gate1573(.a(s_147), .O(gate113inter4));
  nand2 gate1574(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate1575(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate1576(.a(G378), .O(gate113inter7));
  inv1  gate1577(.a(G379), .O(gate113inter8));
  nand2 gate1578(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate1579(.a(s_147), .b(gate113inter3), .O(gate113inter10));
  nor2  gate1580(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate1581(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate1582(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );
nand2 gate116( .a(G384), .b(G385), .O(G459) );
nand2 gate117( .a(G386), .b(G387), .O(G462) );

  xor2  gate953(.a(G389), .b(G388), .O(gate118inter0));
  nand2 gate954(.a(gate118inter0), .b(s_58), .O(gate118inter1));
  and2  gate955(.a(G389), .b(G388), .O(gate118inter2));
  inv1  gate956(.a(s_58), .O(gate118inter3));
  inv1  gate957(.a(s_59), .O(gate118inter4));
  nand2 gate958(.a(gate118inter4), .b(gate118inter3), .O(gate118inter5));
  nor2  gate959(.a(gate118inter5), .b(gate118inter2), .O(gate118inter6));
  inv1  gate960(.a(G388), .O(gate118inter7));
  inv1  gate961(.a(G389), .O(gate118inter8));
  nand2 gate962(.a(gate118inter8), .b(gate118inter7), .O(gate118inter9));
  nand2 gate963(.a(s_59), .b(gate118inter3), .O(gate118inter10));
  nor2  gate964(.a(gate118inter10), .b(gate118inter9), .O(gate118inter11));
  nor2  gate965(.a(gate118inter11), .b(gate118inter6), .O(gate118inter12));
  nand2 gate966(.a(gate118inter12), .b(gate118inter1), .O(G465));
nand2 gate119( .a(G390), .b(G391), .O(G468) );

  xor2  gate631(.a(G393), .b(G392), .O(gate120inter0));
  nand2 gate632(.a(gate120inter0), .b(s_12), .O(gate120inter1));
  and2  gate633(.a(G393), .b(G392), .O(gate120inter2));
  inv1  gate634(.a(s_12), .O(gate120inter3));
  inv1  gate635(.a(s_13), .O(gate120inter4));
  nand2 gate636(.a(gate120inter4), .b(gate120inter3), .O(gate120inter5));
  nor2  gate637(.a(gate120inter5), .b(gate120inter2), .O(gate120inter6));
  inv1  gate638(.a(G392), .O(gate120inter7));
  inv1  gate639(.a(G393), .O(gate120inter8));
  nand2 gate640(.a(gate120inter8), .b(gate120inter7), .O(gate120inter9));
  nand2 gate641(.a(s_13), .b(gate120inter3), .O(gate120inter10));
  nor2  gate642(.a(gate120inter10), .b(gate120inter9), .O(gate120inter11));
  nor2  gate643(.a(gate120inter11), .b(gate120inter6), .O(gate120inter12));
  nand2 gate644(.a(gate120inter12), .b(gate120inter1), .O(G471));
nand2 gate121( .a(G394), .b(G395), .O(G474) );

  xor2  gate1135(.a(G397), .b(G396), .O(gate122inter0));
  nand2 gate1136(.a(gate122inter0), .b(s_84), .O(gate122inter1));
  and2  gate1137(.a(G397), .b(G396), .O(gate122inter2));
  inv1  gate1138(.a(s_84), .O(gate122inter3));
  inv1  gate1139(.a(s_85), .O(gate122inter4));
  nand2 gate1140(.a(gate122inter4), .b(gate122inter3), .O(gate122inter5));
  nor2  gate1141(.a(gate122inter5), .b(gate122inter2), .O(gate122inter6));
  inv1  gate1142(.a(G396), .O(gate122inter7));
  inv1  gate1143(.a(G397), .O(gate122inter8));
  nand2 gate1144(.a(gate122inter8), .b(gate122inter7), .O(gate122inter9));
  nand2 gate1145(.a(s_85), .b(gate122inter3), .O(gate122inter10));
  nor2  gate1146(.a(gate122inter10), .b(gate122inter9), .O(gate122inter11));
  nor2  gate1147(.a(gate122inter11), .b(gate122inter6), .O(gate122inter12));
  nand2 gate1148(.a(gate122inter12), .b(gate122inter1), .O(G477));
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );

  xor2  gate1527(.a(G405), .b(G404), .O(gate126inter0));
  nand2 gate1528(.a(gate126inter0), .b(s_140), .O(gate126inter1));
  and2  gate1529(.a(G405), .b(G404), .O(gate126inter2));
  inv1  gate1530(.a(s_140), .O(gate126inter3));
  inv1  gate1531(.a(s_141), .O(gate126inter4));
  nand2 gate1532(.a(gate126inter4), .b(gate126inter3), .O(gate126inter5));
  nor2  gate1533(.a(gate126inter5), .b(gate126inter2), .O(gate126inter6));
  inv1  gate1534(.a(G404), .O(gate126inter7));
  inv1  gate1535(.a(G405), .O(gate126inter8));
  nand2 gate1536(.a(gate126inter8), .b(gate126inter7), .O(gate126inter9));
  nand2 gate1537(.a(s_141), .b(gate126inter3), .O(gate126inter10));
  nor2  gate1538(.a(gate126inter10), .b(gate126inter9), .O(gate126inter11));
  nor2  gate1539(.a(gate126inter11), .b(gate126inter6), .O(gate126inter12));
  nand2 gate1540(.a(gate126inter12), .b(gate126inter1), .O(G489));
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );

  xor2  gate1443(.a(G411), .b(G410), .O(gate129inter0));
  nand2 gate1444(.a(gate129inter0), .b(s_128), .O(gate129inter1));
  and2  gate1445(.a(G411), .b(G410), .O(gate129inter2));
  inv1  gate1446(.a(s_128), .O(gate129inter3));
  inv1  gate1447(.a(s_129), .O(gate129inter4));
  nand2 gate1448(.a(gate129inter4), .b(gate129inter3), .O(gate129inter5));
  nor2  gate1449(.a(gate129inter5), .b(gate129inter2), .O(gate129inter6));
  inv1  gate1450(.a(G410), .O(gate129inter7));
  inv1  gate1451(.a(G411), .O(gate129inter8));
  nand2 gate1452(.a(gate129inter8), .b(gate129inter7), .O(gate129inter9));
  nand2 gate1453(.a(s_129), .b(gate129inter3), .O(gate129inter10));
  nor2  gate1454(.a(gate129inter10), .b(gate129inter9), .O(gate129inter11));
  nor2  gate1455(.a(gate129inter11), .b(gate129inter6), .O(gate129inter12));
  nand2 gate1456(.a(gate129inter12), .b(gate129inter1), .O(G498));
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );
nand2 gate137( .a(G426), .b(G429), .O(G522) );
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate1317(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate1318(.a(gate144inter0), .b(s_110), .O(gate144inter1));
  and2  gate1319(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate1320(.a(s_110), .O(gate144inter3));
  inv1  gate1321(.a(s_111), .O(gate144inter4));
  nand2 gate1322(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate1323(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate1324(.a(G468), .O(gate144inter7));
  inv1  gate1325(.a(G471), .O(gate144inter8));
  nand2 gate1326(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate1327(.a(s_111), .b(gate144inter3), .O(gate144inter10));
  nor2  gate1328(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate1329(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate1330(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );

  xor2  gate743(.a(G483), .b(G480), .O(gate146inter0));
  nand2 gate744(.a(gate146inter0), .b(s_28), .O(gate146inter1));
  and2  gate745(.a(G483), .b(G480), .O(gate146inter2));
  inv1  gate746(.a(s_28), .O(gate146inter3));
  inv1  gate747(.a(s_29), .O(gate146inter4));
  nand2 gate748(.a(gate146inter4), .b(gate146inter3), .O(gate146inter5));
  nor2  gate749(.a(gate146inter5), .b(gate146inter2), .O(gate146inter6));
  inv1  gate750(.a(G480), .O(gate146inter7));
  inv1  gate751(.a(G483), .O(gate146inter8));
  nand2 gate752(.a(gate146inter8), .b(gate146inter7), .O(gate146inter9));
  nand2 gate753(.a(s_29), .b(gate146inter3), .O(gate146inter10));
  nor2  gate754(.a(gate146inter10), .b(gate146inter9), .O(gate146inter11));
  nor2  gate755(.a(gate146inter11), .b(gate146inter6), .O(gate146inter12));
  nand2 gate756(.a(gate146inter12), .b(gate146inter1), .O(G549));

  xor2  gate1597(.a(G489), .b(G486), .O(gate147inter0));
  nand2 gate1598(.a(gate147inter0), .b(s_150), .O(gate147inter1));
  and2  gate1599(.a(G489), .b(G486), .O(gate147inter2));
  inv1  gate1600(.a(s_150), .O(gate147inter3));
  inv1  gate1601(.a(s_151), .O(gate147inter4));
  nand2 gate1602(.a(gate147inter4), .b(gate147inter3), .O(gate147inter5));
  nor2  gate1603(.a(gate147inter5), .b(gate147inter2), .O(gate147inter6));
  inv1  gate1604(.a(G486), .O(gate147inter7));
  inv1  gate1605(.a(G489), .O(gate147inter8));
  nand2 gate1606(.a(gate147inter8), .b(gate147inter7), .O(gate147inter9));
  nand2 gate1607(.a(s_151), .b(gate147inter3), .O(gate147inter10));
  nor2  gate1608(.a(gate147inter10), .b(gate147inter9), .O(gate147inter11));
  nor2  gate1609(.a(gate147inter11), .b(gate147inter6), .O(gate147inter12));
  nand2 gate1610(.a(gate147inter12), .b(gate147inter1), .O(G552));
nand2 gate148( .a(G492), .b(G495), .O(G555) );

  xor2  gate1247(.a(G501), .b(G498), .O(gate149inter0));
  nand2 gate1248(.a(gate149inter0), .b(s_100), .O(gate149inter1));
  and2  gate1249(.a(G501), .b(G498), .O(gate149inter2));
  inv1  gate1250(.a(s_100), .O(gate149inter3));
  inv1  gate1251(.a(s_101), .O(gate149inter4));
  nand2 gate1252(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate1253(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate1254(.a(G498), .O(gate149inter7));
  inv1  gate1255(.a(G501), .O(gate149inter8));
  nand2 gate1256(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate1257(.a(s_101), .b(gate149inter3), .O(gate149inter10));
  nor2  gate1258(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate1259(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate1260(.a(gate149inter12), .b(gate149inter1), .O(G558));
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );

  xor2  gate603(.a(G525), .b(G435), .O(gate156inter0));
  nand2 gate604(.a(gate156inter0), .b(s_8), .O(gate156inter1));
  and2  gate605(.a(G525), .b(G435), .O(gate156inter2));
  inv1  gate606(.a(s_8), .O(gate156inter3));
  inv1  gate607(.a(s_9), .O(gate156inter4));
  nand2 gate608(.a(gate156inter4), .b(gate156inter3), .O(gate156inter5));
  nor2  gate609(.a(gate156inter5), .b(gate156inter2), .O(gate156inter6));
  inv1  gate610(.a(G435), .O(gate156inter7));
  inv1  gate611(.a(G525), .O(gate156inter8));
  nand2 gate612(.a(gate156inter8), .b(gate156inter7), .O(gate156inter9));
  nand2 gate613(.a(s_9), .b(gate156inter3), .O(gate156inter10));
  nor2  gate614(.a(gate156inter10), .b(gate156inter9), .O(gate156inter11));
  nor2  gate615(.a(gate156inter11), .b(gate156inter6), .O(gate156inter12));
  nand2 gate616(.a(gate156inter12), .b(gate156inter1), .O(G573));
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate1401(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate1402(.a(gate160inter0), .b(s_122), .O(gate160inter1));
  and2  gate1403(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate1404(.a(s_122), .O(gate160inter3));
  inv1  gate1405(.a(s_123), .O(gate160inter4));
  nand2 gate1406(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate1407(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate1408(.a(G447), .O(gate160inter7));
  inv1  gate1409(.a(G531), .O(gate160inter8));
  nand2 gate1410(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate1411(.a(s_123), .b(gate160inter3), .O(gate160inter10));
  nor2  gate1412(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate1413(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate1414(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate701(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate702(.a(gate162inter0), .b(s_22), .O(gate162inter1));
  and2  gate703(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate704(.a(s_22), .O(gate162inter3));
  inv1  gate705(.a(s_23), .O(gate162inter4));
  nand2 gate706(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate707(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate708(.a(G453), .O(gate162inter7));
  inv1  gate709(.a(G534), .O(gate162inter8));
  nand2 gate710(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate711(.a(s_23), .b(gate162inter3), .O(gate162inter10));
  nor2  gate712(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate713(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate714(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );

  xor2  gate1261(.a(G555), .b(G492), .O(gate175inter0));
  nand2 gate1262(.a(gate175inter0), .b(s_102), .O(gate175inter1));
  and2  gate1263(.a(G555), .b(G492), .O(gate175inter2));
  inv1  gate1264(.a(s_102), .O(gate175inter3));
  inv1  gate1265(.a(s_103), .O(gate175inter4));
  nand2 gate1266(.a(gate175inter4), .b(gate175inter3), .O(gate175inter5));
  nor2  gate1267(.a(gate175inter5), .b(gate175inter2), .O(gate175inter6));
  inv1  gate1268(.a(G492), .O(gate175inter7));
  inv1  gate1269(.a(G555), .O(gate175inter8));
  nand2 gate1270(.a(gate175inter8), .b(gate175inter7), .O(gate175inter9));
  nand2 gate1271(.a(s_103), .b(gate175inter3), .O(gate175inter10));
  nor2  gate1272(.a(gate175inter10), .b(gate175inter9), .O(gate175inter11));
  nor2  gate1273(.a(gate175inter11), .b(gate175inter6), .O(gate175inter12));
  nand2 gate1274(.a(gate175inter12), .b(gate175inter1), .O(G592));
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );

  xor2  gate757(.a(G585), .b(G584), .O(gate192inter0));
  nand2 gate758(.a(gate192inter0), .b(s_30), .O(gate192inter1));
  and2  gate759(.a(G585), .b(G584), .O(gate192inter2));
  inv1  gate760(.a(s_30), .O(gate192inter3));
  inv1  gate761(.a(s_31), .O(gate192inter4));
  nand2 gate762(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate763(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate764(.a(G584), .O(gate192inter7));
  inv1  gate765(.a(G585), .O(gate192inter8));
  nand2 gate766(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate767(.a(s_31), .b(gate192inter3), .O(gate192inter10));
  nor2  gate768(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate769(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate770(.a(gate192inter12), .b(gate192inter1), .O(G637));
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate897(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate898(.a(gate198inter0), .b(s_50), .O(gate198inter1));
  and2  gate899(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate900(.a(s_50), .O(gate198inter3));
  inv1  gate901(.a(s_51), .O(gate198inter4));
  nand2 gate902(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate903(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate904(.a(G596), .O(gate198inter7));
  inv1  gate905(.a(G597), .O(gate198inter8));
  nand2 gate906(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate907(.a(s_51), .b(gate198inter3), .O(gate198inter10));
  nor2  gate908(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate909(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate910(.a(gate198inter12), .b(gate198inter1), .O(G657));
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );

  xor2  gate1457(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate1458(.a(gate202inter0), .b(s_130), .O(gate202inter1));
  and2  gate1459(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate1460(.a(s_130), .O(gate202inter3));
  inv1  gate1461(.a(s_131), .O(gate202inter4));
  nand2 gate1462(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate1463(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate1464(.a(G612), .O(gate202inter7));
  inv1  gate1465(.a(G617), .O(gate202inter8));
  nand2 gate1466(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate1467(.a(s_131), .b(gate202inter3), .O(gate202inter10));
  nor2  gate1468(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate1469(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate1470(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );

  xor2  gate841(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate842(.a(gate204inter0), .b(s_42), .O(gate204inter1));
  and2  gate843(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate844(.a(s_42), .O(gate204inter3));
  inv1  gate845(.a(s_43), .O(gate204inter4));
  nand2 gate846(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate847(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate848(.a(G607), .O(gate204inter7));
  inv1  gate849(.a(G617), .O(gate204inter8));
  nand2 gate850(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate851(.a(s_43), .b(gate204inter3), .O(gate204inter10));
  nor2  gate852(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate853(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate854(.a(gate204inter12), .b(gate204inter1), .O(G675));
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );

  xor2  gate1107(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate1108(.a(gate210inter0), .b(s_80), .O(gate210inter1));
  and2  gate1109(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate1110(.a(s_80), .O(gate210inter3));
  inv1  gate1111(.a(s_81), .O(gate210inter4));
  nand2 gate1112(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate1113(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate1114(.a(G607), .O(gate210inter7));
  inv1  gate1115(.a(G666), .O(gate210inter8));
  nand2 gate1116(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate1117(.a(s_81), .b(gate210inter3), .O(gate210inter10));
  nor2  gate1118(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate1119(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate1120(.a(gate210inter12), .b(gate210inter1), .O(G691));

  xor2  gate1023(.a(G669), .b(G612), .O(gate211inter0));
  nand2 gate1024(.a(gate211inter0), .b(s_68), .O(gate211inter1));
  and2  gate1025(.a(G669), .b(G612), .O(gate211inter2));
  inv1  gate1026(.a(s_68), .O(gate211inter3));
  inv1  gate1027(.a(s_69), .O(gate211inter4));
  nand2 gate1028(.a(gate211inter4), .b(gate211inter3), .O(gate211inter5));
  nor2  gate1029(.a(gate211inter5), .b(gate211inter2), .O(gate211inter6));
  inv1  gate1030(.a(G612), .O(gate211inter7));
  inv1  gate1031(.a(G669), .O(gate211inter8));
  nand2 gate1032(.a(gate211inter8), .b(gate211inter7), .O(gate211inter9));
  nand2 gate1033(.a(s_69), .b(gate211inter3), .O(gate211inter10));
  nor2  gate1034(.a(gate211inter10), .b(gate211inter9), .O(gate211inter11));
  nor2  gate1035(.a(gate211inter11), .b(gate211inter6), .O(gate211inter12));
  nand2 gate1036(.a(gate211inter12), .b(gate211inter1), .O(G692));
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate575(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate576(.a(gate231inter0), .b(s_4), .O(gate231inter1));
  and2  gate577(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate578(.a(s_4), .O(gate231inter3));
  inv1  gate579(.a(s_5), .O(gate231inter4));
  nand2 gate580(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate581(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate582(.a(G702), .O(gate231inter7));
  inv1  gate583(.a(G703), .O(gate231inter8));
  nand2 gate584(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate585(.a(s_5), .b(gate231inter3), .O(gate231inter10));
  nor2  gate586(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate587(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate588(.a(gate231inter12), .b(gate231inter1), .O(G724));
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate1639(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate1640(.a(gate236inter0), .b(s_156), .O(gate236inter1));
  and2  gate1641(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate1642(.a(s_156), .O(gate236inter3));
  inv1  gate1643(.a(s_157), .O(gate236inter4));
  nand2 gate1644(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate1645(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate1646(.a(G251), .O(gate236inter7));
  inv1  gate1647(.a(G727), .O(gate236inter8));
  nand2 gate1648(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate1649(.a(s_157), .b(gate236inter3), .O(gate236inter10));
  nor2  gate1650(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate1651(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate1652(.a(gate236inter12), .b(gate236inter1), .O(G739));
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );

  xor2  gate1345(.a(G730), .b(G242), .O(gate241inter0));
  nand2 gate1346(.a(gate241inter0), .b(s_114), .O(gate241inter1));
  and2  gate1347(.a(G730), .b(G242), .O(gate241inter2));
  inv1  gate1348(.a(s_114), .O(gate241inter3));
  inv1  gate1349(.a(s_115), .O(gate241inter4));
  nand2 gate1350(.a(gate241inter4), .b(gate241inter3), .O(gate241inter5));
  nor2  gate1351(.a(gate241inter5), .b(gate241inter2), .O(gate241inter6));
  inv1  gate1352(.a(G242), .O(gate241inter7));
  inv1  gate1353(.a(G730), .O(gate241inter8));
  nand2 gate1354(.a(gate241inter8), .b(gate241inter7), .O(gate241inter9));
  nand2 gate1355(.a(s_115), .b(gate241inter3), .O(gate241inter10));
  nor2  gate1356(.a(gate241inter10), .b(gate241inter9), .O(gate241inter11));
  nor2  gate1357(.a(gate241inter11), .b(gate241inter6), .O(gate241inter12));
  nand2 gate1358(.a(gate241inter12), .b(gate241inter1), .O(G754));
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );

  xor2  gate561(.a(G742), .b(G254), .O(gate249inter0));
  nand2 gate562(.a(gate249inter0), .b(s_2), .O(gate249inter1));
  and2  gate563(.a(G742), .b(G254), .O(gate249inter2));
  inv1  gate564(.a(s_2), .O(gate249inter3));
  inv1  gate565(.a(s_3), .O(gate249inter4));
  nand2 gate566(.a(gate249inter4), .b(gate249inter3), .O(gate249inter5));
  nor2  gate567(.a(gate249inter5), .b(gate249inter2), .O(gate249inter6));
  inv1  gate568(.a(G254), .O(gate249inter7));
  inv1  gate569(.a(G742), .O(gate249inter8));
  nand2 gate570(.a(gate249inter8), .b(gate249inter7), .O(gate249inter9));
  nand2 gate571(.a(s_3), .b(gate249inter3), .O(gate249inter10));
  nor2  gate572(.a(gate249inter10), .b(gate249inter9), .O(gate249inter11));
  nor2  gate573(.a(gate249inter11), .b(gate249inter6), .O(gate249inter12));
  nand2 gate574(.a(gate249inter12), .b(gate249inter1), .O(G762));
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate1037(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate1038(.a(gate257inter0), .b(s_70), .O(gate257inter1));
  and2  gate1039(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate1040(.a(s_70), .O(gate257inter3));
  inv1  gate1041(.a(s_71), .O(gate257inter4));
  nand2 gate1042(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate1043(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate1044(.a(G754), .O(gate257inter7));
  inv1  gate1045(.a(G755), .O(gate257inter8));
  nand2 gate1046(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate1047(.a(s_71), .b(gate257inter3), .O(gate257inter10));
  nor2  gate1048(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate1049(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate1050(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );

  xor2  gate659(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate660(.a(gate263inter0), .b(s_16), .O(gate263inter1));
  and2  gate661(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate662(.a(s_16), .O(gate263inter3));
  inv1  gate663(.a(s_17), .O(gate263inter4));
  nand2 gate664(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate665(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate666(.a(G766), .O(gate263inter7));
  inv1  gate667(.a(G767), .O(gate263inter8));
  nand2 gate668(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate669(.a(s_17), .b(gate263inter3), .O(gate263inter10));
  nor2  gate670(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate671(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate672(.a(gate263inter12), .b(gate263inter1), .O(G788));

  xor2  gate1359(.a(G769), .b(G768), .O(gate264inter0));
  nand2 gate1360(.a(gate264inter0), .b(s_116), .O(gate264inter1));
  and2  gate1361(.a(G769), .b(G768), .O(gate264inter2));
  inv1  gate1362(.a(s_116), .O(gate264inter3));
  inv1  gate1363(.a(s_117), .O(gate264inter4));
  nand2 gate1364(.a(gate264inter4), .b(gate264inter3), .O(gate264inter5));
  nor2  gate1365(.a(gate264inter5), .b(gate264inter2), .O(gate264inter6));
  inv1  gate1366(.a(G768), .O(gate264inter7));
  inv1  gate1367(.a(G769), .O(gate264inter8));
  nand2 gate1368(.a(gate264inter8), .b(gate264inter7), .O(gate264inter9));
  nand2 gate1369(.a(s_117), .b(gate264inter3), .O(gate264inter10));
  nor2  gate1370(.a(gate264inter10), .b(gate264inter9), .O(gate264inter11));
  nor2  gate1371(.a(gate264inter11), .b(gate264inter6), .O(gate264inter12));
  nand2 gate1372(.a(gate264inter12), .b(gate264inter1), .O(G791));
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate925(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate926(.a(gate272inter0), .b(s_54), .O(gate272inter1));
  and2  gate927(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate928(.a(s_54), .O(gate272inter3));
  inv1  gate929(.a(s_55), .O(gate272inter4));
  nand2 gate930(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate931(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate932(.a(G663), .O(gate272inter7));
  inv1  gate933(.a(G791), .O(gate272inter8));
  nand2 gate934(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate935(.a(s_55), .b(gate272inter3), .O(gate272inter10));
  nor2  gate936(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate937(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate938(.a(gate272inter12), .b(gate272inter1), .O(G815));

  xor2  gate1611(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate1612(.a(gate273inter0), .b(s_152), .O(gate273inter1));
  and2  gate1613(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate1614(.a(s_152), .O(gate273inter3));
  inv1  gate1615(.a(s_153), .O(gate273inter4));
  nand2 gate1616(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate1617(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate1618(.a(G642), .O(gate273inter7));
  inv1  gate1619(.a(G794), .O(gate273inter8));
  nand2 gate1620(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate1621(.a(s_153), .b(gate273inter3), .O(gate273inter10));
  nor2  gate1622(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate1623(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate1624(.a(gate273inter12), .b(gate273inter1), .O(G818));
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );

  xor2  gate1051(.a(G800), .b(G776), .O(gate278inter0));
  nand2 gate1052(.a(gate278inter0), .b(s_72), .O(gate278inter1));
  and2  gate1053(.a(G800), .b(G776), .O(gate278inter2));
  inv1  gate1054(.a(s_72), .O(gate278inter3));
  inv1  gate1055(.a(s_73), .O(gate278inter4));
  nand2 gate1056(.a(gate278inter4), .b(gate278inter3), .O(gate278inter5));
  nor2  gate1057(.a(gate278inter5), .b(gate278inter2), .O(gate278inter6));
  inv1  gate1058(.a(G776), .O(gate278inter7));
  inv1  gate1059(.a(G800), .O(gate278inter8));
  nand2 gate1060(.a(gate278inter8), .b(gate278inter7), .O(gate278inter9));
  nand2 gate1061(.a(s_73), .b(gate278inter3), .O(gate278inter10));
  nor2  gate1062(.a(gate278inter10), .b(gate278inter9), .O(gate278inter11));
  nor2  gate1063(.a(gate278inter11), .b(gate278inter6), .O(gate278inter12));
  nand2 gate1064(.a(gate278inter12), .b(gate278inter1), .O(G823));
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate1485(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate1486(.a(gate287inter0), .b(s_134), .O(gate287inter1));
  and2  gate1487(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate1488(.a(s_134), .O(gate287inter3));
  inv1  gate1489(.a(s_135), .O(gate287inter4));
  nand2 gate1490(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate1491(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate1492(.a(G663), .O(gate287inter7));
  inv1  gate1493(.a(G815), .O(gate287inter8));
  nand2 gate1494(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate1495(.a(s_135), .b(gate287inter3), .O(gate287inter10));
  nor2  gate1496(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate1497(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate1498(.a(gate287inter12), .b(gate287inter1), .O(G832));

  xor2  gate589(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate590(.a(gate288inter0), .b(s_6), .O(gate288inter1));
  and2  gate591(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate592(.a(s_6), .O(gate288inter3));
  inv1  gate593(.a(s_7), .O(gate288inter4));
  nand2 gate594(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate595(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate596(.a(G791), .O(gate288inter7));
  inv1  gate597(.a(G815), .O(gate288inter8));
  nand2 gate598(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate599(.a(s_7), .b(gate288inter3), .O(gate288inter10));
  nor2  gate600(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate601(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate602(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate939(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate940(.a(gate292inter0), .b(s_56), .O(gate292inter1));
  and2  gate941(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate942(.a(s_56), .O(gate292inter3));
  inv1  gate943(.a(s_57), .O(gate292inter4));
  nand2 gate944(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate945(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate946(.a(G824), .O(gate292inter7));
  inv1  gate947(.a(G825), .O(gate292inter8));
  nand2 gate948(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate949(.a(s_57), .b(gate292inter3), .O(gate292inter10));
  nor2  gate950(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate951(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate952(.a(gate292inter12), .b(gate292inter1), .O(G873));
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate715(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate716(.a(gate295inter0), .b(s_24), .O(gate295inter1));
  and2  gate717(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate718(.a(s_24), .O(gate295inter3));
  inv1  gate719(.a(s_25), .O(gate295inter4));
  nand2 gate720(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate721(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate722(.a(G830), .O(gate295inter7));
  inv1  gate723(.a(G831), .O(gate295inter8));
  nand2 gate724(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate725(.a(s_25), .b(gate295inter3), .O(gate295inter10));
  nor2  gate726(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate727(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate728(.a(gate295inter12), .b(gate295inter1), .O(G912));
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate1625(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate1626(.a(gate390inter0), .b(s_154), .O(gate390inter1));
  and2  gate1627(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate1628(.a(s_154), .O(gate390inter3));
  inv1  gate1629(.a(s_155), .O(gate390inter4));
  nand2 gate1630(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate1631(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate1632(.a(G4), .O(gate390inter7));
  inv1  gate1633(.a(G1045), .O(gate390inter8));
  nand2 gate1634(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate1635(.a(s_155), .b(gate390inter3), .O(gate390inter10));
  nor2  gate1636(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate1637(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate1638(.a(gate390inter12), .b(gate390inter1), .O(G1141));
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );

  xor2  gate1499(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate1500(.a(gate404inter0), .b(s_136), .O(gate404inter1));
  and2  gate1501(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate1502(.a(s_136), .O(gate404inter3));
  inv1  gate1503(.a(s_137), .O(gate404inter4));
  nand2 gate1504(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate1505(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate1506(.a(G18), .O(gate404inter7));
  inv1  gate1507(.a(G1087), .O(gate404inter8));
  nand2 gate1508(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate1509(.a(s_137), .b(gate404inter3), .O(gate404inter10));
  nor2  gate1510(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate1511(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate1512(.a(gate404inter12), .b(gate404inter1), .O(G1183));
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );

  xor2  gate1387(.a(G1093), .b(G20), .O(gate406inter0));
  nand2 gate1388(.a(gate406inter0), .b(s_120), .O(gate406inter1));
  and2  gate1389(.a(G1093), .b(G20), .O(gate406inter2));
  inv1  gate1390(.a(s_120), .O(gate406inter3));
  inv1  gate1391(.a(s_121), .O(gate406inter4));
  nand2 gate1392(.a(gate406inter4), .b(gate406inter3), .O(gate406inter5));
  nor2  gate1393(.a(gate406inter5), .b(gate406inter2), .O(gate406inter6));
  inv1  gate1394(.a(G20), .O(gate406inter7));
  inv1  gate1395(.a(G1093), .O(gate406inter8));
  nand2 gate1396(.a(gate406inter8), .b(gate406inter7), .O(gate406inter9));
  nand2 gate1397(.a(s_121), .b(gate406inter3), .O(gate406inter10));
  nor2  gate1398(.a(gate406inter10), .b(gate406inter9), .O(gate406inter11));
  nor2  gate1399(.a(gate406inter11), .b(gate406inter6), .O(gate406inter12));
  nand2 gate1400(.a(gate406inter12), .b(gate406inter1), .O(G1189));
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );

  xor2  gate855(.a(G1108), .b(G25), .O(gate411inter0));
  nand2 gate856(.a(gate411inter0), .b(s_44), .O(gate411inter1));
  and2  gate857(.a(G1108), .b(G25), .O(gate411inter2));
  inv1  gate858(.a(s_44), .O(gate411inter3));
  inv1  gate859(.a(s_45), .O(gate411inter4));
  nand2 gate860(.a(gate411inter4), .b(gate411inter3), .O(gate411inter5));
  nor2  gate861(.a(gate411inter5), .b(gate411inter2), .O(gate411inter6));
  inv1  gate862(.a(G25), .O(gate411inter7));
  inv1  gate863(.a(G1108), .O(gate411inter8));
  nand2 gate864(.a(gate411inter8), .b(gate411inter7), .O(gate411inter9));
  nand2 gate865(.a(s_45), .b(gate411inter3), .O(gate411inter10));
  nor2  gate866(.a(gate411inter10), .b(gate411inter9), .O(gate411inter11));
  nor2  gate867(.a(gate411inter11), .b(gate411inter6), .O(gate411inter12));
  nand2 gate868(.a(gate411inter12), .b(gate411inter1), .O(G1204));
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );

  xor2  gate687(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate688(.a(gate425inter0), .b(s_20), .O(gate425inter1));
  and2  gate689(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate690(.a(s_20), .O(gate425inter3));
  inv1  gate691(.a(s_21), .O(gate425inter4));
  nand2 gate692(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate693(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate694(.a(G4), .O(gate425inter7));
  inv1  gate695(.a(G1141), .O(gate425inter8));
  nand2 gate696(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate697(.a(s_21), .b(gate425inter3), .O(gate425inter10));
  nor2  gate698(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate699(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate700(.a(gate425inter12), .b(gate425inter1), .O(G1234));

  xor2  gate1191(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate1192(.a(gate426inter0), .b(s_92), .O(gate426inter1));
  and2  gate1193(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate1194(.a(s_92), .O(gate426inter3));
  inv1  gate1195(.a(s_93), .O(gate426inter4));
  nand2 gate1196(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate1197(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate1198(.a(G1045), .O(gate426inter7));
  inv1  gate1199(.a(G1141), .O(gate426inter8));
  nand2 gate1200(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate1201(.a(s_93), .b(gate426inter3), .O(gate426inter10));
  nor2  gate1202(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate1203(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate1204(.a(gate426inter12), .b(gate426inter1), .O(G1235));

  xor2  gate1373(.a(G1144), .b(G5), .O(gate427inter0));
  nand2 gate1374(.a(gate427inter0), .b(s_118), .O(gate427inter1));
  and2  gate1375(.a(G1144), .b(G5), .O(gate427inter2));
  inv1  gate1376(.a(s_118), .O(gate427inter3));
  inv1  gate1377(.a(s_119), .O(gate427inter4));
  nand2 gate1378(.a(gate427inter4), .b(gate427inter3), .O(gate427inter5));
  nor2  gate1379(.a(gate427inter5), .b(gate427inter2), .O(gate427inter6));
  inv1  gate1380(.a(G5), .O(gate427inter7));
  inv1  gate1381(.a(G1144), .O(gate427inter8));
  nand2 gate1382(.a(gate427inter8), .b(gate427inter7), .O(gate427inter9));
  nand2 gate1383(.a(s_119), .b(gate427inter3), .O(gate427inter10));
  nor2  gate1384(.a(gate427inter10), .b(gate427inter9), .O(gate427inter11));
  nor2  gate1385(.a(gate427inter11), .b(gate427inter6), .O(gate427inter12));
  nand2 gate1386(.a(gate427inter12), .b(gate427inter1), .O(G1236));
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );

  xor2  gate1093(.a(G1147), .b(G1051), .O(gate430inter0));
  nand2 gate1094(.a(gate430inter0), .b(s_78), .O(gate430inter1));
  and2  gate1095(.a(G1147), .b(G1051), .O(gate430inter2));
  inv1  gate1096(.a(s_78), .O(gate430inter3));
  inv1  gate1097(.a(s_79), .O(gate430inter4));
  nand2 gate1098(.a(gate430inter4), .b(gate430inter3), .O(gate430inter5));
  nor2  gate1099(.a(gate430inter5), .b(gate430inter2), .O(gate430inter6));
  inv1  gate1100(.a(G1051), .O(gate430inter7));
  inv1  gate1101(.a(G1147), .O(gate430inter8));
  nand2 gate1102(.a(gate430inter8), .b(gate430inter7), .O(gate430inter9));
  nand2 gate1103(.a(s_79), .b(gate430inter3), .O(gate430inter10));
  nor2  gate1104(.a(gate430inter10), .b(gate430inter9), .O(gate430inter11));
  nor2  gate1105(.a(gate430inter11), .b(gate430inter6), .O(gate430inter12));
  nand2 gate1106(.a(gate430inter12), .b(gate430inter1), .O(G1239));

  xor2  gate1163(.a(G1150), .b(G7), .O(gate431inter0));
  nand2 gate1164(.a(gate431inter0), .b(s_88), .O(gate431inter1));
  and2  gate1165(.a(G1150), .b(G7), .O(gate431inter2));
  inv1  gate1166(.a(s_88), .O(gate431inter3));
  inv1  gate1167(.a(s_89), .O(gate431inter4));
  nand2 gate1168(.a(gate431inter4), .b(gate431inter3), .O(gate431inter5));
  nor2  gate1169(.a(gate431inter5), .b(gate431inter2), .O(gate431inter6));
  inv1  gate1170(.a(G7), .O(gate431inter7));
  inv1  gate1171(.a(G1150), .O(gate431inter8));
  nand2 gate1172(.a(gate431inter8), .b(gate431inter7), .O(gate431inter9));
  nand2 gate1173(.a(s_89), .b(gate431inter3), .O(gate431inter10));
  nor2  gate1174(.a(gate431inter10), .b(gate431inter9), .O(gate431inter11));
  nor2  gate1175(.a(gate431inter11), .b(gate431inter6), .O(gate431inter12));
  nand2 gate1176(.a(gate431inter12), .b(gate431inter1), .O(G1240));
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );

  xor2  gate1513(.a(G1159), .b(G10), .O(gate437inter0));
  nand2 gate1514(.a(gate437inter0), .b(s_138), .O(gate437inter1));
  and2  gate1515(.a(G1159), .b(G10), .O(gate437inter2));
  inv1  gate1516(.a(s_138), .O(gate437inter3));
  inv1  gate1517(.a(s_139), .O(gate437inter4));
  nand2 gate1518(.a(gate437inter4), .b(gate437inter3), .O(gate437inter5));
  nor2  gate1519(.a(gate437inter5), .b(gate437inter2), .O(gate437inter6));
  inv1  gate1520(.a(G10), .O(gate437inter7));
  inv1  gate1521(.a(G1159), .O(gate437inter8));
  nand2 gate1522(.a(gate437inter8), .b(gate437inter7), .O(gate437inter9));
  nand2 gate1523(.a(s_139), .b(gate437inter3), .O(gate437inter10));
  nor2  gate1524(.a(gate437inter10), .b(gate437inter9), .O(gate437inter11));
  nor2  gate1525(.a(gate437inter11), .b(gate437inter6), .O(gate437inter12));
  nand2 gate1526(.a(gate437inter12), .b(gate437inter1), .O(G1246));

  xor2  gate645(.a(G1159), .b(G1063), .O(gate438inter0));
  nand2 gate646(.a(gate438inter0), .b(s_14), .O(gate438inter1));
  and2  gate647(.a(G1159), .b(G1063), .O(gate438inter2));
  inv1  gate648(.a(s_14), .O(gate438inter3));
  inv1  gate649(.a(s_15), .O(gate438inter4));
  nand2 gate650(.a(gate438inter4), .b(gate438inter3), .O(gate438inter5));
  nor2  gate651(.a(gate438inter5), .b(gate438inter2), .O(gate438inter6));
  inv1  gate652(.a(G1063), .O(gate438inter7));
  inv1  gate653(.a(G1159), .O(gate438inter8));
  nand2 gate654(.a(gate438inter8), .b(gate438inter7), .O(gate438inter9));
  nand2 gate655(.a(s_15), .b(gate438inter3), .O(gate438inter10));
  nor2  gate656(.a(gate438inter10), .b(gate438inter9), .O(gate438inter11));
  nor2  gate657(.a(gate438inter11), .b(gate438inter6), .O(gate438inter12));
  nand2 gate658(.a(gate438inter12), .b(gate438inter1), .O(G1247));

  xor2  gate1429(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate1430(.a(gate439inter0), .b(s_126), .O(gate439inter1));
  and2  gate1431(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate1432(.a(s_126), .O(gate439inter3));
  inv1  gate1433(.a(s_127), .O(gate439inter4));
  nand2 gate1434(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate1435(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate1436(.a(G11), .O(gate439inter7));
  inv1  gate1437(.a(G1162), .O(gate439inter8));
  nand2 gate1438(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate1439(.a(s_127), .b(gate439inter3), .O(gate439inter10));
  nor2  gate1440(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate1441(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate1442(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );

  xor2  gate869(.a(G1168), .b(G1072), .O(gate444inter0));
  nand2 gate870(.a(gate444inter0), .b(s_46), .O(gate444inter1));
  and2  gate871(.a(G1168), .b(G1072), .O(gate444inter2));
  inv1  gate872(.a(s_46), .O(gate444inter3));
  inv1  gate873(.a(s_47), .O(gate444inter4));
  nand2 gate874(.a(gate444inter4), .b(gate444inter3), .O(gate444inter5));
  nor2  gate875(.a(gate444inter5), .b(gate444inter2), .O(gate444inter6));
  inv1  gate876(.a(G1072), .O(gate444inter7));
  inv1  gate877(.a(G1168), .O(gate444inter8));
  nand2 gate878(.a(gate444inter8), .b(gate444inter7), .O(gate444inter9));
  nand2 gate879(.a(s_47), .b(gate444inter3), .O(gate444inter10));
  nor2  gate880(.a(gate444inter10), .b(gate444inter9), .O(gate444inter11));
  nor2  gate881(.a(gate444inter11), .b(gate444inter6), .O(gate444inter12));
  nand2 gate882(.a(gate444inter12), .b(gate444inter1), .O(G1253));
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );

  xor2  gate1331(.a(G1189), .b(G1093), .O(gate458inter0));
  nand2 gate1332(.a(gate458inter0), .b(s_112), .O(gate458inter1));
  and2  gate1333(.a(G1189), .b(G1093), .O(gate458inter2));
  inv1  gate1334(.a(s_112), .O(gate458inter3));
  inv1  gate1335(.a(s_113), .O(gate458inter4));
  nand2 gate1336(.a(gate458inter4), .b(gate458inter3), .O(gate458inter5));
  nor2  gate1337(.a(gate458inter5), .b(gate458inter2), .O(gate458inter6));
  inv1  gate1338(.a(G1093), .O(gate458inter7));
  inv1  gate1339(.a(G1189), .O(gate458inter8));
  nand2 gate1340(.a(gate458inter8), .b(gate458inter7), .O(gate458inter9));
  nand2 gate1341(.a(s_113), .b(gate458inter3), .O(gate458inter10));
  nor2  gate1342(.a(gate458inter10), .b(gate458inter9), .O(gate458inter11));
  nor2  gate1343(.a(gate458inter11), .b(gate458inter6), .O(gate458inter12));
  nand2 gate1344(.a(gate458inter12), .b(gate458inter1), .O(G1267));
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate1177(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate1178(.a(gate460inter0), .b(s_90), .O(gate460inter1));
  and2  gate1179(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate1180(.a(s_90), .O(gate460inter3));
  inv1  gate1181(.a(s_91), .O(gate460inter4));
  nand2 gate1182(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate1183(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate1184(.a(G1096), .O(gate460inter7));
  inv1  gate1185(.a(G1192), .O(gate460inter8));
  nand2 gate1186(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate1187(.a(s_91), .b(gate460inter3), .O(gate460inter10));
  nor2  gate1188(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate1189(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate1190(.a(gate460inter12), .b(gate460inter1), .O(G1269));

  xor2  gate967(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate968(.a(gate461inter0), .b(s_60), .O(gate461inter1));
  and2  gate969(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate970(.a(s_60), .O(gate461inter3));
  inv1  gate971(.a(s_61), .O(gate461inter4));
  nand2 gate972(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate973(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate974(.a(G22), .O(gate461inter7));
  inv1  gate975(.a(G1195), .O(gate461inter8));
  nand2 gate976(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate977(.a(s_61), .b(gate461inter3), .O(gate461inter10));
  nor2  gate978(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate979(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate980(.a(gate461inter12), .b(gate461inter1), .O(G1270));

  xor2  gate771(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate772(.a(gate462inter0), .b(s_32), .O(gate462inter1));
  and2  gate773(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate774(.a(s_32), .O(gate462inter3));
  inv1  gate775(.a(s_33), .O(gate462inter4));
  nand2 gate776(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate777(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate778(.a(G1099), .O(gate462inter7));
  inv1  gate779(.a(G1195), .O(gate462inter8));
  nand2 gate780(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate781(.a(s_33), .b(gate462inter3), .O(gate462inter10));
  nor2  gate782(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate783(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate784(.a(gate462inter12), .b(gate462inter1), .O(G1271));
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );

  xor2  gate1415(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate1416(.a(gate464inter0), .b(s_124), .O(gate464inter1));
  and2  gate1417(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate1418(.a(s_124), .O(gate464inter3));
  inv1  gate1419(.a(s_125), .O(gate464inter4));
  nand2 gate1420(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate1421(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate1422(.a(G1102), .O(gate464inter7));
  inv1  gate1423(.a(G1198), .O(gate464inter8));
  nand2 gate1424(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate1425(.a(s_125), .b(gate464inter3), .O(gate464inter10));
  nor2  gate1426(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate1427(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate1428(.a(gate464inter12), .b(gate464inter1), .O(G1273));

  xor2  gate673(.a(G1201), .b(G24), .O(gate465inter0));
  nand2 gate674(.a(gate465inter0), .b(s_18), .O(gate465inter1));
  and2  gate675(.a(G1201), .b(G24), .O(gate465inter2));
  inv1  gate676(.a(s_18), .O(gate465inter3));
  inv1  gate677(.a(s_19), .O(gate465inter4));
  nand2 gate678(.a(gate465inter4), .b(gate465inter3), .O(gate465inter5));
  nor2  gate679(.a(gate465inter5), .b(gate465inter2), .O(gate465inter6));
  inv1  gate680(.a(G24), .O(gate465inter7));
  inv1  gate681(.a(G1201), .O(gate465inter8));
  nand2 gate682(.a(gate465inter8), .b(gate465inter7), .O(gate465inter9));
  nand2 gate683(.a(s_19), .b(gate465inter3), .O(gate465inter10));
  nor2  gate684(.a(gate465inter10), .b(gate465inter9), .O(gate465inter11));
  nor2  gate685(.a(gate465inter11), .b(gate465inter6), .O(gate465inter12));
  nand2 gate686(.a(gate465inter12), .b(gate465inter1), .O(G1274));
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate1471(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate1472(.a(gate480inter0), .b(s_132), .O(gate480inter1));
  and2  gate1473(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate1474(.a(s_132), .O(gate480inter3));
  inv1  gate1475(.a(s_133), .O(gate480inter4));
  nand2 gate1476(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate1477(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate1478(.a(G1126), .O(gate480inter7));
  inv1  gate1479(.a(G1222), .O(gate480inter8));
  nand2 gate1480(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate1481(.a(s_133), .b(gate480inter3), .O(gate480inter10));
  nor2  gate1482(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate1483(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate1484(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );

  xor2  gate1555(.a(G1245), .b(G1244), .O(gate491inter0));
  nand2 gate1556(.a(gate491inter0), .b(s_144), .O(gate491inter1));
  and2  gate1557(.a(G1245), .b(G1244), .O(gate491inter2));
  inv1  gate1558(.a(s_144), .O(gate491inter3));
  inv1  gate1559(.a(s_145), .O(gate491inter4));
  nand2 gate1560(.a(gate491inter4), .b(gate491inter3), .O(gate491inter5));
  nor2  gate1561(.a(gate491inter5), .b(gate491inter2), .O(gate491inter6));
  inv1  gate1562(.a(G1244), .O(gate491inter7));
  inv1  gate1563(.a(G1245), .O(gate491inter8));
  nand2 gate1564(.a(gate491inter8), .b(gate491inter7), .O(gate491inter9));
  nand2 gate1565(.a(s_145), .b(gate491inter3), .O(gate491inter10));
  nor2  gate1566(.a(gate491inter10), .b(gate491inter9), .O(gate491inter11));
  nor2  gate1567(.a(gate491inter11), .b(gate491inter6), .O(gate491inter12));
  nand2 gate1568(.a(gate491inter12), .b(gate491inter1), .O(G1300));
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );

  xor2  gate547(.a(G1253), .b(G1252), .O(gate495inter0));
  nand2 gate548(.a(gate495inter0), .b(s_0), .O(gate495inter1));
  and2  gate549(.a(G1253), .b(G1252), .O(gate495inter2));
  inv1  gate550(.a(s_0), .O(gate495inter3));
  inv1  gate551(.a(s_1), .O(gate495inter4));
  nand2 gate552(.a(gate495inter4), .b(gate495inter3), .O(gate495inter5));
  nor2  gate553(.a(gate495inter5), .b(gate495inter2), .O(gate495inter6));
  inv1  gate554(.a(G1252), .O(gate495inter7));
  inv1  gate555(.a(G1253), .O(gate495inter8));
  nand2 gate556(.a(gate495inter8), .b(gate495inter7), .O(gate495inter9));
  nand2 gate557(.a(s_1), .b(gate495inter3), .O(gate495inter10));
  nor2  gate558(.a(gate495inter10), .b(gate495inter9), .O(gate495inter11));
  nor2  gate559(.a(gate495inter11), .b(gate495inter6), .O(gate495inter12));
  nand2 gate560(.a(gate495inter12), .b(gate495inter1), .O(G1304));
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate1149(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate1150(.a(gate510inter0), .b(s_86), .O(gate510inter1));
  and2  gate1151(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate1152(.a(s_86), .O(gate510inter3));
  inv1  gate1153(.a(s_87), .O(gate510inter4));
  nand2 gate1154(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate1155(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate1156(.a(G1282), .O(gate510inter7));
  inv1  gate1157(.a(G1283), .O(gate510inter8));
  nand2 gate1158(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate1159(.a(s_87), .b(gate510inter3), .O(gate510inter10));
  nor2  gate1160(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate1161(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate1162(.a(gate510inter12), .b(gate510inter1), .O(G1319));
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule