module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate98inter0, gate98inter1, gate98inter2, gate98inter3, gate98inter4, gate98inter5, gate98inter6, gate98inter7, gate98inter8, gate98inter9, gate98inter10, gate98inter11, gate98inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate12inter0, gate12inter1, gate12inter2, gate12inter3, gate12inter4, gate12inter5, gate12inter6, gate12inter7, gate12inter8, gate12inter9, gate12inter10, gate12inter11, gate12inter12, gate484inter0, gate484inter1, gate484inter2, gate484inter3, gate484inter4, gate484inter5, gate484inter6, gate484inter7, gate484inter8, gate484inter9, gate484inter10, gate484inter11, gate484inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate113inter0, gate113inter1, gate113inter2, gate113inter3, gate113inter4, gate113inter5, gate113inter6, gate113inter7, gate113inter8, gate113inter9, gate113inter10, gate113inter11, gate113inter12, gate479inter0, gate479inter1, gate479inter2, gate479inter3, gate479inter4, gate479inter5, gate479inter6, gate479inter7, gate479inter8, gate479inter9, gate479inter10, gate479inter11, gate479inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate494inter0, gate494inter1, gate494inter2, gate494inter3, gate494inter4, gate494inter5, gate494inter6, gate494inter7, gate494inter8, gate494inter9, gate494inter10, gate494inter11, gate494inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate88inter0, gate88inter1, gate88inter2, gate88inter3, gate88inter4, gate88inter5, gate88inter6, gate88inter7, gate88inter8, gate88inter9, gate88inter10, gate88inter11, gate88inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate229inter0, gate229inter1, gate229inter2, gate229inter3, gate229inter4, gate229inter5, gate229inter6, gate229inter7, gate229inter8, gate229inter9, gate229inter10, gate229inter11, gate229inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate133inter0, gate133inter1, gate133inter2, gate133inter3, gate133inter4, gate133inter5, gate133inter6, gate133inter7, gate133inter8, gate133inter9, gate133inter10, gate133inter11, gate133inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate257inter0, gate257inter1, gate257inter2, gate257inter3, gate257inter4, gate257inter5, gate257inter6, gate257inter7, gate257inter8, gate257inter9, gate257inter10, gate257inter11, gate257inter12, gate154inter0, gate154inter1, gate154inter2, gate154inter3, gate154inter4, gate154inter5, gate154inter6, gate154inter7, gate154inter8, gate154inter9, gate154inter10, gate154inter11, gate154inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate487inter0, gate487inter1, gate487inter2, gate487inter3, gate487inter4, gate487inter5, gate487inter6, gate487inter7, gate487inter8, gate487inter9, gate487inter10, gate487inter11, gate487inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate117inter0, gate117inter1, gate117inter2, gate117inter3, gate117inter4, gate117inter5, gate117inter6, gate117inter7, gate117inter8, gate117inter9, gate117inter10, gate117inter11, gate117inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate94inter0, gate94inter1, gate94inter2, gate94inter3, gate94inter4, gate94inter5, gate94inter6, gate94inter7, gate94inter8, gate94inter9, gate94inter10, gate94inter11, gate94inter12, gate460inter0, gate460inter1, gate460inter2, gate460inter3, gate460inter4, gate460inter5, gate460inter6, gate460inter7, gate460inter8, gate460inter9, gate460inter10, gate460inter11, gate460inter12, gate48inter0, gate48inter1, gate48inter2, gate48inter3, gate48inter4, gate48inter5, gate48inter6, gate48inter7, gate48inter8, gate48inter9, gate48inter10, gate48inter11, gate48inter12, gate488inter0, gate488inter1, gate488inter2, gate488inter3, gate488inter4, gate488inter5, gate488inter6, gate488inter7, gate488inter8, gate488inter9, gate488inter10, gate488inter11, gate488inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate489inter0, gate489inter1, gate489inter2, gate489inter3, gate489inter4, gate489inter5, gate489inter6, gate489inter7, gate489inter8, gate489inter9, gate489inter10, gate489inter11, gate489inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate204inter0, gate204inter1, gate204inter2, gate204inter3, gate204inter4, gate204inter5, gate204inter6, gate204inter7, gate204inter8, gate204inter9, gate204inter10, gate204inter11, gate204inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate41inter0, gate41inter1, gate41inter2, gate41inter3, gate41inter4, gate41inter5, gate41inter6, gate41inter7, gate41inter8, gate41inter9, gate41inter10, gate41inter11, gate41inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );

  xor2  gate603(.a(G8), .b(G7), .O(gate12inter0));
  nand2 gate604(.a(gate12inter0), .b(s_8), .O(gate12inter1));
  and2  gate605(.a(G8), .b(G7), .O(gate12inter2));
  inv1  gate606(.a(s_8), .O(gate12inter3));
  inv1  gate607(.a(s_9), .O(gate12inter4));
  nand2 gate608(.a(gate12inter4), .b(gate12inter3), .O(gate12inter5));
  nor2  gate609(.a(gate12inter5), .b(gate12inter2), .O(gate12inter6));
  inv1  gate610(.a(G7), .O(gate12inter7));
  inv1  gate611(.a(G8), .O(gate12inter8));
  nand2 gate612(.a(gate12inter8), .b(gate12inter7), .O(gate12inter9));
  nand2 gate613(.a(s_9), .b(gate12inter3), .O(gate12inter10));
  nor2  gate614(.a(gate12inter10), .b(gate12inter9), .O(gate12inter11));
  nor2  gate615(.a(gate12inter11), .b(gate12inter6), .O(gate12inter12));
  nand2 gate616(.a(gate12inter12), .b(gate12inter1), .O(G275));

  xor2  gate1121(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate1122(.a(gate13inter0), .b(s_82), .O(gate13inter1));
  and2  gate1123(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate1124(.a(s_82), .O(gate13inter3));
  inv1  gate1125(.a(s_83), .O(gate13inter4));
  nand2 gate1126(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate1127(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate1128(.a(G9), .O(gate13inter7));
  inv1  gate1129(.a(G10), .O(gate13inter8));
  nand2 gate1130(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate1131(.a(s_83), .b(gate13inter3), .O(gate13inter10));
  nor2  gate1132(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate1133(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate1134(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate575(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate576(.a(gate15inter0), .b(s_4), .O(gate15inter1));
  and2  gate577(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate578(.a(s_4), .O(gate15inter3));
  inv1  gate579(.a(s_5), .O(gate15inter4));
  nand2 gate580(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate581(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate582(.a(G13), .O(gate15inter7));
  inv1  gate583(.a(G14), .O(gate15inter8));
  nand2 gate584(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate585(.a(s_5), .b(gate15inter3), .O(gate15inter10));
  nor2  gate586(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate587(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate588(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );
nand2 gate20( .a(G23), .b(G24), .O(G299) );
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate785(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate786(.a(gate31inter0), .b(s_34), .O(gate31inter1));
  and2  gate787(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate788(.a(s_34), .O(gate31inter3));
  inv1  gate789(.a(s_35), .O(gate31inter4));
  nand2 gate790(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate791(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate792(.a(G4), .O(gate31inter7));
  inv1  gate793(.a(G8), .O(gate31inter8));
  nand2 gate794(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate795(.a(s_35), .b(gate31inter3), .O(gate31inter10));
  nor2  gate796(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate797(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate798(.a(gate31inter12), .b(gate31inter1), .O(G332));
nand2 gate32( .a(G12), .b(G16), .O(G335) );
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );

  xor2  gate1163(.a(G266), .b(G1), .O(gate41inter0));
  nand2 gate1164(.a(gate41inter0), .b(s_88), .O(gate41inter1));
  and2  gate1165(.a(G266), .b(G1), .O(gate41inter2));
  inv1  gate1166(.a(s_88), .O(gate41inter3));
  inv1  gate1167(.a(s_89), .O(gate41inter4));
  nand2 gate1168(.a(gate41inter4), .b(gate41inter3), .O(gate41inter5));
  nor2  gate1169(.a(gate41inter5), .b(gate41inter2), .O(gate41inter6));
  inv1  gate1170(.a(G1), .O(gate41inter7));
  inv1  gate1171(.a(G266), .O(gate41inter8));
  nand2 gate1172(.a(gate41inter8), .b(gate41inter7), .O(gate41inter9));
  nand2 gate1173(.a(s_89), .b(gate41inter3), .O(gate41inter10));
  nor2  gate1174(.a(gate41inter10), .b(gate41inter9), .O(gate41inter11));
  nor2  gate1175(.a(gate41inter11), .b(gate41inter6), .O(gate41inter12));
  nand2 gate1176(.a(gate41inter12), .b(gate41inter1), .O(G362));
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate1051(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate1052(.a(gate43inter0), .b(s_72), .O(gate43inter1));
  and2  gate1053(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate1054(.a(s_72), .O(gate43inter3));
  inv1  gate1055(.a(s_73), .O(gate43inter4));
  nand2 gate1056(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate1057(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate1058(.a(G3), .O(gate43inter7));
  inv1  gate1059(.a(G269), .O(gate43inter8));
  nand2 gate1060(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate1061(.a(s_73), .b(gate43inter3), .O(gate43inter10));
  nor2  gate1062(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate1063(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate1064(.a(gate43inter12), .b(gate43inter1), .O(G364));
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );
nand2 gate47( .a(G7), .b(G275), .O(G368) );

  xor2  gate1009(.a(G275), .b(G8), .O(gate48inter0));
  nand2 gate1010(.a(gate48inter0), .b(s_66), .O(gate48inter1));
  and2  gate1011(.a(G275), .b(G8), .O(gate48inter2));
  inv1  gate1012(.a(s_66), .O(gate48inter3));
  inv1  gate1013(.a(s_67), .O(gate48inter4));
  nand2 gate1014(.a(gate48inter4), .b(gate48inter3), .O(gate48inter5));
  nor2  gate1015(.a(gate48inter5), .b(gate48inter2), .O(gate48inter6));
  inv1  gate1016(.a(G8), .O(gate48inter7));
  inv1  gate1017(.a(G275), .O(gate48inter8));
  nand2 gate1018(.a(gate48inter8), .b(gate48inter7), .O(gate48inter9));
  nand2 gate1019(.a(s_67), .b(gate48inter3), .O(gate48inter10));
  nor2  gate1020(.a(gate48inter10), .b(gate48inter9), .O(gate48inter11));
  nor2  gate1021(.a(gate48inter11), .b(gate48inter6), .O(gate48inter12));
  nand2 gate1022(.a(gate48inter12), .b(gate48inter1), .O(G369));
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );
nand2 gate53( .a(G13), .b(G284), .O(G374) );
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate897(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate898(.a(gate67inter0), .b(s_50), .O(gate67inter1));
  and2  gate899(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate900(.a(s_50), .O(gate67inter3));
  inv1  gate901(.a(s_51), .O(gate67inter4));
  nand2 gate902(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate903(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate904(.a(G27), .O(gate67inter7));
  inv1  gate905(.a(G305), .O(gate67inter8));
  nand2 gate906(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate907(.a(s_51), .b(gate67inter3), .O(gate67inter10));
  nor2  gate908(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate909(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate910(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );
nand2 gate71( .a(G31), .b(G311), .O(G392) );
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );
nand2 gate84( .a(G15), .b(G329), .O(G405) );
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );

  xor2  gate771(.a(G335), .b(G16), .O(gate88inter0));
  nand2 gate772(.a(gate88inter0), .b(s_32), .O(gate88inter1));
  and2  gate773(.a(G335), .b(G16), .O(gate88inter2));
  inv1  gate774(.a(s_32), .O(gate88inter3));
  inv1  gate775(.a(s_33), .O(gate88inter4));
  nand2 gate776(.a(gate88inter4), .b(gate88inter3), .O(gate88inter5));
  nor2  gate777(.a(gate88inter5), .b(gate88inter2), .O(gate88inter6));
  inv1  gate778(.a(G16), .O(gate88inter7));
  inv1  gate779(.a(G335), .O(gate88inter8));
  nand2 gate780(.a(gate88inter8), .b(gate88inter7), .O(gate88inter9));
  nand2 gate781(.a(s_33), .b(gate88inter3), .O(gate88inter10));
  nor2  gate782(.a(gate88inter10), .b(gate88inter9), .O(gate88inter11));
  nor2  gate783(.a(gate88inter11), .b(gate88inter6), .O(gate88inter12));
  nand2 gate784(.a(gate88inter12), .b(gate88inter1), .O(G409));
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );

  xor2  gate981(.a(G344), .b(G22), .O(gate94inter0));
  nand2 gate982(.a(gate94inter0), .b(s_62), .O(gate94inter1));
  and2  gate983(.a(G344), .b(G22), .O(gate94inter2));
  inv1  gate984(.a(s_62), .O(gate94inter3));
  inv1  gate985(.a(s_63), .O(gate94inter4));
  nand2 gate986(.a(gate94inter4), .b(gate94inter3), .O(gate94inter5));
  nor2  gate987(.a(gate94inter5), .b(gate94inter2), .O(gate94inter6));
  inv1  gate988(.a(G22), .O(gate94inter7));
  inv1  gate989(.a(G344), .O(gate94inter8));
  nand2 gate990(.a(gate94inter8), .b(gate94inter7), .O(gate94inter9));
  nand2 gate991(.a(s_63), .b(gate94inter3), .O(gate94inter10));
  nor2  gate992(.a(gate94inter10), .b(gate94inter9), .O(gate94inter11));
  nor2  gate993(.a(gate94inter11), .b(gate94inter6), .O(gate94inter12));
  nand2 gate994(.a(gate94inter12), .b(gate94inter1), .O(G415));
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );

  xor2  gate547(.a(G350), .b(G23), .O(gate98inter0));
  nand2 gate548(.a(gate98inter0), .b(s_0), .O(gate98inter1));
  and2  gate549(.a(G350), .b(G23), .O(gate98inter2));
  inv1  gate550(.a(s_0), .O(gate98inter3));
  inv1  gate551(.a(s_1), .O(gate98inter4));
  nand2 gate552(.a(gate98inter4), .b(gate98inter3), .O(gate98inter5));
  nor2  gate553(.a(gate98inter5), .b(gate98inter2), .O(gate98inter6));
  inv1  gate554(.a(G23), .O(gate98inter7));
  inv1  gate555(.a(G350), .O(gate98inter8));
  nand2 gate556(.a(gate98inter8), .b(gate98inter7), .O(gate98inter9));
  nand2 gate557(.a(s_1), .b(gate98inter3), .O(gate98inter10));
  nor2  gate558(.a(gate98inter10), .b(gate98inter9), .O(gate98inter11));
  nor2  gate559(.a(gate98inter11), .b(gate98inter6), .O(gate98inter12));
  nand2 gate560(.a(gate98inter12), .b(gate98inter1), .O(G419));
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );

  xor2  gate1093(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate1094(.a(gate103inter0), .b(s_78), .O(gate103inter1));
  and2  gate1095(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate1096(.a(s_78), .O(gate103inter3));
  inv1  gate1097(.a(s_79), .O(gate103inter4));
  nand2 gate1098(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate1099(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate1100(.a(G28), .O(gate103inter7));
  inv1  gate1101(.a(G359), .O(gate103inter8));
  nand2 gate1102(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate1103(.a(s_79), .b(gate103inter3), .O(gate103inter10));
  nor2  gate1104(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate1105(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate1106(.a(gate103inter12), .b(gate103inter1), .O(G424));
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );

  xor2  gate659(.a(G379), .b(G378), .O(gate113inter0));
  nand2 gate660(.a(gate113inter0), .b(s_16), .O(gate113inter1));
  and2  gate661(.a(G379), .b(G378), .O(gate113inter2));
  inv1  gate662(.a(s_16), .O(gate113inter3));
  inv1  gate663(.a(s_17), .O(gate113inter4));
  nand2 gate664(.a(gate113inter4), .b(gate113inter3), .O(gate113inter5));
  nor2  gate665(.a(gate113inter5), .b(gate113inter2), .O(gate113inter6));
  inv1  gate666(.a(G378), .O(gate113inter7));
  inv1  gate667(.a(G379), .O(gate113inter8));
  nand2 gate668(.a(gate113inter8), .b(gate113inter7), .O(gate113inter9));
  nand2 gate669(.a(s_17), .b(gate113inter3), .O(gate113inter10));
  nor2  gate670(.a(gate113inter10), .b(gate113inter9), .O(gate113inter11));
  nor2  gate671(.a(gate113inter11), .b(gate113inter6), .O(gate113inter12));
  nand2 gate672(.a(gate113inter12), .b(gate113inter1), .O(G450));
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate701(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate702(.a(gate116inter0), .b(s_22), .O(gate116inter1));
  and2  gate703(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate704(.a(s_22), .O(gate116inter3));
  inv1  gate705(.a(s_23), .O(gate116inter4));
  nand2 gate706(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate707(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate708(.a(G384), .O(gate116inter7));
  inv1  gate709(.a(G385), .O(gate116inter8));
  nand2 gate710(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate711(.a(s_23), .b(gate116inter3), .O(gate116inter10));
  nor2  gate712(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate713(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate714(.a(gate116inter12), .b(gate116inter1), .O(G459));

  xor2  gate953(.a(G387), .b(G386), .O(gate117inter0));
  nand2 gate954(.a(gate117inter0), .b(s_58), .O(gate117inter1));
  and2  gate955(.a(G387), .b(G386), .O(gate117inter2));
  inv1  gate956(.a(s_58), .O(gate117inter3));
  inv1  gate957(.a(s_59), .O(gate117inter4));
  nand2 gate958(.a(gate117inter4), .b(gate117inter3), .O(gate117inter5));
  nor2  gate959(.a(gate117inter5), .b(gate117inter2), .O(gate117inter6));
  inv1  gate960(.a(G386), .O(gate117inter7));
  inv1  gate961(.a(G387), .O(gate117inter8));
  nand2 gate962(.a(gate117inter8), .b(gate117inter7), .O(gate117inter9));
  nand2 gate963(.a(s_59), .b(gate117inter3), .O(gate117inter10));
  nor2  gate964(.a(gate117inter10), .b(gate117inter9), .O(gate117inter11));
  nor2  gate965(.a(gate117inter11), .b(gate117inter6), .O(gate117inter12));
  nand2 gate966(.a(gate117inter12), .b(gate117inter1), .O(G462));
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );

  xor2  gate827(.a(G419), .b(G418), .O(gate133inter0));
  nand2 gate828(.a(gate133inter0), .b(s_40), .O(gate133inter1));
  and2  gate829(.a(G419), .b(G418), .O(gate133inter2));
  inv1  gate830(.a(s_40), .O(gate133inter3));
  inv1  gate831(.a(s_41), .O(gate133inter4));
  nand2 gate832(.a(gate133inter4), .b(gate133inter3), .O(gate133inter5));
  nor2  gate833(.a(gate133inter5), .b(gate133inter2), .O(gate133inter6));
  inv1  gate834(.a(G418), .O(gate133inter7));
  inv1  gate835(.a(G419), .O(gate133inter8));
  nand2 gate836(.a(gate133inter8), .b(gate133inter7), .O(gate133inter9));
  nand2 gate837(.a(s_41), .b(gate133inter3), .O(gate133inter10));
  nor2  gate838(.a(gate133inter10), .b(gate133inter9), .O(gate133inter11));
  nor2  gate839(.a(gate133inter11), .b(gate133inter6), .O(gate133inter12));
  nand2 gate840(.a(gate133inter12), .b(gate133inter1), .O(G510));
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate757(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate758(.a(gate137inter0), .b(s_30), .O(gate137inter1));
  and2  gate759(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate760(.a(s_30), .O(gate137inter3));
  inv1  gate761(.a(s_31), .O(gate137inter4));
  nand2 gate762(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate763(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate764(.a(G426), .O(gate137inter7));
  inv1  gate765(.a(G429), .O(gate137inter8));
  nand2 gate766(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate767(.a(s_31), .b(gate137inter3), .O(gate137inter10));
  nor2  gate768(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate769(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate770(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );

  xor2  gate687(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate688(.a(gate140inter0), .b(s_20), .O(gate140inter1));
  and2  gate689(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate690(.a(s_20), .O(gate140inter3));
  inv1  gate691(.a(s_21), .O(gate140inter4));
  nand2 gate692(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate693(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate694(.a(G444), .O(gate140inter7));
  inv1  gate695(.a(G447), .O(gate140inter8));
  nand2 gate696(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate697(.a(s_21), .b(gate140inter3), .O(gate140inter10));
  nor2  gate698(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate699(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate700(.a(gate140inter12), .b(gate140inter1), .O(G531));
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );

  xor2  gate1037(.a(G522), .b(G426), .O(gate153inter0));
  nand2 gate1038(.a(gate153inter0), .b(s_70), .O(gate153inter1));
  and2  gate1039(.a(G522), .b(G426), .O(gate153inter2));
  inv1  gate1040(.a(s_70), .O(gate153inter3));
  inv1  gate1041(.a(s_71), .O(gate153inter4));
  nand2 gate1042(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate1043(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate1044(.a(G426), .O(gate153inter7));
  inv1  gate1045(.a(G522), .O(gate153inter8));
  nand2 gate1046(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate1047(.a(s_71), .b(gate153inter3), .O(gate153inter10));
  nor2  gate1048(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate1049(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate1050(.a(gate153inter12), .b(gate153inter1), .O(G570));

  xor2  gate869(.a(G522), .b(G429), .O(gate154inter0));
  nand2 gate870(.a(gate154inter0), .b(s_46), .O(gate154inter1));
  and2  gate871(.a(G522), .b(G429), .O(gate154inter2));
  inv1  gate872(.a(s_46), .O(gate154inter3));
  inv1  gate873(.a(s_47), .O(gate154inter4));
  nand2 gate874(.a(gate154inter4), .b(gate154inter3), .O(gate154inter5));
  nor2  gate875(.a(gate154inter5), .b(gate154inter2), .O(gate154inter6));
  inv1  gate876(.a(G429), .O(gate154inter7));
  inv1  gate877(.a(G522), .O(gate154inter8));
  nand2 gate878(.a(gate154inter8), .b(gate154inter7), .O(gate154inter9));
  nand2 gate879(.a(s_47), .b(gate154inter3), .O(gate154inter10));
  nor2  gate880(.a(gate154inter10), .b(gate154inter9), .O(gate154inter11));
  nor2  gate881(.a(gate154inter11), .b(gate154inter6), .O(gate154inter12));
  nand2 gate882(.a(gate154inter12), .b(gate154inter1), .O(G571));
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );
nand2 gate165( .a(G462), .b(G540), .O(G582) );
nand2 gate166( .a(G465), .b(G540), .O(G583) );
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );
nand2 gate173( .a(G486), .b(G552), .O(G590) );
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );
nand2 gate183( .a(G516), .b(G567), .O(G600) );
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate967(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate968(.a(gate197inter0), .b(s_60), .O(gate197inter1));
  and2  gate969(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate970(.a(s_60), .O(gate197inter3));
  inv1  gate971(.a(s_61), .O(gate197inter4));
  nand2 gate972(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate973(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate974(.a(G594), .O(gate197inter7));
  inv1  gate975(.a(G595), .O(gate197inter8));
  nand2 gate976(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate977(.a(s_61), .b(gate197inter3), .O(gate197inter10));
  nor2  gate978(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate979(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate980(.a(gate197inter12), .b(gate197inter1), .O(G654));

  xor2  gate1107(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate1108(.a(gate198inter0), .b(s_80), .O(gate198inter1));
  and2  gate1109(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate1110(.a(s_80), .O(gate198inter3));
  inv1  gate1111(.a(s_81), .O(gate198inter4));
  nand2 gate1112(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate1113(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate1114(.a(G596), .O(gate198inter7));
  inv1  gate1115(.a(G597), .O(gate198inter8));
  nand2 gate1116(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate1117(.a(s_81), .b(gate198inter3), .O(gate198inter10));
  nor2  gate1118(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate1119(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate1120(.a(gate198inter12), .b(gate198inter1), .O(G657));
nand2 gate199( .a(G598), .b(G599), .O(G660) );
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate1065(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate1066(.a(gate203inter0), .b(s_74), .O(gate203inter1));
  and2  gate1067(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate1068(.a(s_74), .O(gate203inter3));
  inv1  gate1069(.a(s_75), .O(gate203inter4));
  nand2 gate1070(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate1071(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate1072(.a(G602), .O(gate203inter7));
  inv1  gate1073(.a(G612), .O(gate203inter8));
  nand2 gate1074(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate1075(.a(s_75), .b(gate203inter3), .O(gate203inter10));
  nor2  gate1076(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate1077(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate1078(.a(gate203inter12), .b(gate203inter1), .O(G672));

  xor2  gate1135(.a(G617), .b(G607), .O(gate204inter0));
  nand2 gate1136(.a(gate204inter0), .b(s_84), .O(gate204inter1));
  and2  gate1137(.a(G617), .b(G607), .O(gate204inter2));
  inv1  gate1138(.a(s_84), .O(gate204inter3));
  inv1  gate1139(.a(s_85), .O(gate204inter4));
  nand2 gate1140(.a(gate204inter4), .b(gate204inter3), .O(gate204inter5));
  nor2  gate1141(.a(gate204inter5), .b(gate204inter2), .O(gate204inter6));
  inv1  gate1142(.a(G607), .O(gate204inter7));
  inv1  gate1143(.a(G617), .O(gate204inter8));
  nand2 gate1144(.a(gate204inter8), .b(gate204inter7), .O(gate204inter9));
  nand2 gate1145(.a(s_85), .b(gate204inter3), .O(gate204inter10));
  nor2  gate1146(.a(gate204inter10), .b(gate204inter9), .O(gate204inter11));
  nor2  gate1147(.a(gate204inter11), .b(gate204inter6), .O(gate204inter12));
  nand2 gate1148(.a(gate204inter12), .b(gate204inter1), .O(G675));
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );
nand2 gate220( .a(G637), .b(G681), .O(G701) );
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );
nand2 gate227( .a(G694), .b(G695), .O(G712) );
nand2 gate228( .a(G696), .b(G697), .O(G715) );

  xor2  gate799(.a(G699), .b(G698), .O(gate229inter0));
  nand2 gate800(.a(gate229inter0), .b(s_36), .O(gate229inter1));
  and2  gate801(.a(G699), .b(G698), .O(gate229inter2));
  inv1  gate802(.a(s_36), .O(gate229inter3));
  inv1  gate803(.a(s_37), .O(gate229inter4));
  nand2 gate804(.a(gate229inter4), .b(gate229inter3), .O(gate229inter5));
  nor2  gate805(.a(gate229inter5), .b(gate229inter2), .O(gate229inter6));
  inv1  gate806(.a(G698), .O(gate229inter7));
  inv1  gate807(.a(G699), .O(gate229inter8));
  nand2 gate808(.a(gate229inter8), .b(gate229inter7), .O(gate229inter9));
  nand2 gate809(.a(s_37), .b(gate229inter3), .O(gate229inter10));
  nor2  gate810(.a(gate229inter10), .b(gate229inter9), .O(gate229inter11));
  nor2  gate811(.a(gate229inter11), .b(gate229inter6), .O(gate229inter12));
  nand2 gate812(.a(gate229inter12), .b(gate229inter1), .O(G718));
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );

  xor2  gate1177(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate1178(.a(gate242inter0), .b(s_90), .O(gate242inter1));
  and2  gate1179(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate1180(.a(s_90), .O(gate242inter3));
  inv1  gate1181(.a(s_91), .O(gate242inter4));
  nand2 gate1182(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate1183(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate1184(.a(G718), .O(gate242inter7));
  inv1  gate1185(.a(G730), .O(gate242inter8));
  nand2 gate1186(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate1187(.a(s_91), .b(gate242inter3), .O(gate242inter10));
  nor2  gate1188(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate1189(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate1190(.a(gate242inter12), .b(gate242inter1), .O(G755));
nand2 gate243( .a(G245), .b(G733), .O(G756) );

  xor2  gate561(.a(G733), .b(G721), .O(gate244inter0));
  nand2 gate562(.a(gate244inter0), .b(s_2), .O(gate244inter1));
  and2  gate563(.a(G733), .b(G721), .O(gate244inter2));
  inv1  gate564(.a(s_2), .O(gate244inter3));
  inv1  gate565(.a(s_3), .O(gate244inter4));
  nand2 gate566(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate567(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate568(.a(G721), .O(gate244inter7));
  inv1  gate569(.a(G733), .O(gate244inter8));
  nand2 gate570(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate571(.a(s_3), .b(gate244inter3), .O(gate244inter10));
  nor2  gate572(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate573(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate574(.a(gate244inter12), .b(gate244inter1), .O(G757));
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );
nand2 gate252( .a(G709), .b(G745), .O(G765) );
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );

  xor2  gate855(.a(G755), .b(G754), .O(gate257inter0));
  nand2 gate856(.a(gate257inter0), .b(s_44), .O(gate257inter1));
  and2  gate857(.a(G755), .b(G754), .O(gate257inter2));
  inv1  gate858(.a(s_44), .O(gate257inter3));
  inv1  gate859(.a(s_45), .O(gate257inter4));
  nand2 gate860(.a(gate257inter4), .b(gate257inter3), .O(gate257inter5));
  nor2  gate861(.a(gate257inter5), .b(gate257inter2), .O(gate257inter6));
  inv1  gate862(.a(G754), .O(gate257inter7));
  inv1  gate863(.a(G755), .O(gate257inter8));
  nand2 gate864(.a(gate257inter8), .b(gate257inter7), .O(gate257inter9));
  nand2 gate865(.a(s_45), .b(gate257inter3), .O(gate257inter10));
  nor2  gate866(.a(gate257inter10), .b(gate257inter9), .O(gate257inter11));
  nor2  gate867(.a(gate257inter11), .b(gate257inter6), .O(gate257inter12));
  nand2 gate868(.a(gate257inter12), .b(gate257inter1), .O(G770));
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate1149(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate1150(.a(gate268inter0), .b(s_86), .O(gate268inter1));
  and2  gate1151(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate1152(.a(s_86), .O(gate268inter3));
  inv1  gate1153(.a(s_87), .O(gate268inter4));
  nand2 gate1154(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1155(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1156(.a(G651), .O(gate268inter7));
  inv1  gate1157(.a(G779), .O(gate268inter8));
  nand2 gate1158(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1159(.a(s_87), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1160(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1161(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1162(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );
nand2 gate273( .a(G642), .b(G794), .O(G818) );
nand2 gate274( .a(G770), .b(G794), .O(G819) );
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );
nand2 gate279( .a(G651), .b(G803), .O(G824) );
nand2 gate280( .a(G779), .b(G803), .O(G825) );
nand2 gate281( .a(G654), .b(G806), .O(G826) );

  xor2  gate645(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate646(.a(gate282inter0), .b(s_14), .O(gate282inter1));
  and2  gate647(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate648(.a(s_14), .O(gate282inter3));
  inv1  gate649(.a(s_15), .O(gate282inter4));
  nand2 gate650(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate651(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate652(.a(G782), .O(gate282inter7));
  inv1  gate653(.a(G806), .O(gate282inter8));
  nand2 gate654(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate655(.a(s_15), .b(gate282inter3), .O(gate282inter10));
  nor2  gate656(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate657(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate658(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );
nand2 gate284( .a(G785), .b(G809), .O(G829) );

  xor2  gate841(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate842(.a(gate285inter0), .b(s_42), .O(gate285inter1));
  and2  gate843(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate844(.a(s_42), .O(gate285inter3));
  inv1  gate845(.a(s_43), .O(gate285inter4));
  nand2 gate846(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate847(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate848(.a(G660), .O(gate285inter7));
  inv1  gate849(.a(G812), .O(gate285inter8));
  nand2 gate850(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate851(.a(s_43), .b(gate285inter3), .O(gate285inter10));
  nor2  gate852(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate853(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate854(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );
nand2 gate291( .a(G822), .b(G823), .O(G860) );
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );

  xor2  gate729(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate730(.a(gate391inter0), .b(s_26), .O(gate391inter1));
  and2  gate731(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate732(.a(s_26), .O(gate391inter3));
  inv1  gate733(.a(s_27), .O(gate391inter4));
  nand2 gate734(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate735(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate736(.a(G5), .O(gate391inter7));
  inv1  gate737(.a(G1048), .O(gate391inter8));
  nand2 gate738(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate739(.a(s_27), .b(gate391inter3), .O(gate391inter10));
  nor2  gate740(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate741(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate742(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );
nand2 gate408( .a(G22), .b(G1099), .O(G1195) );
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );
nand2 gate418( .a(G32), .b(G1129), .O(G1225) );
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );

  xor2  gate743(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate744(.a(gate420inter0), .b(s_28), .O(gate420inter1));
  and2  gate745(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate746(.a(s_28), .O(gate420inter3));
  inv1  gate747(.a(s_29), .O(gate420inter4));
  nand2 gate748(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate749(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate750(.a(G1036), .O(gate420inter7));
  inv1  gate751(.a(G1132), .O(gate420inter8));
  nand2 gate752(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate753(.a(s_29), .b(gate420inter3), .O(gate420inter10));
  nor2  gate754(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate755(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate756(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );

  xor2  gate631(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate632(.a(gate423inter0), .b(s_12), .O(gate423inter1));
  and2  gate633(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate634(.a(s_12), .O(gate423inter3));
  inv1  gate635(.a(s_13), .O(gate423inter4));
  nand2 gate636(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate637(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate638(.a(G3), .O(gate423inter7));
  inv1  gate639(.a(G1138), .O(gate423inter8));
  nand2 gate640(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate641(.a(s_13), .b(gate423inter3), .O(gate423inter10));
  nor2  gate642(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate643(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate644(.a(gate423inter12), .b(gate423inter1), .O(G1232));
nand2 gate424( .a(G1042), .b(G1138), .O(G1233) );
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );
nand2 gate442( .a(G1069), .b(G1165), .O(G1251) );
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );

  xor2  gate883(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate884(.a(gate449inter0), .b(s_48), .O(gate449inter1));
  and2  gate885(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate886(.a(s_48), .O(gate449inter3));
  inv1  gate887(.a(s_49), .O(gate449inter4));
  nand2 gate888(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate889(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate890(.a(G16), .O(gate449inter7));
  inv1  gate891(.a(G1177), .O(gate449inter8));
  nand2 gate892(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate893(.a(s_49), .b(gate449inter3), .O(gate449inter10));
  nor2  gate894(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate895(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate896(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );

  xor2  gate995(.a(G1192), .b(G1096), .O(gate460inter0));
  nand2 gate996(.a(gate460inter0), .b(s_64), .O(gate460inter1));
  and2  gate997(.a(G1192), .b(G1096), .O(gate460inter2));
  inv1  gate998(.a(s_64), .O(gate460inter3));
  inv1  gate999(.a(s_65), .O(gate460inter4));
  nand2 gate1000(.a(gate460inter4), .b(gate460inter3), .O(gate460inter5));
  nor2  gate1001(.a(gate460inter5), .b(gate460inter2), .O(gate460inter6));
  inv1  gate1002(.a(G1096), .O(gate460inter7));
  inv1  gate1003(.a(G1192), .O(gate460inter8));
  nand2 gate1004(.a(gate460inter8), .b(gate460inter7), .O(gate460inter9));
  nand2 gate1005(.a(s_65), .b(gate460inter3), .O(gate460inter10));
  nor2  gate1006(.a(gate460inter10), .b(gate460inter9), .O(gate460inter11));
  nor2  gate1007(.a(gate460inter11), .b(gate460inter6), .O(gate460inter12));
  nand2 gate1008(.a(gate460inter12), .b(gate460inter1), .O(G1269));
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );

  xor2  gate939(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate940(.a(gate462inter0), .b(s_56), .O(gate462inter1));
  and2  gate941(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate942(.a(s_56), .O(gate462inter3));
  inv1  gate943(.a(s_57), .O(gate462inter4));
  nand2 gate944(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate945(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate946(.a(G1099), .O(gate462inter7));
  inv1  gate947(.a(G1195), .O(gate462inter8));
  nand2 gate948(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate949(.a(s_57), .b(gate462inter3), .O(gate462inter10));
  nor2  gate950(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate951(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate952(.a(gate462inter12), .b(gate462inter1), .O(G1271));

  xor2  gate589(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate590(.a(gate463inter0), .b(s_6), .O(gate463inter1));
  and2  gate591(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate592(.a(s_6), .O(gate463inter3));
  inv1  gate593(.a(s_7), .O(gate463inter4));
  nand2 gate594(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate595(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate596(.a(G23), .O(gate463inter7));
  inv1  gate597(.a(G1198), .O(gate463inter8));
  nand2 gate598(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate599(.a(s_7), .b(gate463inter3), .O(gate463inter10));
  nor2  gate600(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate601(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate602(.a(gate463inter12), .b(gate463inter1), .O(G1272));
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );
nand2 gate466( .a(G1105), .b(G1201), .O(G1275) );
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );

  xor2  gate813(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate814(.a(gate472inter0), .b(s_38), .O(gate472inter1));
  and2  gate815(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate816(.a(s_38), .O(gate472inter3));
  inv1  gate817(.a(s_39), .O(gate472inter4));
  nand2 gate818(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate819(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate820(.a(G1114), .O(gate472inter7));
  inv1  gate821(.a(G1210), .O(gate472inter8));
  nand2 gate822(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate823(.a(s_39), .b(gate472inter3), .O(gate472inter10));
  nor2  gate824(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate825(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate826(.a(gate472inter12), .b(gate472inter1), .O(G1281));
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );

  xor2  gate673(.a(G1222), .b(G31), .O(gate479inter0));
  nand2 gate674(.a(gate479inter0), .b(s_18), .O(gate479inter1));
  and2  gate675(.a(G1222), .b(G31), .O(gate479inter2));
  inv1  gate676(.a(s_18), .O(gate479inter3));
  inv1  gate677(.a(s_19), .O(gate479inter4));
  nand2 gate678(.a(gate479inter4), .b(gate479inter3), .O(gate479inter5));
  nor2  gate679(.a(gate479inter5), .b(gate479inter2), .O(gate479inter6));
  inv1  gate680(.a(G31), .O(gate479inter7));
  inv1  gate681(.a(G1222), .O(gate479inter8));
  nand2 gate682(.a(gate479inter8), .b(gate479inter7), .O(gate479inter9));
  nand2 gate683(.a(s_19), .b(gate479inter3), .O(gate479inter10));
  nor2  gate684(.a(gate479inter10), .b(gate479inter9), .O(gate479inter11));
  nor2  gate685(.a(gate479inter11), .b(gate479inter6), .O(gate479inter12));
  nand2 gate686(.a(gate479inter12), .b(gate479inter1), .O(G1288));
nand2 gate480( .a(G1126), .b(G1222), .O(G1289) );
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );

  xor2  gate617(.a(G1231), .b(G1230), .O(gate484inter0));
  nand2 gate618(.a(gate484inter0), .b(s_10), .O(gate484inter1));
  and2  gate619(.a(G1231), .b(G1230), .O(gate484inter2));
  inv1  gate620(.a(s_10), .O(gate484inter3));
  inv1  gate621(.a(s_11), .O(gate484inter4));
  nand2 gate622(.a(gate484inter4), .b(gate484inter3), .O(gate484inter5));
  nor2  gate623(.a(gate484inter5), .b(gate484inter2), .O(gate484inter6));
  inv1  gate624(.a(G1230), .O(gate484inter7));
  inv1  gate625(.a(G1231), .O(gate484inter8));
  nand2 gate626(.a(gate484inter8), .b(gate484inter7), .O(gate484inter9));
  nand2 gate627(.a(s_11), .b(gate484inter3), .O(gate484inter10));
  nor2  gate628(.a(gate484inter10), .b(gate484inter9), .O(gate484inter11));
  nor2  gate629(.a(gate484inter11), .b(gate484inter6), .O(gate484inter12));
  nand2 gate630(.a(gate484inter12), .b(gate484inter1), .O(G1293));
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );

  xor2  gate911(.a(G1237), .b(G1236), .O(gate487inter0));
  nand2 gate912(.a(gate487inter0), .b(s_52), .O(gate487inter1));
  and2  gate913(.a(G1237), .b(G1236), .O(gate487inter2));
  inv1  gate914(.a(s_52), .O(gate487inter3));
  inv1  gate915(.a(s_53), .O(gate487inter4));
  nand2 gate916(.a(gate487inter4), .b(gate487inter3), .O(gate487inter5));
  nor2  gate917(.a(gate487inter5), .b(gate487inter2), .O(gate487inter6));
  inv1  gate918(.a(G1236), .O(gate487inter7));
  inv1  gate919(.a(G1237), .O(gate487inter8));
  nand2 gate920(.a(gate487inter8), .b(gate487inter7), .O(gate487inter9));
  nand2 gate921(.a(s_53), .b(gate487inter3), .O(gate487inter10));
  nor2  gate922(.a(gate487inter10), .b(gate487inter9), .O(gate487inter11));
  nor2  gate923(.a(gate487inter11), .b(gate487inter6), .O(gate487inter12));
  nand2 gate924(.a(gate487inter12), .b(gate487inter1), .O(G1296));

  xor2  gate1023(.a(G1239), .b(G1238), .O(gate488inter0));
  nand2 gate1024(.a(gate488inter0), .b(s_68), .O(gate488inter1));
  and2  gate1025(.a(G1239), .b(G1238), .O(gate488inter2));
  inv1  gate1026(.a(s_68), .O(gate488inter3));
  inv1  gate1027(.a(s_69), .O(gate488inter4));
  nand2 gate1028(.a(gate488inter4), .b(gate488inter3), .O(gate488inter5));
  nor2  gate1029(.a(gate488inter5), .b(gate488inter2), .O(gate488inter6));
  inv1  gate1030(.a(G1238), .O(gate488inter7));
  inv1  gate1031(.a(G1239), .O(gate488inter8));
  nand2 gate1032(.a(gate488inter8), .b(gate488inter7), .O(gate488inter9));
  nand2 gate1033(.a(s_69), .b(gate488inter3), .O(gate488inter10));
  nor2  gate1034(.a(gate488inter10), .b(gate488inter9), .O(gate488inter11));
  nor2  gate1035(.a(gate488inter11), .b(gate488inter6), .O(gate488inter12));
  nand2 gate1036(.a(gate488inter12), .b(gate488inter1), .O(G1297));

  xor2  gate1079(.a(G1241), .b(G1240), .O(gate489inter0));
  nand2 gate1080(.a(gate489inter0), .b(s_76), .O(gate489inter1));
  and2  gate1081(.a(G1241), .b(G1240), .O(gate489inter2));
  inv1  gate1082(.a(s_76), .O(gate489inter3));
  inv1  gate1083(.a(s_77), .O(gate489inter4));
  nand2 gate1084(.a(gate489inter4), .b(gate489inter3), .O(gate489inter5));
  nor2  gate1085(.a(gate489inter5), .b(gate489inter2), .O(gate489inter6));
  inv1  gate1086(.a(G1240), .O(gate489inter7));
  inv1  gate1087(.a(G1241), .O(gate489inter8));
  nand2 gate1088(.a(gate489inter8), .b(gate489inter7), .O(gate489inter9));
  nand2 gate1089(.a(s_77), .b(gate489inter3), .O(gate489inter10));
  nor2  gate1090(.a(gate489inter10), .b(gate489inter9), .O(gate489inter11));
  nor2  gate1091(.a(gate489inter11), .b(gate489inter6), .O(gate489inter12));
  nand2 gate1092(.a(gate489inter12), .b(gate489inter1), .O(G1298));
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );

  xor2  gate715(.a(G1251), .b(G1250), .O(gate494inter0));
  nand2 gate716(.a(gate494inter0), .b(s_24), .O(gate494inter1));
  and2  gate717(.a(G1251), .b(G1250), .O(gate494inter2));
  inv1  gate718(.a(s_24), .O(gate494inter3));
  inv1  gate719(.a(s_25), .O(gate494inter4));
  nand2 gate720(.a(gate494inter4), .b(gate494inter3), .O(gate494inter5));
  nor2  gate721(.a(gate494inter5), .b(gate494inter2), .O(gate494inter6));
  inv1  gate722(.a(G1250), .O(gate494inter7));
  inv1  gate723(.a(G1251), .O(gate494inter8));
  nand2 gate724(.a(gate494inter8), .b(gate494inter7), .O(gate494inter9));
  nand2 gate725(.a(s_25), .b(gate494inter3), .O(gate494inter10));
  nor2  gate726(.a(gate494inter10), .b(gate494inter9), .O(gate494inter11));
  nor2  gate727(.a(gate494inter11), .b(gate494inter6), .O(gate494inter12));
  nand2 gate728(.a(gate494inter12), .b(gate494inter1), .O(G1303));
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );

  xor2  gate925(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate926(.a(gate511inter0), .b(s_54), .O(gate511inter1));
  and2  gate927(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate928(.a(s_54), .O(gate511inter3));
  inv1  gate929(.a(s_55), .O(gate511inter4));
  nand2 gate930(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate931(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate932(.a(G1284), .O(gate511inter7));
  inv1  gate933(.a(G1285), .O(gate511inter8));
  nand2 gate934(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate935(.a(s_55), .b(gate511inter3), .O(gate511inter10));
  nor2  gate936(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate937(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate938(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule