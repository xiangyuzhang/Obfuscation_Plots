module c880 (N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,
             N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,
             N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,
             N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,
             N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,
             N219,N228,N237,N246,N255,N259,N260,N261,N267,N268,
             N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,
             N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,
             N865,N866,N874,N878,N879,N880);
input N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,
      N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,
      N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,
      N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,
      N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,
      N219,N228,N237,N246,N255,N259,N260,N261,N267,N268;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81;
output N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,
       N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,
       N865,N866,N874,N878,N879,N880;
wire N269,N270,N273,N276,N279,N280,N284,N285,N286,N287,
     N290,N291,N292,N293,N294,N295,N296,N297,N298,N301,
     N302,N303,N304,N305,N306,N307,N308,N309,N310,N316,
     N317,N318,N319,N322,N323,N324,N325,N326,N327,N328,
     N329,N330,N331,N332,N333,N334,N335,N336,N337,N338,
     N339,N340,N341,N342,N343,N344,N345,N346,N347,N348,
     N349,N350,N351,N352,N353,N354,N355,N356,N357,N360,
     N363,N366,N369,N375,N376,N379,N382,N385,N392,N393,
     N399,N400,N401,N402,N403,N404,N405,N406,N407,N408,
     N409,N410,N411,N412,N413,N414,N415,N416,N417,N424,
     N425,N426,N427,N432,N437,N442,N443,N444,N445,N451,
     N460,N463,N466,N475,N476,N477,N478,N479,N480,N481,
     N482,N483,N488,N489,N490,N491,N492,N495,N498,N499,
     N500,N501,N502,N503,N504,N505,N506,N507,N508,N509,
     N510,N511,N512,N513,N514,N515,N516,N517,N518,N519,
     N520,N521,N522,N523,N524,N525,N526,N527,N528,N529,
     N530,N533,N536,N537,N538,N539,N540,N541,N542,N543,
     N544,N547,N550,N551,N552,N553,N557,N561,N565,N569,
     N573,N577,N581,N585,N586,N587,N588,N589,N590,N593,
     N596,N597,N600,N605,N606,N609,N615,N616,N619,N624,
     N625,N628,N631,N632,N635,N640,N641,N644,N650,N651,
     N654,N659,N660,N661,N662,N665,N669,N670,N673,N677,
     N678,N682,N686,N687,N692,N696,N697,N700,N704,N705,
     N708,N712,N713,N717,N721,N722,N727,N731,N732,N733,
     N734,N735,N736,N737,N738,N739,N740,N741,N742,N743,
     N744,N745,N746,N747,N748,N749,N750,N751,N752,N753,
     N754,N755,N756,N757,N758,N759,N760,N761,N762,N763,
     N764,N765,N766,N769,N770,N771,N772,N773,N777,N778,
     N781,N782,N785,N786,N787,N788,N789,N790,N791,N792,
     N793,N794,N795,N796,N802,N803,N804,N805,N806,N807,
     N808,N809,N810,N811,N812,N813,N814,N815,N819,N822,
     N825,N826,N827,N828,N829,N830,N831,N832,N833,N834,
     N835,N836,N837,N838,N839,N840,N841,N842,N843,N844,
     N845,N846,N847,N848,N849,N851,N852,N853,N854,N855,
     N856,N857,N858,N859,N860,N861,N862,N867,N868,N869,
     N870,N871,N872,N873,N875,N876,N877, gate180inter0, gate180inter1, gate180inter2, gate180inter3, gate180inter4, gate180inter5, gate180inter6, gate180inter7, gate180inter8, gate180inter9, gate180inter10, gate180inter11, gate180inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate244inter0, gate244inter1, gate244inter2, gate244inter3, gate244inter4, gate244inter5, gate244inter6, gate244inter7, gate244inter8, gate244inter9, gate244inter10, gate244inter11, gate244inter12, gate238inter0, gate238inter1, gate238inter2, gate238inter3, gate238inter4, gate238inter5, gate238inter6, gate238inter7, gate238inter8, gate238inter9, gate238inter10, gate238inter11, gate238inter12, gate315inter0, gate315inter1, gate315inter2, gate315inter3, gate315inter4, gate315inter5, gate315inter6, gate315inter7, gate315inter8, gate315inter9, gate315inter10, gate315inter11, gate315inter12, gate181inter0, gate181inter1, gate181inter2, gate181inter3, gate181inter4, gate181inter5, gate181inter6, gate181inter7, gate181inter8, gate181inter9, gate181inter10, gate181inter11, gate181inter12, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate254inter0, gate254inter1, gate254inter2, gate254inter3, gate254inter4, gate254inter5, gate254inter6, gate254inter7, gate254inter8, gate254inter9, gate254inter10, gate254inter11, gate254inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate235inter0, gate235inter1, gate235inter2, gate235inter3, gate235inter4, gate235inter5, gate235inter6, gate235inter7, gate235inter8, gate235inter9, gate235inter10, gate235inter11, gate235inter12, gate42inter0, gate42inter1, gate42inter2, gate42inter3, gate42inter4, gate42inter5, gate42inter6, gate42inter7, gate42inter8, gate42inter9, gate42inter10, gate42inter11, gate42inter12, gate216inter0, gate216inter1, gate216inter2, gate216inter3, gate216inter4, gate216inter5, gate216inter6, gate216inter7, gate216inter8, gate216inter9, gate216inter10, gate216inter11, gate216inter12, gate337inter0, gate337inter1, gate337inter2, gate337inter3, gate337inter4, gate337inter5, gate337inter6, gate337inter7, gate337inter8, gate337inter9, gate337inter10, gate337inter11, gate337inter12, gate294inter0, gate294inter1, gate294inter2, gate294inter3, gate294inter4, gate294inter5, gate294inter6, gate294inter7, gate294inter8, gate294inter9, gate294inter10, gate294inter11, gate294inter12, gate310inter0, gate310inter1, gate310inter2, gate310inter3, gate310inter4, gate310inter5, gate310inter6, gate310inter7, gate310inter8, gate310inter9, gate310inter10, gate310inter11, gate310inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate192inter0, gate192inter1, gate192inter2, gate192inter3, gate192inter4, gate192inter5, gate192inter6, gate192inter7, gate192inter8, gate192inter9, gate192inter10, gate192inter11, gate192inter12, gate314inter0, gate314inter1, gate314inter2, gate314inter3, gate314inter4, gate314inter5, gate314inter6, gate314inter7, gate314inter8, gate314inter9, gate314inter10, gate314inter11, gate314inter12, gate151inter0, gate151inter1, gate151inter2, gate151inter3, gate151inter4, gate151inter5, gate151inter6, gate151inter7, gate151inter8, gate151inter9, gate151inter10, gate151inter11, gate151inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate333inter0, gate333inter1, gate333inter2, gate333inter3, gate333inter4, gate333inter5, gate333inter6, gate333inter7, gate333inter8, gate333inter9, gate333inter10, gate333inter11, gate333inter12, gate70inter0, gate70inter1, gate70inter2, gate70inter3, gate70inter4, gate70inter5, gate70inter6, gate70inter7, gate70inter8, gate70inter9, gate70inter10, gate70inter11, gate70inter12, gate186inter0, gate186inter1, gate186inter2, gate186inter3, gate186inter4, gate186inter5, gate186inter6, gate186inter7, gate186inter8, gate186inter9, gate186inter10, gate186inter11, gate186inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate26inter0, gate26inter1, gate26inter2, gate26inter3, gate26inter4, gate26inter5, gate26inter6, gate26inter7, gate26inter8, gate26inter9, gate26inter10, gate26inter11, gate26inter12, gate128inter0, gate128inter1, gate128inter2, gate128inter3, gate128inter4, gate128inter5, gate128inter6, gate128inter7, gate128inter8, gate128inter9, gate128inter10, gate128inter11, gate128inter12, gate348inter0, gate348inter1, gate348inter2, gate348inter3, gate348inter4, gate348inter5, gate348inter6, gate348inter7, gate348inter8, gate348inter9, gate348inter10, gate348inter11, gate348inter12, gate191inter0, gate191inter1, gate191inter2, gate191inter3, gate191inter4, gate191inter5, gate191inter6, gate191inter7, gate191inter8, gate191inter9, gate191inter10, gate191inter11, gate191inter12, gate155inter0, gate155inter1, gate155inter2, gate155inter3, gate155inter4, gate155inter5, gate155inter6, gate155inter7, gate155inter8, gate155inter9, gate155inter10, gate155inter11, gate155inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate149inter0, gate149inter1, gate149inter2, gate149inter3, gate149inter4, gate149inter5, gate149inter6, gate149inter7, gate149inter8, gate149inter9, gate149inter10, gate149inter11, gate149inter12, gate36inter0, gate36inter1, gate36inter2, gate36inter3, gate36inter4, gate36inter5, gate36inter6, gate36inter7, gate36inter8, gate36inter9, gate36inter10, gate36inter11, gate36inter12, gate177inter0, gate177inter1, gate177inter2, gate177inter3, gate177inter4, gate177inter5, gate177inter6, gate177inter7, gate177inter8, gate177inter9, gate177inter10, gate177inter11, gate177inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate153inter0, gate153inter1, gate153inter2, gate153inter3, gate153inter4, gate153inter5, gate153inter6, gate153inter7, gate153inter8, gate153inter9, gate153inter10, gate153inter11, gate153inter12, gate299inter0, gate299inter1, gate299inter2, gate299inter3, gate299inter4, gate299inter5, gate299inter6, gate299inter7, gate299inter8, gate299inter9, gate299inter10, gate299inter11, gate299inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate225inter0, gate225inter1, gate225inter2, gate225inter3, gate225inter4, gate225inter5, gate225inter6, gate225inter7, gate225inter8, gate225inter9, gate225inter10, gate225inter11, gate225inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12;


nand4 gate1( .a(N1), .b(N8), .c(N13), .d(N17), .O(N269) );
nand4 gate2( .a(N1), .b(N26), .c(N13), .d(N17), .O(N270) );
and3 gate3( .a(N29), .b(N36), .c(N42), .O(N273) );
and3 gate4( .a(N1), .b(N26), .c(N51), .O(N276) );
nand4 gate5( .a(N1), .b(N8), .c(N51), .d(N17), .O(N279) );
nand4 gate6( .a(N1), .b(N8), .c(N13), .d(N55), .O(N280) );
nand4 gate7( .a(N59), .b(N42), .c(N68), .d(N72), .O(N284) );
nand2 gate8( .a(N29), .b(N68), .O(N285) );
nand3 gate9( .a(N59), .b(N68), .c(N74), .O(N286) );
and3 gate10( .a(N29), .b(N75), .c(N80), .O(N287) );
and3 gate11( .a(N29), .b(N75), .c(N42), .O(N290) );
and3 gate12( .a(N29), .b(N36), .c(N80), .O(N291) );
and3 gate13( .a(N29), .b(N36), .c(N42), .O(N292) );
and3 gate14( .a(N59), .b(N75), .c(N80), .O(N293) );
and3 gate15( .a(N59), .b(N75), .c(N42), .O(N294) );
and3 gate16( .a(N59), .b(N36), .c(N80), .O(N295) );
and3 gate17( .a(N59), .b(N36), .c(N42), .O(N296) );
and2 gate18( .a(N85), .b(N86), .O(N297) );
or2 gate19( .a(N87), .b(N88), .O(N298) );
nand2 gate20( .a(N91), .b(N96), .O(N301) );
or2 gate21( .a(N91), .b(N96), .O(N302) );
nand2 gate22( .a(N101), .b(N106), .O(N303) );
or2 gate23( .a(N101), .b(N106), .O(N304) );
nand2 gate24( .a(N111), .b(N116), .O(N305) );
or2 gate25( .a(N111), .b(N116), .O(N306) );

  xor2  gate734(.a(N126), .b(N121), .O(gate26inter0));
  nand2 gate735(.a(gate26inter0), .b(s_50), .O(gate26inter1));
  and2  gate736(.a(N126), .b(N121), .O(gate26inter2));
  inv1  gate737(.a(s_50), .O(gate26inter3));
  inv1  gate738(.a(s_51), .O(gate26inter4));
  nand2 gate739(.a(gate26inter4), .b(gate26inter3), .O(gate26inter5));
  nor2  gate740(.a(gate26inter5), .b(gate26inter2), .O(gate26inter6));
  inv1  gate741(.a(N121), .O(gate26inter7));
  inv1  gate742(.a(N126), .O(gate26inter8));
  nand2 gate743(.a(gate26inter8), .b(gate26inter7), .O(gate26inter9));
  nand2 gate744(.a(s_51), .b(gate26inter3), .O(gate26inter10));
  nor2  gate745(.a(gate26inter10), .b(gate26inter9), .O(gate26inter11));
  nor2  gate746(.a(gate26inter11), .b(gate26inter6), .O(gate26inter12));
  nand2 gate747(.a(gate26inter12), .b(gate26inter1), .O(N307));
or2 gate27( .a(N121), .b(N126), .O(N308) );
and2 gate28( .a(N8), .b(N138), .O(N309) );
inv1 gate29( .a(N268), .O(N310) );
and2 gate30( .a(N51), .b(N138), .O(N316) );
and2 gate31( .a(N17), .b(N138), .O(N317) );
and2 gate32( .a(N152), .b(N138), .O(N318) );
nand2 gate33( .a(N59), .b(N156), .O(N319) );
nor2 gate34( .a(N17), .b(N42), .O(N322) );
and2 gate35( .a(N17), .b(N42), .O(N323) );

  xor2  gate846(.a(N165), .b(N159), .O(gate36inter0));
  nand2 gate847(.a(gate36inter0), .b(s_66), .O(gate36inter1));
  and2  gate848(.a(N165), .b(N159), .O(gate36inter2));
  inv1  gate849(.a(s_66), .O(gate36inter3));
  inv1  gate850(.a(s_67), .O(gate36inter4));
  nand2 gate851(.a(gate36inter4), .b(gate36inter3), .O(gate36inter5));
  nor2  gate852(.a(gate36inter5), .b(gate36inter2), .O(gate36inter6));
  inv1  gate853(.a(N159), .O(gate36inter7));
  inv1  gate854(.a(N165), .O(gate36inter8));
  nand2 gate855(.a(gate36inter8), .b(gate36inter7), .O(gate36inter9));
  nand2 gate856(.a(s_67), .b(gate36inter3), .O(gate36inter10));
  nor2  gate857(.a(gate36inter10), .b(gate36inter9), .O(gate36inter11));
  nor2  gate858(.a(gate36inter11), .b(gate36inter6), .O(gate36inter12));
  nand2 gate859(.a(gate36inter12), .b(gate36inter1), .O(N324));
or2 gate37( .a(N159), .b(N165), .O(N325) );
nand2 gate38( .a(N171), .b(N177), .O(N326) );
or2 gate39( .a(N171), .b(N177), .O(N327) );
nand2 gate40( .a(N183), .b(N189), .O(N328) );
or2 gate41( .a(N183), .b(N189), .O(N329) );

  xor2  gate538(.a(N201), .b(N195), .O(gate42inter0));
  nand2 gate539(.a(gate42inter0), .b(s_22), .O(gate42inter1));
  and2  gate540(.a(N201), .b(N195), .O(gate42inter2));
  inv1  gate541(.a(s_22), .O(gate42inter3));
  inv1  gate542(.a(s_23), .O(gate42inter4));
  nand2 gate543(.a(gate42inter4), .b(gate42inter3), .O(gate42inter5));
  nor2  gate544(.a(gate42inter5), .b(gate42inter2), .O(gate42inter6));
  inv1  gate545(.a(N195), .O(gate42inter7));
  inv1  gate546(.a(N201), .O(gate42inter8));
  nand2 gate547(.a(gate42inter8), .b(gate42inter7), .O(gate42inter9));
  nand2 gate548(.a(s_23), .b(gate42inter3), .O(gate42inter10));
  nor2  gate549(.a(gate42inter10), .b(gate42inter9), .O(gate42inter11));
  nor2  gate550(.a(gate42inter11), .b(gate42inter6), .O(gate42inter12));
  nand2 gate551(.a(gate42inter12), .b(gate42inter1), .O(N330));
or2 gate43( .a(N195), .b(N201), .O(N331) );
and2 gate44( .a(N210), .b(N91), .O(N332) );
and2 gate45( .a(N210), .b(N96), .O(N333) );
and2 gate46( .a(N210), .b(N101), .O(N334) );
and2 gate47( .a(N210), .b(N106), .O(N335) );
and2 gate48( .a(N210), .b(N111), .O(N336) );
and2 gate49( .a(N255), .b(N259), .O(N337) );
and2 gate50( .a(N210), .b(N116), .O(N338) );
and2 gate51( .a(N255), .b(N260), .O(N339) );
and2 gate52( .a(N210), .b(N121), .O(N340) );
and2 gate53( .a(N255), .b(N267), .O(N341) );
inv1 gate54( .a(N269), .O(N342) );
inv1 gate55( .a(N273), .O(N343) );
or2 gate56( .a(N270), .b(N273), .O(N344) );
inv1 gate57( .a(N276), .O(N345) );
inv1 gate58( .a(N276), .O(N346) );
inv1 gate59( .a(N279), .O(N347) );
nor2 gate60( .a(N280), .b(N284), .O(N348) );
or2 gate61( .a(N280), .b(N285), .O(N349) );
or2 gate62( .a(N280), .b(N286), .O(N350) );
inv1 gate63( .a(N293), .O(N351) );
inv1 gate64( .a(N294), .O(N352) );
inv1 gate65( .a(N295), .O(N353) );
inv1 gate66( .a(N296), .O(N354) );
nand2 gate67( .a(N89), .b(N298), .O(N355) );
and2 gate68( .a(N90), .b(N298), .O(N356) );

  xor2  gate398(.a(N302), .b(N301), .O(gate69inter0));
  nand2 gate399(.a(gate69inter0), .b(s_2), .O(gate69inter1));
  and2  gate400(.a(N302), .b(N301), .O(gate69inter2));
  inv1  gate401(.a(s_2), .O(gate69inter3));
  inv1  gate402(.a(s_3), .O(gate69inter4));
  nand2 gate403(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate404(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate405(.a(N301), .O(gate69inter7));
  inv1  gate406(.a(N302), .O(gate69inter8));
  nand2 gate407(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate408(.a(s_3), .b(gate69inter3), .O(gate69inter10));
  nor2  gate409(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate410(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate411(.a(gate69inter12), .b(gate69inter1), .O(N357));

  xor2  gate692(.a(N304), .b(N303), .O(gate70inter0));
  nand2 gate693(.a(gate70inter0), .b(s_44), .O(gate70inter1));
  and2  gate694(.a(N304), .b(N303), .O(gate70inter2));
  inv1  gate695(.a(s_44), .O(gate70inter3));
  inv1  gate696(.a(s_45), .O(gate70inter4));
  nand2 gate697(.a(gate70inter4), .b(gate70inter3), .O(gate70inter5));
  nor2  gate698(.a(gate70inter5), .b(gate70inter2), .O(gate70inter6));
  inv1  gate699(.a(N303), .O(gate70inter7));
  inv1  gate700(.a(N304), .O(gate70inter8));
  nand2 gate701(.a(gate70inter8), .b(gate70inter7), .O(gate70inter9));
  nand2 gate702(.a(s_45), .b(gate70inter3), .O(gate70inter10));
  nor2  gate703(.a(gate70inter10), .b(gate70inter9), .O(gate70inter11));
  nor2  gate704(.a(gate70inter11), .b(gate70inter6), .O(gate70inter12));
  nand2 gate705(.a(gate70inter12), .b(gate70inter1), .O(N360));

  xor2  gate664(.a(N306), .b(N305), .O(gate71inter0));
  nand2 gate665(.a(gate71inter0), .b(s_40), .O(gate71inter1));
  and2  gate666(.a(N306), .b(N305), .O(gate71inter2));
  inv1  gate667(.a(s_40), .O(gate71inter3));
  inv1  gate668(.a(s_41), .O(gate71inter4));
  nand2 gate669(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate670(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate671(.a(N305), .O(gate71inter7));
  inv1  gate672(.a(N306), .O(gate71inter8));
  nand2 gate673(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate674(.a(s_41), .b(gate71inter3), .O(gate71inter10));
  nor2  gate675(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate676(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate677(.a(gate71inter12), .b(gate71inter1), .O(N363));
nand2 gate72( .a(N307), .b(N308), .O(N366) );
inv1 gate73( .a(N310), .O(N369) );
nor2 gate74( .a(N322), .b(N323), .O(N375) );
nand2 gate75( .a(N324), .b(N325), .O(N376) );
nand2 gate76( .a(N326), .b(N327), .O(N379) );
nand2 gate77( .a(N328), .b(N329), .O(N382) );
nand2 gate78( .a(N330), .b(N331), .O(N385) );
buf1 gate79( .a(N290), .O(N388) );
buf1 gate80( .a(N291), .O(N389) );
buf1 gate81( .a(N292), .O(N390) );
buf1 gate82( .a(N297), .O(N391) );
or2 gate83( .a(N270), .b(N343), .O(N392) );
inv1 gate84( .a(N345), .O(N393) );
inv1 gate85( .a(N346), .O(N399) );
and2 gate86( .a(N348), .b(N73), .O(N400) );
inv1 gate87( .a(N349), .O(N401) );
inv1 gate88( .a(N350), .O(N402) );
inv1 gate89( .a(N355), .O(N403) );
inv1 gate90( .a(N357), .O(N404) );
inv1 gate91( .a(N360), .O(N405) );
and2 gate92( .a(N357), .b(N360), .O(N406) );
inv1 gate93( .a(N363), .O(N407) );
inv1 gate94( .a(N366), .O(N408) );
and2 gate95( .a(N363), .b(N366), .O(N409) );
nand2 gate96( .a(N347), .b(N352), .O(N410) );
inv1 gate97( .a(N376), .O(N411) );
inv1 gate98( .a(N379), .O(N412) );
and2 gate99( .a(N376), .b(N379), .O(N413) );
inv1 gate100( .a(N382), .O(N414) );
inv1 gate101( .a(N385), .O(N415) );
and2 gate102( .a(N382), .b(N385), .O(N416) );
and2 gate103( .a(N210), .b(N369), .O(N417) );
buf1 gate104( .a(N342), .O(N418) );
buf1 gate105( .a(N344), .O(N419) );
buf1 gate106( .a(N351), .O(N420) );
buf1 gate107( .a(N353), .O(N421) );
buf1 gate108( .a(N354), .O(N422) );
buf1 gate109( .a(N356), .O(N423) );
inv1 gate110( .a(N400), .O(N424) );
and2 gate111( .a(N404), .b(N405), .O(N425) );
and2 gate112( .a(N407), .b(N408), .O(N426) );
and3 gate113( .a(N319), .b(N393), .c(N55), .O(N427) );
and3 gate114( .a(N393), .b(N17), .c(N287), .O(N432) );
nand3 gate115( .a(N393), .b(N287), .c(N55), .O(N437) );
nand4 gate116( .a(N375), .b(N59), .c(N156), .d(N393), .O(N442) );
nand3 gate117( .a(N393), .b(N319), .c(N17), .O(N443) );
and2 gate118( .a(N411), .b(N412), .O(N444) );
and2 gate119( .a(N414), .b(N415), .O(N445) );
buf1 gate120( .a(N392), .O(N446) );
buf1 gate121( .a(N399), .O(N447) );
buf1 gate122( .a(N401), .O(N448) );
buf1 gate123( .a(N402), .O(N449) );
buf1 gate124( .a(N403), .O(N450) );
inv1 gate125( .a(N424), .O(N451) );
nor2 gate126( .a(N406), .b(N425), .O(N460) );
nor2 gate127( .a(N409), .b(N426), .O(N463) );

  xor2  gate748(.a(N410), .b(N442), .O(gate128inter0));
  nand2 gate749(.a(gate128inter0), .b(s_52), .O(gate128inter1));
  and2  gate750(.a(N410), .b(N442), .O(gate128inter2));
  inv1  gate751(.a(s_52), .O(gate128inter3));
  inv1  gate752(.a(s_53), .O(gate128inter4));
  nand2 gate753(.a(gate128inter4), .b(gate128inter3), .O(gate128inter5));
  nor2  gate754(.a(gate128inter5), .b(gate128inter2), .O(gate128inter6));
  inv1  gate755(.a(N442), .O(gate128inter7));
  inv1  gate756(.a(N410), .O(gate128inter8));
  nand2 gate757(.a(gate128inter8), .b(gate128inter7), .O(gate128inter9));
  nand2 gate758(.a(s_53), .b(gate128inter3), .O(gate128inter10));
  nor2  gate759(.a(gate128inter10), .b(gate128inter9), .O(gate128inter11));
  nor2  gate760(.a(gate128inter11), .b(gate128inter6), .O(gate128inter12));
  nand2 gate761(.a(gate128inter12), .b(gate128inter1), .O(N466));
and2 gate129( .a(N143), .b(N427), .O(N475) );
and2 gate130( .a(N310), .b(N432), .O(N476) );
and2 gate131( .a(N146), .b(N427), .O(N477) );
and2 gate132( .a(N310), .b(N432), .O(N478) );
and2 gate133( .a(N149), .b(N427), .O(N479) );
and2 gate134( .a(N310), .b(N432), .O(N480) );
and2 gate135( .a(N153), .b(N427), .O(N481) );
and2 gate136( .a(N310), .b(N432), .O(N482) );

  xor2  gate510(.a(N1), .b(N443), .O(gate137inter0));
  nand2 gate511(.a(gate137inter0), .b(s_18), .O(gate137inter1));
  and2  gate512(.a(N1), .b(N443), .O(gate137inter2));
  inv1  gate513(.a(s_18), .O(gate137inter3));
  inv1  gate514(.a(s_19), .O(gate137inter4));
  nand2 gate515(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate516(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate517(.a(N443), .O(gate137inter7));
  inv1  gate518(.a(N1), .O(gate137inter8));
  nand2 gate519(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate520(.a(s_19), .b(gate137inter3), .O(gate137inter10));
  nor2  gate521(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate522(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate523(.a(gate137inter12), .b(gate137inter1), .O(N483));
or2 gate138( .a(N369), .b(N437), .O(N488) );
or2 gate139( .a(N369), .b(N437), .O(N489) );
or2 gate140( .a(N369), .b(N437), .O(N490) );
or2 gate141( .a(N369), .b(N437), .O(N491) );
nor2 gate142( .a(N413), .b(N444), .O(N492) );
nor2 gate143( .a(N416), .b(N445), .O(N495) );

  xor2  gate804(.a(N460), .b(N130), .O(gate144inter0));
  nand2 gate805(.a(gate144inter0), .b(s_60), .O(gate144inter1));
  and2  gate806(.a(N460), .b(N130), .O(gate144inter2));
  inv1  gate807(.a(s_60), .O(gate144inter3));
  inv1  gate808(.a(s_61), .O(gate144inter4));
  nand2 gate809(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate810(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate811(.a(N130), .O(gate144inter7));
  inv1  gate812(.a(N460), .O(gate144inter8));
  nand2 gate813(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate814(.a(s_61), .b(gate144inter3), .O(gate144inter10));
  nor2  gate815(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate816(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate817(.a(gate144inter12), .b(gate144inter1), .O(N498));
or2 gate145( .a(N130), .b(N460), .O(N499) );
nand2 gate146( .a(N463), .b(N135), .O(N500) );
or2 gate147( .a(N463), .b(N135), .O(N501) );
and2 gate148( .a(N91), .b(N466), .O(N502) );

  xor2  gate832(.a(N476), .b(N475), .O(gate149inter0));
  nand2 gate833(.a(gate149inter0), .b(s_64), .O(gate149inter1));
  and2  gate834(.a(N476), .b(N475), .O(gate149inter2));
  inv1  gate835(.a(s_64), .O(gate149inter3));
  inv1  gate836(.a(s_65), .O(gate149inter4));
  nand2 gate837(.a(gate149inter4), .b(gate149inter3), .O(gate149inter5));
  nor2  gate838(.a(gate149inter5), .b(gate149inter2), .O(gate149inter6));
  inv1  gate839(.a(N475), .O(gate149inter7));
  inv1  gate840(.a(N476), .O(gate149inter8));
  nand2 gate841(.a(gate149inter8), .b(gate149inter7), .O(gate149inter9));
  nand2 gate842(.a(s_65), .b(gate149inter3), .O(gate149inter10));
  nor2  gate843(.a(gate149inter10), .b(gate149inter9), .O(gate149inter11));
  nor2  gate844(.a(gate149inter11), .b(gate149inter6), .O(gate149inter12));
  nand2 gate845(.a(gate149inter12), .b(gate149inter1), .O(N503));
and2 gate150( .a(N96), .b(N466), .O(N504) );

  xor2  gate650(.a(N478), .b(N477), .O(gate151inter0));
  nand2 gate651(.a(gate151inter0), .b(s_38), .O(gate151inter1));
  and2  gate652(.a(N478), .b(N477), .O(gate151inter2));
  inv1  gate653(.a(s_38), .O(gate151inter3));
  inv1  gate654(.a(s_39), .O(gate151inter4));
  nand2 gate655(.a(gate151inter4), .b(gate151inter3), .O(gate151inter5));
  nor2  gate656(.a(gate151inter5), .b(gate151inter2), .O(gate151inter6));
  inv1  gate657(.a(N477), .O(gate151inter7));
  inv1  gate658(.a(N478), .O(gate151inter8));
  nand2 gate659(.a(gate151inter8), .b(gate151inter7), .O(gate151inter9));
  nand2 gate660(.a(s_39), .b(gate151inter3), .O(gate151inter10));
  nor2  gate661(.a(gate151inter10), .b(gate151inter9), .O(gate151inter11));
  nor2  gate662(.a(gate151inter11), .b(gate151inter6), .O(gate151inter12));
  nand2 gate663(.a(gate151inter12), .b(gate151inter1), .O(N505));
and2 gate152( .a(N101), .b(N466), .O(N506) );

  xor2  gate888(.a(N480), .b(N479), .O(gate153inter0));
  nand2 gate889(.a(gate153inter0), .b(s_72), .O(gate153inter1));
  and2  gate890(.a(N480), .b(N479), .O(gate153inter2));
  inv1  gate891(.a(s_72), .O(gate153inter3));
  inv1  gate892(.a(s_73), .O(gate153inter4));
  nand2 gate893(.a(gate153inter4), .b(gate153inter3), .O(gate153inter5));
  nor2  gate894(.a(gate153inter5), .b(gate153inter2), .O(gate153inter6));
  inv1  gate895(.a(N479), .O(gate153inter7));
  inv1  gate896(.a(N480), .O(gate153inter8));
  nand2 gate897(.a(gate153inter8), .b(gate153inter7), .O(gate153inter9));
  nand2 gate898(.a(s_73), .b(gate153inter3), .O(gate153inter10));
  nor2  gate899(.a(gate153inter10), .b(gate153inter9), .O(gate153inter11));
  nor2  gate900(.a(gate153inter11), .b(gate153inter6), .O(gate153inter12));
  nand2 gate901(.a(gate153inter12), .b(gate153inter1), .O(N507));
and2 gate154( .a(N106), .b(N466), .O(N508) );

  xor2  gate790(.a(N482), .b(N481), .O(gate155inter0));
  nand2 gate791(.a(gate155inter0), .b(s_58), .O(gate155inter1));
  and2  gate792(.a(N482), .b(N481), .O(gate155inter2));
  inv1  gate793(.a(s_58), .O(gate155inter3));
  inv1  gate794(.a(s_59), .O(gate155inter4));
  nand2 gate795(.a(gate155inter4), .b(gate155inter3), .O(gate155inter5));
  nor2  gate796(.a(gate155inter5), .b(gate155inter2), .O(gate155inter6));
  inv1  gate797(.a(N481), .O(gate155inter7));
  inv1  gate798(.a(N482), .O(gate155inter8));
  nand2 gate799(.a(gate155inter8), .b(gate155inter7), .O(gate155inter9));
  nand2 gate800(.a(s_59), .b(gate155inter3), .O(gate155inter10));
  nor2  gate801(.a(gate155inter10), .b(gate155inter9), .O(gate155inter11));
  nor2  gate802(.a(gate155inter11), .b(gate155inter6), .O(gate155inter12));
  nand2 gate803(.a(gate155inter12), .b(gate155inter1), .O(N509));
and2 gate156( .a(N143), .b(N483), .O(N510) );
and2 gate157( .a(N111), .b(N466), .O(N511) );
and2 gate158( .a(N146), .b(N483), .O(N512) );
and2 gate159( .a(N116), .b(N466), .O(N513) );
and2 gate160( .a(N149), .b(N483), .O(N514) );
and2 gate161( .a(N121), .b(N466), .O(N515) );
and2 gate162( .a(N153), .b(N483), .O(N516) );
and2 gate163( .a(N126), .b(N466), .O(N517) );
nand2 gate164( .a(N130), .b(N492), .O(N518) );
or2 gate165( .a(N130), .b(N492), .O(N519) );

  xor2  gate874(.a(N207), .b(N495), .O(gate166inter0));
  nand2 gate875(.a(gate166inter0), .b(s_70), .O(gate166inter1));
  and2  gate876(.a(N207), .b(N495), .O(gate166inter2));
  inv1  gate877(.a(s_70), .O(gate166inter3));
  inv1  gate878(.a(s_71), .O(gate166inter4));
  nand2 gate879(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate880(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate881(.a(N495), .O(gate166inter7));
  inv1  gate882(.a(N207), .O(gate166inter8));
  nand2 gate883(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate884(.a(s_71), .b(gate166inter3), .O(gate166inter10));
  nor2  gate885(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate886(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate887(.a(gate166inter12), .b(gate166inter1), .O(N520));
or2 gate167( .a(N495), .b(N207), .O(N521) );
and2 gate168( .a(N451), .b(N159), .O(N522) );
and2 gate169( .a(N451), .b(N165), .O(N523) );
and2 gate170( .a(N451), .b(N171), .O(N524) );
and2 gate171( .a(N451), .b(N177), .O(N525) );
and2 gate172( .a(N451), .b(N183), .O(N526) );
nand2 gate173( .a(N451), .b(N189), .O(N527) );

  xor2  gate944(.a(N195), .b(N451), .O(gate174inter0));
  nand2 gate945(.a(gate174inter0), .b(s_80), .O(gate174inter1));
  and2  gate946(.a(N195), .b(N451), .O(gate174inter2));
  inv1  gate947(.a(s_80), .O(gate174inter3));
  inv1  gate948(.a(s_81), .O(gate174inter4));
  nand2 gate949(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate950(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate951(.a(N451), .O(gate174inter7));
  inv1  gate952(.a(N195), .O(gate174inter8));
  nand2 gate953(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate954(.a(s_81), .b(gate174inter3), .O(gate174inter10));
  nor2  gate955(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate956(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate957(.a(gate174inter12), .b(gate174inter1), .O(N528));
nand2 gate175( .a(N451), .b(N201), .O(N529) );
nand2 gate176( .a(N498), .b(N499), .O(N530) );

  xor2  gate860(.a(N501), .b(N500), .O(gate177inter0));
  nand2 gate861(.a(gate177inter0), .b(s_68), .O(gate177inter1));
  and2  gate862(.a(N501), .b(N500), .O(gate177inter2));
  inv1  gate863(.a(s_68), .O(gate177inter3));
  inv1  gate864(.a(s_69), .O(gate177inter4));
  nand2 gate865(.a(gate177inter4), .b(gate177inter3), .O(gate177inter5));
  nor2  gate866(.a(gate177inter5), .b(gate177inter2), .O(gate177inter6));
  inv1  gate867(.a(N500), .O(gate177inter7));
  inv1  gate868(.a(N501), .O(gate177inter8));
  nand2 gate869(.a(gate177inter8), .b(gate177inter7), .O(gate177inter9));
  nand2 gate870(.a(s_69), .b(gate177inter3), .O(gate177inter10));
  nor2  gate871(.a(gate177inter10), .b(gate177inter9), .O(gate177inter11));
  nor2  gate872(.a(gate177inter11), .b(gate177inter6), .O(gate177inter12));
  nand2 gate873(.a(gate177inter12), .b(gate177inter1), .O(N533));
nor2 gate178( .a(N309), .b(N502), .O(N536) );
nor2 gate179( .a(N316), .b(N504), .O(N537) );

  xor2  gate384(.a(N506), .b(N317), .O(gate180inter0));
  nand2 gate385(.a(gate180inter0), .b(s_0), .O(gate180inter1));
  and2  gate386(.a(N506), .b(N317), .O(gate180inter2));
  inv1  gate387(.a(s_0), .O(gate180inter3));
  inv1  gate388(.a(s_1), .O(gate180inter4));
  nand2 gate389(.a(gate180inter4), .b(gate180inter3), .O(gate180inter5));
  nor2  gate390(.a(gate180inter5), .b(gate180inter2), .O(gate180inter6));
  inv1  gate391(.a(N317), .O(gate180inter7));
  inv1  gate392(.a(N506), .O(gate180inter8));
  nand2 gate393(.a(gate180inter8), .b(gate180inter7), .O(gate180inter9));
  nand2 gate394(.a(s_1), .b(gate180inter3), .O(gate180inter10));
  nor2  gate395(.a(gate180inter10), .b(gate180inter9), .O(gate180inter11));
  nor2  gate396(.a(gate180inter11), .b(gate180inter6), .O(gate180inter12));
  nand2 gate397(.a(gate180inter12), .b(gate180inter1), .O(N538));

  xor2  gate454(.a(N508), .b(N318), .O(gate181inter0));
  nand2 gate455(.a(gate181inter0), .b(s_10), .O(gate181inter1));
  and2  gate456(.a(N508), .b(N318), .O(gate181inter2));
  inv1  gate457(.a(s_10), .O(gate181inter3));
  inv1  gate458(.a(s_11), .O(gate181inter4));
  nand2 gate459(.a(gate181inter4), .b(gate181inter3), .O(gate181inter5));
  nor2  gate460(.a(gate181inter5), .b(gate181inter2), .O(gate181inter6));
  inv1  gate461(.a(N318), .O(gate181inter7));
  inv1  gate462(.a(N508), .O(gate181inter8));
  nand2 gate463(.a(gate181inter8), .b(gate181inter7), .O(gate181inter9));
  nand2 gate464(.a(s_11), .b(gate181inter3), .O(gate181inter10));
  nor2  gate465(.a(gate181inter10), .b(gate181inter9), .O(gate181inter11));
  nor2  gate466(.a(gate181inter11), .b(gate181inter6), .O(gate181inter12));
  nand2 gate467(.a(gate181inter12), .b(gate181inter1), .O(N539));
nor2 gate182( .a(N510), .b(N511), .O(N540) );

  xor2  gate608(.a(N513), .b(N512), .O(gate183inter0));
  nand2 gate609(.a(gate183inter0), .b(s_32), .O(gate183inter1));
  and2  gate610(.a(N513), .b(N512), .O(gate183inter2));
  inv1  gate611(.a(s_32), .O(gate183inter3));
  inv1  gate612(.a(s_33), .O(gate183inter4));
  nand2 gate613(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate614(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate615(.a(N512), .O(gate183inter7));
  inv1  gate616(.a(N513), .O(gate183inter8));
  nand2 gate617(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate618(.a(s_33), .b(gate183inter3), .O(gate183inter10));
  nor2  gate619(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate620(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate621(.a(gate183inter12), .b(gate183inter1), .O(N541));

  xor2  gate496(.a(N515), .b(N514), .O(gate184inter0));
  nand2 gate497(.a(gate184inter0), .b(s_16), .O(gate184inter1));
  and2  gate498(.a(N515), .b(N514), .O(gate184inter2));
  inv1  gate499(.a(s_16), .O(gate184inter3));
  inv1  gate500(.a(s_17), .O(gate184inter4));
  nand2 gate501(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate502(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate503(.a(N514), .O(gate184inter7));
  inv1  gate504(.a(N515), .O(gate184inter8));
  nand2 gate505(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate506(.a(s_17), .b(gate184inter3), .O(gate184inter10));
  nor2  gate507(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate508(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate509(.a(gate184inter12), .b(gate184inter1), .O(N542));
nor2 gate185( .a(N516), .b(N517), .O(N543) );

  xor2  gate706(.a(N519), .b(N518), .O(gate186inter0));
  nand2 gate707(.a(gate186inter0), .b(s_46), .O(gate186inter1));
  and2  gate708(.a(N519), .b(N518), .O(gate186inter2));
  inv1  gate709(.a(s_46), .O(gate186inter3));
  inv1  gate710(.a(s_47), .O(gate186inter4));
  nand2 gate711(.a(gate186inter4), .b(gate186inter3), .O(gate186inter5));
  nor2  gate712(.a(gate186inter5), .b(gate186inter2), .O(gate186inter6));
  inv1  gate713(.a(N518), .O(gate186inter7));
  inv1  gate714(.a(N519), .O(gate186inter8));
  nand2 gate715(.a(gate186inter8), .b(gate186inter7), .O(gate186inter9));
  nand2 gate716(.a(s_47), .b(gate186inter3), .O(gate186inter10));
  nor2  gate717(.a(gate186inter10), .b(gate186inter9), .O(gate186inter11));
  nor2  gate718(.a(gate186inter11), .b(gate186inter6), .O(gate186inter12));
  nand2 gate719(.a(gate186inter12), .b(gate186inter1), .O(N544));
nand2 gate187( .a(N520), .b(N521), .O(N547) );
inv1 gate188( .a(N530), .O(N550) );
inv1 gate189( .a(N533), .O(N551) );
and2 gate190( .a(N530), .b(N533), .O(N552) );

  xor2  gate776(.a(N503), .b(N536), .O(gate191inter0));
  nand2 gate777(.a(gate191inter0), .b(s_56), .O(gate191inter1));
  and2  gate778(.a(N503), .b(N536), .O(gate191inter2));
  inv1  gate779(.a(s_56), .O(gate191inter3));
  inv1  gate780(.a(s_57), .O(gate191inter4));
  nand2 gate781(.a(gate191inter4), .b(gate191inter3), .O(gate191inter5));
  nor2  gate782(.a(gate191inter5), .b(gate191inter2), .O(gate191inter6));
  inv1  gate783(.a(N536), .O(gate191inter7));
  inv1  gate784(.a(N503), .O(gate191inter8));
  nand2 gate785(.a(gate191inter8), .b(gate191inter7), .O(gate191inter9));
  nand2 gate786(.a(s_57), .b(gate191inter3), .O(gate191inter10));
  nor2  gate787(.a(gate191inter10), .b(gate191inter9), .O(gate191inter11));
  nor2  gate788(.a(gate191inter11), .b(gate191inter6), .O(gate191inter12));
  nand2 gate789(.a(gate191inter12), .b(gate191inter1), .O(N553));

  xor2  gate622(.a(N505), .b(N537), .O(gate192inter0));
  nand2 gate623(.a(gate192inter0), .b(s_34), .O(gate192inter1));
  and2  gate624(.a(N505), .b(N537), .O(gate192inter2));
  inv1  gate625(.a(s_34), .O(gate192inter3));
  inv1  gate626(.a(s_35), .O(gate192inter4));
  nand2 gate627(.a(gate192inter4), .b(gate192inter3), .O(gate192inter5));
  nor2  gate628(.a(gate192inter5), .b(gate192inter2), .O(gate192inter6));
  inv1  gate629(.a(N537), .O(gate192inter7));
  inv1  gate630(.a(N505), .O(gate192inter8));
  nand2 gate631(.a(gate192inter8), .b(gate192inter7), .O(gate192inter9));
  nand2 gate632(.a(s_35), .b(gate192inter3), .O(gate192inter10));
  nor2  gate633(.a(gate192inter10), .b(gate192inter9), .O(gate192inter11));
  nor2  gate634(.a(gate192inter11), .b(gate192inter6), .O(gate192inter12));
  nand2 gate635(.a(gate192inter12), .b(gate192inter1), .O(N557));
nand2 gate193( .a(N538), .b(N507), .O(N561) );
nand2 gate194( .a(N539), .b(N509), .O(N565) );
nand2 gate195( .a(N488), .b(N540), .O(N569) );
nand2 gate196( .a(N489), .b(N541), .O(N573) );

  xor2  gate916(.a(N542), .b(N490), .O(gate197inter0));
  nand2 gate917(.a(gate197inter0), .b(s_76), .O(gate197inter1));
  and2  gate918(.a(N542), .b(N490), .O(gate197inter2));
  inv1  gate919(.a(s_76), .O(gate197inter3));
  inv1  gate920(.a(s_77), .O(gate197inter4));
  nand2 gate921(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate922(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate923(.a(N490), .O(gate197inter7));
  inv1  gate924(.a(N542), .O(gate197inter8));
  nand2 gate925(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate926(.a(s_77), .b(gate197inter3), .O(gate197inter10));
  nor2  gate927(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate928(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate929(.a(gate197inter12), .b(gate197inter1), .O(N577));
nand2 gate198( .a(N491), .b(N543), .O(N581) );
inv1 gate199( .a(N544), .O(N585) );
inv1 gate200( .a(N547), .O(N586) );
and2 gate201( .a(N544), .b(N547), .O(N587) );
and2 gate202( .a(N550), .b(N551), .O(N588) );
and2 gate203( .a(N585), .b(N586), .O(N589) );
nand2 gate204( .a(N553), .b(N159), .O(N590) );
or2 gate205( .a(N553), .b(N159), .O(N593) );
and2 gate206( .a(N246), .b(N553), .O(N596) );
nand2 gate207( .a(N557), .b(N165), .O(N597) );
or2 gate208( .a(N557), .b(N165), .O(N600) );
and2 gate209( .a(N246), .b(N557), .O(N605) );
nand2 gate210( .a(N561), .b(N171), .O(N606) );
or2 gate211( .a(N561), .b(N171), .O(N609) );
and2 gate212( .a(N246), .b(N561), .O(N615) );
nand2 gate213( .a(N565), .b(N177), .O(N616) );
or2 gate214( .a(N565), .b(N177), .O(N619) );
and2 gate215( .a(N246), .b(N565), .O(N624) );

  xor2  gate552(.a(N183), .b(N569), .O(gate216inter0));
  nand2 gate553(.a(gate216inter0), .b(s_24), .O(gate216inter1));
  and2  gate554(.a(N183), .b(N569), .O(gate216inter2));
  inv1  gate555(.a(s_24), .O(gate216inter3));
  inv1  gate556(.a(s_25), .O(gate216inter4));
  nand2 gate557(.a(gate216inter4), .b(gate216inter3), .O(gate216inter5));
  nor2  gate558(.a(gate216inter5), .b(gate216inter2), .O(gate216inter6));
  inv1  gate559(.a(N569), .O(gate216inter7));
  inv1  gate560(.a(N183), .O(gate216inter8));
  nand2 gate561(.a(gate216inter8), .b(gate216inter7), .O(gate216inter9));
  nand2 gate562(.a(s_25), .b(gate216inter3), .O(gate216inter10));
  nor2  gate563(.a(gate216inter10), .b(gate216inter9), .O(gate216inter11));
  nor2  gate564(.a(gate216inter11), .b(gate216inter6), .O(gate216inter12));
  nand2 gate565(.a(gate216inter12), .b(gate216inter1), .O(N625));
or2 gate217( .a(N569), .b(N183), .O(N628) );
and2 gate218( .a(N246), .b(N569), .O(N631) );
nand2 gate219( .a(N573), .b(N189), .O(N632) );
or2 gate220( .a(N573), .b(N189), .O(N635) );
and2 gate221( .a(N246), .b(N573), .O(N640) );
nand2 gate222( .a(N577), .b(N195), .O(N641) );
or2 gate223( .a(N577), .b(N195), .O(N644) );
and2 gate224( .a(N246), .b(N577), .O(N650) );

  xor2  gate930(.a(N201), .b(N581), .O(gate225inter0));
  nand2 gate931(.a(gate225inter0), .b(s_78), .O(gate225inter1));
  and2  gate932(.a(N201), .b(N581), .O(gate225inter2));
  inv1  gate933(.a(s_78), .O(gate225inter3));
  inv1  gate934(.a(s_79), .O(gate225inter4));
  nand2 gate935(.a(gate225inter4), .b(gate225inter3), .O(gate225inter5));
  nor2  gate936(.a(gate225inter5), .b(gate225inter2), .O(gate225inter6));
  inv1  gate937(.a(N581), .O(gate225inter7));
  inv1  gate938(.a(N201), .O(gate225inter8));
  nand2 gate939(.a(gate225inter8), .b(gate225inter7), .O(gate225inter9));
  nand2 gate940(.a(s_79), .b(gate225inter3), .O(gate225inter10));
  nor2  gate941(.a(gate225inter10), .b(gate225inter9), .O(gate225inter11));
  nor2  gate942(.a(gate225inter11), .b(gate225inter6), .O(gate225inter12));
  nand2 gate943(.a(gate225inter12), .b(gate225inter1), .O(N651));
or2 gate226( .a(N581), .b(N201), .O(N654) );
and2 gate227( .a(N246), .b(N581), .O(N659) );
nor2 gate228( .a(N552), .b(N588), .O(N660) );
nor2 gate229( .a(N587), .b(N589), .O(N661) );
inv1 gate230( .a(N590), .O(N662) );
and2 gate231( .a(N593), .b(N590), .O(N665) );

  xor2  gate818(.a(N522), .b(N596), .O(gate232inter0));
  nand2 gate819(.a(gate232inter0), .b(s_62), .O(gate232inter1));
  and2  gate820(.a(N522), .b(N596), .O(gate232inter2));
  inv1  gate821(.a(s_62), .O(gate232inter3));
  inv1  gate822(.a(s_63), .O(gate232inter4));
  nand2 gate823(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate824(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate825(.a(N596), .O(gate232inter7));
  inv1  gate826(.a(N522), .O(gate232inter8));
  nand2 gate827(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate828(.a(s_63), .b(gate232inter3), .O(gate232inter10));
  nor2  gate829(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate830(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate831(.a(gate232inter12), .b(gate232inter1), .O(N669));
inv1 gate233( .a(N597), .O(N670) );
and2 gate234( .a(N600), .b(N597), .O(N673) );

  xor2  gate524(.a(N523), .b(N605), .O(gate235inter0));
  nand2 gate525(.a(gate235inter0), .b(s_20), .O(gate235inter1));
  and2  gate526(.a(N523), .b(N605), .O(gate235inter2));
  inv1  gate527(.a(s_20), .O(gate235inter3));
  inv1  gate528(.a(s_21), .O(gate235inter4));
  nand2 gate529(.a(gate235inter4), .b(gate235inter3), .O(gate235inter5));
  nor2  gate530(.a(gate235inter5), .b(gate235inter2), .O(gate235inter6));
  inv1  gate531(.a(N605), .O(gate235inter7));
  inv1  gate532(.a(N523), .O(gate235inter8));
  nand2 gate533(.a(gate235inter8), .b(gate235inter7), .O(gate235inter9));
  nand2 gate534(.a(s_21), .b(gate235inter3), .O(gate235inter10));
  nor2  gate535(.a(gate235inter10), .b(gate235inter9), .O(gate235inter11));
  nor2  gate536(.a(gate235inter11), .b(gate235inter6), .O(gate235inter12));
  nand2 gate537(.a(gate235inter12), .b(gate235inter1), .O(N677));
inv1 gate236( .a(N606), .O(N678) );
and2 gate237( .a(N609), .b(N606), .O(N682) );

  xor2  gate426(.a(N524), .b(N615), .O(gate238inter0));
  nand2 gate427(.a(gate238inter0), .b(s_6), .O(gate238inter1));
  and2  gate428(.a(N524), .b(N615), .O(gate238inter2));
  inv1  gate429(.a(s_6), .O(gate238inter3));
  inv1  gate430(.a(s_7), .O(gate238inter4));
  nand2 gate431(.a(gate238inter4), .b(gate238inter3), .O(gate238inter5));
  nor2  gate432(.a(gate238inter5), .b(gate238inter2), .O(gate238inter6));
  inv1  gate433(.a(N615), .O(gate238inter7));
  inv1  gate434(.a(N524), .O(gate238inter8));
  nand2 gate435(.a(gate238inter8), .b(gate238inter7), .O(gate238inter9));
  nand2 gate436(.a(s_7), .b(gate238inter3), .O(gate238inter10));
  nor2  gate437(.a(gate238inter10), .b(gate238inter9), .O(gate238inter11));
  nor2  gate438(.a(gate238inter11), .b(gate238inter6), .O(gate238inter12));
  nand2 gate439(.a(gate238inter12), .b(gate238inter1), .O(N686));
inv1 gate239( .a(N616), .O(N687) );
and2 gate240( .a(N619), .b(N616), .O(N692) );
nor2 gate241( .a(N624), .b(N525), .O(N696) );
inv1 gate242( .a(N625), .O(N697) );
and2 gate243( .a(N628), .b(N625), .O(N700) );

  xor2  gate412(.a(N526), .b(N631), .O(gate244inter0));
  nand2 gate413(.a(gate244inter0), .b(s_4), .O(gate244inter1));
  and2  gate414(.a(N526), .b(N631), .O(gate244inter2));
  inv1  gate415(.a(s_4), .O(gate244inter3));
  inv1  gate416(.a(s_5), .O(gate244inter4));
  nand2 gate417(.a(gate244inter4), .b(gate244inter3), .O(gate244inter5));
  nor2  gate418(.a(gate244inter5), .b(gate244inter2), .O(gate244inter6));
  inv1  gate419(.a(N631), .O(gate244inter7));
  inv1  gate420(.a(N526), .O(gate244inter8));
  nand2 gate421(.a(gate244inter8), .b(gate244inter7), .O(gate244inter9));
  nand2 gate422(.a(s_5), .b(gate244inter3), .O(gate244inter10));
  nor2  gate423(.a(gate244inter10), .b(gate244inter9), .O(gate244inter11));
  nor2  gate424(.a(gate244inter11), .b(gate244inter6), .O(gate244inter12));
  nand2 gate425(.a(gate244inter12), .b(gate244inter1), .O(N704));
inv1 gate245( .a(N632), .O(N705) );
and2 gate246( .a(N635), .b(N632), .O(N708) );
nor2 gate247( .a(N337), .b(N640), .O(N712) );
inv1 gate248( .a(N641), .O(N713) );
and2 gate249( .a(N644), .b(N641), .O(N717) );
nor2 gate250( .a(N339), .b(N650), .O(N721) );
inv1 gate251( .a(N651), .O(N722) );
and2 gate252( .a(N654), .b(N651), .O(N727) );
nor2 gate253( .a(N341), .b(N659), .O(N731) );

  xor2  gate482(.a(N261), .b(N654), .O(gate254inter0));
  nand2 gate483(.a(gate254inter0), .b(s_14), .O(gate254inter1));
  and2  gate484(.a(N261), .b(N654), .O(gate254inter2));
  inv1  gate485(.a(s_14), .O(gate254inter3));
  inv1  gate486(.a(s_15), .O(gate254inter4));
  nand2 gate487(.a(gate254inter4), .b(gate254inter3), .O(gate254inter5));
  nor2  gate488(.a(gate254inter5), .b(gate254inter2), .O(gate254inter6));
  inv1  gate489(.a(N654), .O(gate254inter7));
  inv1  gate490(.a(N261), .O(gate254inter8));
  nand2 gate491(.a(gate254inter8), .b(gate254inter7), .O(gate254inter9));
  nand2 gate492(.a(s_15), .b(gate254inter3), .O(gate254inter10));
  nor2  gate493(.a(gate254inter10), .b(gate254inter9), .O(gate254inter11));
  nor2  gate494(.a(gate254inter11), .b(gate254inter6), .O(gate254inter12));
  nand2 gate495(.a(gate254inter12), .b(gate254inter1), .O(N732));
nand3 gate255( .a(N644), .b(N654), .c(N261), .O(N733) );
nand4 gate256( .a(N635), .b(N644), .c(N654), .d(N261), .O(N734) );
inv1 gate257( .a(N662), .O(N735) );
and2 gate258( .a(N228), .b(N665), .O(N736) );
and2 gate259( .a(N237), .b(N662), .O(N737) );
inv1 gate260( .a(N670), .O(N738) );
and2 gate261( .a(N228), .b(N673), .O(N739) );
and2 gate262( .a(N237), .b(N670), .O(N740) );
inv1 gate263( .a(N678), .O(N741) );
and2 gate264( .a(N228), .b(N682), .O(N742) );
and2 gate265( .a(N237), .b(N678), .O(N743) );
inv1 gate266( .a(N687), .O(N744) );
and2 gate267( .a(N228), .b(N692), .O(N745) );
and2 gate268( .a(N237), .b(N687), .O(N746) );
inv1 gate269( .a(N697), .O(N747) );
and2 gate270( .a(N228), .b(N700), .O(N748) );
and2 gate271( .a(N237), .b(N697), .O(N749) );
inv1 gate272( .a(N705), .O(N750) );
and2 gate273( .a(N228), .b(N708), .O(N751) );
and2 gate274( .a(N237), .b(N705), .O(N752) );
inv1 gate275( .a(N713), .O(N753) );
and2 gate276( .a(N228), .b(N717), .O(N754) );
and2 gate277( .a(N237), .b(N713), .O(N755) );
inv1 gate278( .a(N722), .O(N756) );
nor2 gate279( .a(N727), .b(N261), .O(N757) );
and2 gate280( .a(N727), .b(N261), .O(N758) );
and2 gate281( .a(N228), .b(N727), .O(N759) );
and2 gate282( .a(N237), .b(N722), .O(N760) );
nand2 gate283( .a(N644), .b(N722), .O(N761) );
nand2 gate284( .a(N635), .b(N713), .O(N762) );
nand3 gate285( .a(N635), .b(N644), .c(N722), .O(N763) );
nand2 gate286( .a(N609), .b(N687), .O(N764) );
nand2 gate287( .a(N600), .b(N678), .O(N765) );
nand3 gate288( .a(N600), .b(N609), .c(N687), .O(N766) );
buf1 gate289( .a(N660), .O(N767) );
buf1 gate290( .a(N661), .O(N768) );
nor2 gate291( .a(N736), .b(N737), .O(N769) );

  xor2  gate468(.a(N740), .b(N739), .O(gate292inter0));
  nand2 gate469(.a(gate292inter0), .b(s_12), .O(gate292inter1));
  and2  gate470(.a(N740), .b(N739), .O(gate292inter2));
  inv1  gate471(.a(s_12), .O(gate292inter3));
  inv1  gate472(.a(s_13), .O(gate292inter4));
  nand2 gate473(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate474(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate475(.a(N739), .O(gate292inter7));
  inv1  gate476(.a(N740), .O(gate292inter8));
  nand2 gate477(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate478(.a(s_13), .b(gate292inter3), .O(gate292inter10));
  nor2  gate479(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate480(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate481(.a(gate292inter12), .b(gate292inter1), .O(N770));

  xor2  gate720(.a(N743), .b(N742), .O(gate293inter0));
  nand2 gate721(.a(gate293inter0), .b(s_48), .O(gate293inter1));
  and2  gate722(.a(N743), .b(N742), .O(gate293inter2));
  inv1  gate723(.a(s_48), .O(gate293inter3));
  inv1  gate724(.a(s_49), .O(gate293inter4));
  nand2 gate725(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate726(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate727(.a(N742), .O(gate293inter7));
  inv1  gate728(.a(N743), .O(gate293inter8));
  nand2 gate729(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate730(.a(s_49), .b(gate293inter3), .O(gate293inter10));
  nor2  gate731(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate732(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate733(.a(gate293inter12), .b(gate293inter1), .O(N771));

  xor2  gate580(.a(N746), .b(N745), .O(gate294inter0));
  nand2 gate581(.a(gate294inter0), .b(s_28), .O(gate294inter1));
  and2  gate582(.a(N746), .b(N745), .O(gate294inter2));
  inv1  gate583(.a(s_28), .O(gate294inter3));
  inv1  gate584(.a(s_29), .O(gate294inter4));
  nand2 gate585(.a(gate294inter4), .b(gate294inter3), .O(gate294inter5));
  nor2  gate586(.a(gate294inter5), .b(gate294inter2), .O(gate294inter6));
  inv1  gate587(.a(N745), .O(gate294inter7));
  inv1  gate588(.a(N746), .O(gate294inter8));
  nand2 gate589(.a(gate294inter8), .b(gate294inter7), .O(gate294inter9));
  nand2 gate590(.a(s_29), .b(gate294inter3), .O(gate294inter10));
  nor2  gate591(.a(gate294inter10), .b(gate294inter9), .O(gate294inter11));
  nor2  gate592(.a(gate294inter11), .b(gate294inter6), .O(gate294inter12));
  nand2 gate593(.a(gate294inter12), .b(gate294inter1), .O(N772));
nand4 gate295( .a(N750), .b(N762), .c(N763), .d(N734), .O(N773) );
nor2 gate296( .a(N748), .b(N749), .O(N777) );
nand3 gate297( .a(N753), .b(N761), .c(N733), .O(N778) );
nor2 gate298( .a(N751), .b(N752), .O(N781) );

  xor2  gate902(.a(N732), .b(N756), .O(gate299inter0));
  nand2 gate903(.a(gate299inter0), .b(s_74), .O(gate299inter1));
  and2  gate904(.a(N732), .b(N756), .O(gate299inter2));
  inv1  gate905(.a(s_74), .O(gate299inter3));
  inv1  gate906(.a(s_75), .O(gate299inter4));
  nand2 gate907(.a(gate299inter4), .b(gate299inter3), .O(gate299inter5));
  nor2  gate908(.a(gate299inter5), .b(gate299inter2), .O(gate299inter6));
  inv1  gate909(.a(N756), .O(gate299inter7));
  inv1  gate910(.a(N732), .O(gate299inter8));
  nand2 gate911(.a(gate299inter8), .b(gate299inter7), .O(gate299inter9));
  nand2 gate912(.a(s_75), .b(gate299inter3), .O(gate299inter10));
  nor2  gate913(.a(gate299inter10), .b(gate299inter9), .O(gate299inter11));
  nor2  gate914(.a(gate299inter11), .b(gate299inter6), .O(gate299inter12));
  nand2 gate915(.a(gate299inter12), .b(gate299inter1), .O(N782));
nor2 gate300( .a(N754), .b(N755), .O(N785) );
nor2 gate301( .a(N757), .b(N758), .O(N786) );
nor2 gate302( .a(N759), .b(N760), .O(N787) );
nor2 gate303( .a(N700), .b(N773), .O(N788) );
and2 gate304( .a(N700), .b(N773), .O(N789) );
nor2 gate305( .a(N708), .b(N778), .O(N790) );
and2 gate306( .a(N708), .b(N778), .O(N791) );
nor2 gate307( .a(N717), .b(N782), .O(N792) );
and2 gate308( .a(N717), .b(N782), .O(N793) );
and2 gate309( .a(N219), .b(N786), .O(N794) );

  xor2  gate594(.a(N773), .b(N628), .O(gate310inter0));
  nand2 gate595(.a(gate310inter0), .b(s_30), .O(gate310inter1));
  and2  gate596(.a(N773), .b(N628), .O(gate310inter2));
  inv1  gate597(.a(s_30), .O(gate310inter3));
  inv1  gate598(.a(s_31), .O(gate310inter4));
  nand2 gate599(.a(gate310inter4), .b(gate310inter3), .O(gate310inter5));
  nor2  gate600(.a(gate310inter5), .b(gate310inter2), .O(gate310inter6));
  inv1  gate601(.a(N628), .O(gate310inter7));
  inv1  gate602(.a(N773), .O(gate310inter8));
  nand2 gate603(.a(gate310inter8), .b(gate310inter7), .O(gate310inter9));
  nand2 gate604(.a(s_31), .b(gate310inter3), .O(gate310inter10));
  nor2  gate605(.a(gate310inter10), .b(gate310inter9), .O(gate310inter11));
  nor2  gate606(.a(gate310inter11), .b(gate310inter6), .O(gate310inter12));
  nand2 gate607(.a(gate310inter12), .b(gate310inter1), .O(N795));
nand2 gate311( .a(N795), .b(N747), .O(N796) );
nor2 gate312( .a(N788), .b(N789), .O(N802) );
nor2 gate313( .a(N790), .b(N791), .O(N803) );

  xor2  gate636(.a(N793), .b(N792), .O(gate314inter0));
  nand2 gate637(.a(gate314inter0), .b(s_36), .O(gate314inter1));
  and2  gate638(.a(N793), .b(N792), .O(gate314inter2));
  inv1  gate639(.a(s_36), .O(gate314inter3));
  inv1  gate640(.a(s_37), .O(gate314inter4));
  nand2 gate641(.a(gate314inter4), .b(gate314inter3), .O(gate314inter5));
  nor2  gate642(.a(gate314inter5), .b(gate314inter2), .O(gate314inter6));
  inv1  gate643(.a(N792), .O(gate314inter7));
  inv1  gate644(.a(N793), .O(gate314inter8));
  nand2 gate645(.a(gate314inter8), .b(gate314inter7), .O(gate314inter9));
  nand2 gate646(.a(s_37), .b(gate314inter3), .O(gate314inter10));
  nor2  gate647(.a(gate314inter10), .b(gate314inter9), .O(gate314inter11));
  nor2  gate648(.a(gate314inter11), .b(gate314inter6), .O(gate314inter12));
  nand2 gate649(.a(gate314inter12), .b(gate314inter1), .O(N804));

  xor2  gate440(.a(N794), .b(N340), .O(gate315inter0));
  nand2 gate441(.a(gate315inter0), .b(s_8), .O(gate315inter1));
  and2  gate442(.a(N794), .b(N340), .O(gate315inter2));
  inv1  gate443(.a(s_8), .O(gate315inter3));
  inv1  gate444(.a(s_9), .O(gate315inter4));
  nand2 gate445(.a(gate315inter4), .b(gate315inter3), .O(gate315inter5));
  nor2  gate446(.a(gate315inter5), .b(gate315inter2), .O(gate315inter6));
  inv1  gate447(.a(N340), .O(gate315inter7));
  inv1  gate448(.a(N794), .O(gate315inter8));
  nand2 gate449(.a(gate315inter8), .b(gate315inter7), .O(gate315inter9));
  nand2 gate450(.a(s_9), .b(gate315inter3), .O(gate315inter10));
  nor2  gate451(.a(gate315inter10), .b(gate315inter9), .O(gate315inter11));
  nor2  gate452(.a(gate315inter11), .b(gate315inter6), .O(gate315inter12));
  nand2 gate453(.a(gate315inter12), .b(gate315inter1), .O(N805));
nor2 gate316( .a(N692), .b(N796), .O(N806) );
and2 gate317( .a(N692), .b(N796), .O(N807) );
and2 gate318( .a(N219), .b(N802), .O(N808) );
and2 gate319( .a(N219), .b(N803), .O(N809) );
and2 gate320( .a(N219), .b(N804), .O(N810) );
nand4 gate321( .a(N805), .b(N787), .c(N731), .d(N529), .O(N811) );
nand2 gate322( .a(N619), .b(N796), .O(N812) );
nand3 gate323( .a(N609), .b(N619), .c(N796), .O(N813) );
nand4 gate324( .a(N600), .b(N609), .c(N619), .d(N796), .O(N814) );
nand4 gate325( .a(N738), .b(N765), .c(N766), .d(N814), .O(N815) );
nand3 gate326( .a(N741), .b(N764), .c(N813), .O(N819) );
nand2 gate327( .a(N744), .b(N812), .O(N822) );
nor2 gate328( .a(N806), .b(N807), .O(N825) );
nor2 gate329( .a(N335), .b(N808), .O(N826) );
nor2 gate330( .a(N336), .b(N809), .O(N827) );
nor2 gate331( .a(N338), .b(N810), .O(N828) );
inv1 gate332( .a(N811), .O(N829) );

  xor2  gate678(.a(N815), .b(N665), .O(gate333inter0));
  nand2 gate679(.a(gate333inter0), .b(s_42), .O(gate333inter1));
  and2  gate680(.a(N815), .b(N665), .O(gate333inter2));
  inv1  gate681(.a(s_42), .O(gate333inter3));
  inv1  gate682(.a(s_43), .O(gate333inter4));
  nand2 gate683(.a(gate333inter4), .b(gate333inter3), .O(gate333inter5));
  nor2  gate684(.a(gate333inter5), .b(gate333inter2), .O(gate333inter6));
  inv1  gate685(.a(N665), .O(gate333inter7));
  inv1  gate686(.a(N815), .O(gate333inter8));
  nand2 gate687(.a(gate333inter8), .b(gate333inter7), .O(gate333inter9));
  nand2 gate688(.a(s_43), .b(gate333inter3), .O(gate333inter10));
  nor2  gate689(.a(gate333inter10), .b(gate333inter9), .O(gate333inter11));
  nor2  gate690(.a(gate333inter11), .b(gate333inter6), .O(gate333inter12));
  nand2 gate691(.a(gate333inter12), .b(gate333inter1), .O(N830));
and2 gate334( .a(N665), .b(N815), .O(N831) );
nor2 gate335( .a(N673), .b(N819), .O(N832) );
and2 gate336( .a(N673), .b(N819), .O(N833) );

  xor2  gate566(.a(N822), .b(N682), .O(gate337inter0));
  nand2 gate567(.a(gate337inter0), .b(s_26), .O(gate337inter1));
  and2  gate568(.a(N822), .b(N682), .O(gate337inter2));
  inv1  gate569(.a(s_26), .O(gate337inter3));
  inv1  gate570(.a(s_27), .O(gate337inter4));
  nand2 gate571(.a(gate337inter4), .b(gate337inter3), .O(gate337inter5));
  nor2  gate572(.a(gate337inter5), .b(gate337inter2), .O(gate337inter6));
  inv1  gate573(.a(N682), .O(gate337inter7));
  inv1  gate574(.a(N822), .O(gate337inter8));
  nand2 gate575(.a(gate337inter8), .b(gate337inter7), .O(gate337inter9));
  nand2 gate576(.a(s_27), .b(gate337inter3), .O(gate337inter10));
  nor2  gate577(.a(gate337inter10), .b(gate337inter9), .O(gate337inter11));
  nor2  gate578(.a(gate337inter11), .b(gate337inter6), .O(gate337inter12));
  nand2 gate579(.a(gate337inter12), .b(gate337inter1), .O(N834));
and2 gate338( .a(N682), .b(N822), .O(N835) );
and2 gate339( .a(N219), .b(N825), .O(N836) );
nand3 gate340( .a(N826), .b(N777), .c(N704), .O(N837) );
nand4 gate341( .a(N827), .b(N781), .c(N712), .d(N527), .O(N838) );
nand4 gate342( .a(N828), .b(N785), .c(N721), .d(N528), .O(N839) );
inv1 gate343( .a(N829), .O(N840) );
nand2 gate344( .a(N815), .b(N593), .O(N841) );
nor2 gate345( .a(N830), .b(N831), .O(N842) );
nor2 gate346( .a(N832), .b(N833), .O(N843) );
nor2 gate347( .a(N834), .b(N835), .O(N844) );

  xor2  gate762(.a(N836), .b(N334), .O(gate348inter0));
  nand2 gate763(.a(gate348inter0), .b(s_54), .O(gate348inter1));
  and2  gate764(.a(N836), .b(N334), .O(gate348inter2));
  inv1  gate765(.a(s_54), .O(gate348inter3));
  inv1  gate766(.a(s_55), .O(gate348inter4));
  nand2 gate767(.a(gate348inter4), .b(gate348inter3), .O(gate348inter5));
  nor2  gate768(.a(gate348inter5), .b(gate348inter2), .O(gate348inter6));
  inv1  gate769(.a(N334), .O(gate348inter7));
  inv1  gate770(.a(N836), .O(gate348inter8));
  nand2 gate771(.a(gate348inter8), .b(gate348inter7), .O(gate348inter9));
  nand2 gate772(.a(s_55), .b(gate348inter3), .O(gate348inter10));
  nor2  gate773(.a(gate348inter10), .b(gate348inter9), .O(gate348inter11));
  nor2  gate774(.a(gate348inter11), .b(gate348inter6), .O(gate348inter12));
  nand2 gate775(.a(gate348inter12), .b(gate348inter1), .O(N845));
inv1 gate349( .a(N837), .O(N846) );
inv1 gate350( .a(N838), .O(N847) );
inv1 gate351( .a(N839), .O(N848) );
and2 gate352( .a(N735), .b(N841), .O(N849) );
buf1 gate353( .a(N840), .O(N850) );
and2 gate354( .a(N219), .b(N842), .O(N851) );
and2 gate355( .a(N219), .b(N843), .O(N852) );
and2 gate356( .a(N219), .b(N844), .O(N853) );
nand3 gate357( .a(N845), .b(N772), .c(N696), .O(N854) );
inv1 gate358( .a(N846), .O(N855) );
inv1 gate359( .a(N847), .O(N856) );
inv1 gate360( .a(N848), .O(N857) );
inv1 gate361( .a(N849), .O(N858) );
nor2 gate362( .a(N417), .b(N851), .O(N859) );
nor2 gate363( .a(N332), .b(N852), .O(N860) );
nor2 gate364( .a(N333), .b(N853), .O(N861) );
inv1 gate365( .a(N854), .O(N862) );
buf1 gate366( .a(N855), .O(N863) );
buf1 gate367( .a(N856), .O(N864) );
buf1 gate368( .a(N857), .O(N865) );
buf1 gate369( .a(N858), .O(N866) );
nand3 gate370( .a(N859), .b(N769), .c(N669), .O(N867) );
nand3 gate371( .a(N860), .b(N770), .c(N677), .O(N868) );
nand3 gate372( .a(N861), .b(N771), .c(N686), .O(N869) );
inv1 gate373( .a(N862), .O(N870) );
inv1 gate374( .a(N867), .O(N871) );
inv1 gate375( .a(N868), .O(N872) );
inv1 gate376( .a(N869), .O(N873) );
buf1 gate377( .a(N870), .O(N874) );
inv1 gate378( .a(N871), .O(N875) );
inv1 gate379( .a(N872), .O(N876) );
inv1 gate380( .a(N873), .O(N877) );
buf1 gate381( .a(N875), .O(N878) );
buf1 gate382( .a(N876), .O(N879) );
buf1 gate383( .a(N877), .O(N880) );

endmodule