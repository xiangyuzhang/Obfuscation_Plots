module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate292inter0, gate292inter1, gate292inter2, gate292inter3, gate292inter4, gate292inter5, gate292inter6, gate292inter7, gate292inter8, gate292inter9, gate292inter10, gate292inter11, gate292inter12, gate165inter0, gate165inter1, gate165inter2, gate165inter3, gate165inter4, gate165inter5, gate165inter6, gate165inter7, gate165inter8, gate165inter9, gate165inter10, gate165inter11, gate165inter12, gate407inter0, gate407inter1, gate407inter2, gate407inter3, gate407inter4, gate407inter5, gate407inter6, gate407inter7, gate407inter8, gate407inter9, gate407inter10, gate407inter11, gate407inter12, gate296inter0, gate296inter1, gate296inter2, gate296inter3, gate296inter4, gate296inter5, gate296inter6, gate296inter7, gate296inter8, gate296inter9, gate296inter10, gate296inter11, gate296inter12, gate265inter0, gate265inter1, gate265inter2, gate265inter3, gate265inter4, gate265inter5, gate265inter6, gate265inter7, gate265inter8, gate265inter9, gate265inter10, gate265inter11, gate265inter12, gate197inter0, gate197inter1, gate197inter2, gate197inter3, gate197inter4, gate197inter5, gate197inter6, gate197inter7, gate197inter8, gate197inter9, gate197inter10, gate197inter11, gate197inter12, gate172inter0, gate172inter1, gate172inter2, gate172inter3, gate172inter4, gate172inter5, gate172inter6, gate172inter7, gate172inter8, gate172inter9, gate172inter10, gate172inter11, gate172inter12, gate77inter0, gate77inter1, gate77inter2, gate77inter3, gate77inter4, gate77inter5, gate77inter6, gate77inter7, gate77inter8, gate77inter9, gate77inter10, gate77inter11, gate77inter12, gate390inter0, gate390inter1, gate390inter2, gate390inter3, gate390inter4, gate390inter5, gate390inter6, gate390inter7, gate390inter8, gate390inter9, gate390inter10, gate390inter11, gate390inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate65inter0, gate65inter1, gate65inter2, gate65inter3, gate65inter4, gate65inter5, gate65inter6, gate65inter7, gate65inter8, gate65inter9, gate65inter10, gate65inter11, gate65inter12, gate446inter0, gate446inter1, gate446inter2, gate446inter3, gate446inter4, gate446inter5, gate446inter6, gate446inter7, gate446inter8, gate446inter9, gate446inter10, gate446inter11, gate446inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate84inter0, gate84inter1, gate84inter2, gate84inter3, gate84inter4, gate84inter5, gate84inter6, gate84inter7, gate84inter8, gate84inter9, gate84inter10, gate84inter11, gate84inter12, gate57inter0, gate57inter1, gate57inter2, gate57inter3, gate57inter4, gate57inter5, gate57inter6, gate57inter7, gate57inter8, gate57inter9, gate57inter10, gate57inter11, gate57inter12, gate463inter0, gate463inter1, gate463inter2, gate463inter3, gate463inter4, gate463inter5, gate463inter6, gate463inter7, gate463inter8, gate463inter9, gate463inter10, gate463inter11, gate463inter12, gate492inter0, gate492inter1, gate492inter2, gate492inter3, gate492inter4, gate492inter5, gate492inter6, gate492inter7, gate492inter8, gate492inter9, gate492inter10, gate492inter11, gate492inter12, gate46inter0, gate46inter1, gate46inter2, gate46inter3, gate46inter4, gate46inter5, gate46inter6, gate46inter7, gate46inter8, gate46inter9, gate46inter10, gate46inter11, gate46inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate496inter0, gate496inter1, gate496inter2, gate496inter3, gate496inter4, gate496inter5, gate496inter6, gate496inter7, gate496inter8, gate496inter9, gate496inter10, gate496inter11, gate496inter12, gate24inter0, gate24inter1, gate24inter2, gate24inter3, gate24inter4, gate24inter5, gate24inter6, gate24inter7, gate24inter8, gate24inter9, gate24inter10, gate24inter11, gate24inter12, gate66inter0, gate66inter1, gate66inter2, gate66inter3, gate66inter4, gate66inter5, gate66inter6, gate66inter7, gate66inter8, gate66inter9, gate66inter10, gate66inter11, gate66inter12, gate99inter0, gate99inter1, gate99inter2, gate99inter3, gate99inter4, gate99inter5, gate99inter6, gate99inter7, gate99inter8, gate99inter9, gate99inter10, gate99inter11, gate99inter12, gate40inter0, gate40inter1, gate40inter2, gate40inter3, gate40inter4, gate40inter5, gate40inter6, gate40inter7, gate40inter8, gate40inter9, gate40inter10, gate40inter11, gate40inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate486inter0, gate486inter1, gate486inter2, gate486inter3, gate486inter4, gate486inter5, gate486inter6, gate486inter7, gate486inter8, gate486inter9, gate486inter10, gate486inter11, gate486inter12, gate277inter0, gate277inter1, gate277inter2, gate277inter3, gate277inter4, gate277inter5, gate277inter6, gate277inter7, gate277inter8, gate277inter9, gate277inter10, gate277inter11, gate277inter12, gate81inter0, gate81inter1, gate81inter2, gate81inter3, gate81inter4, gate81inter5, gate81inter6, gate81inter7, gate81inter8, gate81inter9, gate81inter10, gate81inter11, gate81inter12, gate485inter0, gate485inter1, gate485inter2, gate485inter3, gate485inter4, gate485inter5, gate485inter6, gate485inter7, gate485inter8, gate485inter9, gate485inter10, gate485inter11, gate485inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate103inter0, gate103inter1, gate103inter2, gate103inter3, gate103inter4, gate103inter5, gate103inter6, gate103inter7, gate103inter8, gate103inter9, gate103inter10, gate103inter11, gate103inter12, gate439inter0, gate439inter1, gate439inter2, gate439inter3, gate439inter4, gate439inter5, gate439inter6, gate439inter7, gate439inter8, gate439inter9, gate439inter10, gate439inter11, gate439inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate435inter0, gate435inter1, gate435inter2, gate435inter3, gate435inter4, gate435inter5, gate435inter6, gate435inter7, gate435inter8, gate435inter9, gate435inter10, gate435inter11, gate435inter12, gate37inter0, gate37inter1, gate37inter2, gate37inter3, gate37inter4, gate37inter5, gate37inter6, gate37inter7, gate37inter8, gate37inter9, gate37inter10, gate37inter11, gate37inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate135inter0, gate135inter1, gate135inter2, gate135inter3, gate135inter4, gate135inter5, gate135inter6, gate135inter7, gate135inter8, gate135inter9, gate135inter10, gate135inter11, gate135inter12, gate504inter0, gate504inter1, gate504inter2, gate504inter3, gate504inter4, gate504inter5, gate504inter6, gate504inter7, gate504inter8, gate504inter9, gate504inter10, gate504inter11, gate504inter12, gate145inter0, gate145inter1, gate145inter2, gate145inter3, gate145inter4, gate145inter5, gate145inter6, gate145inter7, gate145inter8, gate145inter9, gate145inter10, gate145inter11, gate145inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate263inter0, gate263inter1, gate263inter2, gate263inter3, gate263inter4, gate263inter5, gate263inter6, gate263inter7, gate263inter8, gate263inter9, gate263inter10, gate263inter11, gate263inter12, gate203inter0, gate203inter1, gate203inter2, gate203inter3, gate203inter4, gate203inter5, gate203inter6, gate203inter7, gate203inter8, gate203inter9, gate203inter10, gate203inter11, gate203inter12, gate258inter0, gate258inter1, gate258inter2, gate258inter3, gate258inter4, gate258inter5, gate258inter6, gate258inter7, gate258inter8, gate258inter9, gate258inter10, gate258inter11, gate258inter12, gate20inter0, gate20inter1, gate20inter2, gate20inter3, gate20inter4, gate20inter5, gate20inter6, gate20inter7, gate20inter8, gate20inter9, gate20inter10, gate20inter11, gate20inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate221inter0, gate221inter1, gate221inter2, gate221inter3, gate221inter4, gate221inter5, gate221inter6, gate221inter7, gate221inter8, gate221inter9, gate221inter10, gate221inter11, gate221inter12, gate464inter0, gate464inter1, gate464inter2, gate464inter3, gate464inter4, gate464inter5, gate464inter6, gate464inter7, gate464inter8, gate464inter9, gate464inter10, gate464inter11, gate464inter12, gate184inter0, gate184inter1, gate184inter2, gate184inter3, gate184inter4, gate184inter5, gate184inter6, gate184inter7, gate184inter8, gate184inter9, gate184inter10, gate184inter11, gate184inter12, gate290inter0, gate290inter1, gate290inter2, gate290inter3, gate290inter4, gate290inter5, gate290inter6, gate290inter7, gate290inter8, gate290inter9, gate290inter10, gate290inter11, gate290inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate441inter0, gate441inter1, gate441inter2, gate441inter3, gate441inter4, gate441inter5, gate441inter6, gate441inter7, gate441inter8, gate441inter9, gate441inter10, gate441inter11, gate441inter12, gate285inter0, gate285inter1, gate285inter2, gate285inter3, gate285inter4, gate285inter5, gate285inter6, gate285inter7, gate285inter8, gate285inter9, gate285inter10, gate285inter11, gate285inter12, gate168inter0, gate168inter1, gate168inter2, gate168inter3, gate168inter4, gate168inter5, gate168inter6, gate168inter7, gate168inter8, gate168inter9, gate168inter10, gate168inter11, gate168inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate89inter0, gate89inter1, gate89inter2, gate89inter3, gate89inter4, gate89inter5, gate89inter6, gate89inter7, gate89inter8, gate89inter9, gate89inter10, gate89inter11, gate89inter12, gate160inter0, gate160inter1, gate160inter2, gate160inter3, gate160inter4, gate160inter5, gate160inter6, gate160inter7, gate160inter8, gate160inter9, gate160inter10, gate160inter11, gate160inter12, gate391inter0, gate391inter1, gate391inter2, gate391inter3, gate391inter4, gate391inter5, gate391inter6, gate391inter7, gate391inter8, gate391inter9, gate391inter10, gate391inter11, gate391inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate511inter0, gate511inter1, gate511inter2, gate511inter3, gate511inter4, gate511inter5, gate511inter6, gate511inter7, gate511inter8, gate511inter9, gate511inter10, gate511inter11, gate511inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate62inter0, gate62inter1, gate62inter2, gate62inter3, gate62inter4, gate62inter5, gate62inter6, gate62inter7, gate62inter8, gate62inter9, gate62inter10, gate62inter11, gate62inter12, gate251inter0, gate251inter1, gate251inter2, gate251inter3, gate251inter4, gate251inter5, gate251inter6, gate251inter7, gate251inter8, gate251inter9, gate251inter10, gate251inter11, gate251inter12, gate293inter0, gate293inter1, gate293inter2, gate293inter3, gate293inter4, gate293inter5, gate293inter6, gate293inter7, gate293inter8, gate293inter9, gate293inter10, gate293inter11, gate293inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate422inter0, gate422inter1, gate422inter2, gate422inter3, gate422inter4, gate422inter5, gate422inter6, gate422inter7, gate422inter8, gate422inter9, gate422inter10, gate422inter11, gate422inter12, gate125inter0, gate125inter1, gate125inter2, gate125inter3, gate125inter4, gate125inter5, gate125inter6, gate125inter7, gate125inter8, gate125inter9, gate125inter10, gate125inter11, gate125inter12, gate403inter0, gate403inter1, gate403inter2, gate403inter3, gate403inter4, gate403inter5, gate403inter6, gate403inter7, gate403inter8, gate403inter9, gate403inter10, gate403inter11, gate403inter12, gate61inter0, gate61inter1, gate61inter2, gate61inter3, gate61inter4, gate61inter5, gate61inter6, gate61inter7, gate61inter8, gate61inter9, gate61inter10, gate61inter11, gate61inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate262inter0, gate262inter1, gate262inter2, gate262inter3, gate262inter4, gate262inter5, gate262inter6, gate262inter7, gate262inter8, gate262inter9, gate262inter10, gate262inter11, gate262inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate162inter0, gate162inter1, gate162inter2, gate162inter3, gate162inter4, gate162inter5, gate162inter6, gate162inter7, gate162inter8, gate162inter9, gate162inter10, gate162inter11, gate162inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate38inter0, gate38inter1, gate38inter2, gate38inter3, gate38inter4, gate38inter5, gate38inter6, gate38inter7, gate38inter8, gate38inter9, gate38inter10, gate38inter11, gate38inter12, gate148inter0, gate148inter1, gate148inter2, gate148inter3, gate148inter4, gate148inter5, gate148inter6, gate148inter7, gate148inter8, gate148inter9, gate148inter10, gate148inter11, gate148inter12, gate400inter0, gate400inter1, gate400inter2, gate400inter3, gate400inter4, gate400inter5, gate400inter6, gate400inter7, gate400inter8, gate400inter9, gate400inter10, gate400inter11, gate400inter12, gate219inter0, gate219inter1, gate219inter2, gate219inter3, gate219inter4, gate219inter5, gate219inter6, gate219inter7, gate219inter8, gate219inter9, gate219inter10, gate219inter11, gate219inter12, gate443inter0, gate443inter1, gate443inter2, gate443inter3, gate443inter4, gate443inter5, gate443inter6, gate443inter7, gate443inter8, gate443inter9, gate443inter10, gate443inter11, gate443inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate453inter0, gate453inter1, gate453inter2, gate453inter3, gate453inter4, gate453inter5, gate453inter6, gate453inter7, gate453inter8, gate453inter9, gate453inter10, gate453inter11, gate453inter12, gate188inter0, gate188inter1, gate188inter2, gate188inter3, gate188inter4, gate188inter5, gate188inter6, gate188inter7, gate188inter8, gate188inter9, gate188inter10, gate188inter11, gate188inter12, gate15inter0, gate15inter1, gate15inter2, gate15inter3, gate15inter4, gate15inter5, gate15inter6, gate15inter7, gate15inter8, gate15inter9, gate15inter10, gate15inter11, gate15inter12, gate218inter0, gate218inter1, gate218inter2, gate218inter3, gate218inter4, gate218inter5, gate218inter6, gate218inter7, gate218inter8, gate218inter9, gate218inter10, gate218inter11, gate218inter12, gate510inter0, gate510inter1, gate510inter2, gate510inter3, gate510inter4, gate510inter5, gate510inter6, gate510inter7, gate510inter8, gate510inter9, gate510inter10, gate510inter11, gate510inter12, gate174inter0, gate174inter1, gate174inter2, gate174inter3, gate174inter4, gate174inter5, gate174inter6, gate174inter7, gate174inter8, gate174inter9, gate174inter10, gate174inter11, gate174inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate478inter0, gate478inter1, gate478inter2, gate478inter3, gate478inter4, gate478inter5, gate478inter6, gate478inter7, gate478inter8, gate478inter9, gate478inter10, gate478inter11, gate478inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );
nand2 gate9( .a(G1), .b(G2), .O(G266) );
nand2 gate10( .a(G3), .b(G4), .O(G269) );
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );
nand2 gate13( .a(G9), .b(G10), .O(G278) );
nand2 gate14( .a(G11), .b(G12), .O(G281) );

  xor2  gate1737(.a(G14), .b(G13), .O(gate15inter0));
  nand2 gate1738(.a(gate15inter0), .b(s_170), .O(gate15inter1));
  and2  gate1739(.a(G14), .b(G13), .O(gate15inter2));
  inv1  gate1740(.a(s_170), .O(gate15inter3));
  inv1  gate1741(.a(s_171), .O(gate15inter4));
  nand2 gate1742(.a(gate15inter4), .b(gate15inter3), .O(gate15inter5));
  nor2  gate1743(.a(gate15inter5), .b(gate15inter2), .O(gate15inter6));
  inv1  gate1744(.a(G13), .O(gate15inter7));
  inv1  gate1745(.a(G14), .O(gate15inter8));
  nand2 gate1746(.a(gate15inter8), .b(gate15inter7), .O(gate15inter9));
  nand2 gate1747(.a(s_171), .b(gate15inter3), .O(gate15inter10));
  nor2  gate1748(.a(gate15inter10), .b(gate15inter9), .O(gate15inter11));
  nor2  gate1749(.a(gate15inter11), .b(gate15inter6), .O(gate15inter12));
  nand2 gate1750(.a(gate15inter12), .b(gate15inter1), .O(G284));
nand2 gate16( .a(G15), .b(G16), .O(G287) );
nand2 gate17( .a(G17), .b(G18), .O(G290) );
nand2 gate18( .a(G19), .b(G20), .O(G293) );
nand2 gate19( .a(G21), .b(G22), .O(G296) );

  xor2  gate1191(.a(G24), .b(G23), .O(gate20inter0));
  nand2 gate1192(.a(gate20inter0), .b(s_92), .O(gate20inter1));
  and2  gate1193(.a(G24), .b(G23), .O(gate20inter2));
  inv1  gate1194(.a(s_92), .O(gate20inter3));
  inv1  gate1195(.a(s_93), .O(gate20inter4));
  nand2 gate1196(.a(gate20inter4), .b(gate20inter3), .O(gate20inter5));
  nor2  gate1197(.a(gate20inter5), .b(gate20inter2), .O(gate20inter6));
  inv1  gate1198(.a(G23), .O(gate20inter7));
  inv1  gate1199(.a(G24), .O(gate20inter8));
  nand2 gate1200(.a(gate20inter8), .b(gate20inter7), .O(gate20inter9));
  nand2 gate1201(.a(s_93), .b(gate20inter3), .O(gate20inter10));
  nor2  gate1202(.a(gate20inter10), .b(gate20inter9), .O(gate20inter11));
  nor2  gate1203(.a(gate20inter11), .b(gate20inter6), .O(gate20inter12));
  nand2 gate1204(.a(gate20inter12), .b(gate20inter1), .O(G299));
nand2 gate21( .a(G25), .b(G26), .O(G302) );
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );

  xor2  gate869(.a(G32), .b(G31), .O(gate24inter0));
  nand2 gate870(.a(gate24inter0), .b(s_46), .O(gate24inter1));
  and2  gate871(.a(G32), .b(G31), .O(gate24inter2));
  inv1  gate872(.a(s_46), .O(gate24inter3));
  inv1  gate873(.a(s_47), .O(gate24inter4));
  nand2 gate874(.a(gate24inter4), .b(gate24inter3), .O(gate24inter5));
  nor2  gate875(.a(gate24inter5), .b(gate24inter2), .O(gate24inter6));
  inv1  gate876(.a(G31), .O(gate24inter7));
  inv1  gate877(.a(G32), .O(gate24inter8));
  nand2 gate878(.a(gate24inter8), .b(gate24inter7), .O(gate24inter9));
  nand2 gate879(.a(s_47), .b(gate24inter3), .O(gate24inter10));
  nor2  gate880(.a(gate24inter10), .b(gate24inter9), .O(gate24inter11));
  nor2  gate881(.a(gate24inter11), .b(gate24inter6), .O(gate24inter12));
  nand2 gate882(.a(gate24inter12), .b(gate24inter1), .O(G311));
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );
nand2 gate27( .a(G2), .b(G6), .O(G320) );
nand2 gate28( .a(G10), .b(G14), .O(G323) );
nand2 gate29( .a(G3), .b(G7), .O(G326) );
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate1205(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate1206(.a(gate31inter0), .b(s_94), .O(gate31inter1));
  and2  gate1207(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate1208(.a(s_94), .O(gate31inter3));
  inv1  gate1209(.a(s_95), .O(gate31inter4));
  nand2 gate1210(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate1211(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate1212(.a(G4), .O(gate31inter7));
  inv1  gate1213(.a(G8), .O(gate31inter8));
  nand2 gate1214(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate1215(.a(s_95), .b(gate31inter3), .O(gate31inter10));
  nor2  gate1216(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate1217(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate1218(.a(gate31inter12), .b(gate31inter1), .O(G332));

  xor2  gate1583(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate1584(.a(gate32inter0), .b(s_148), .O(gate32inter1));
  and2  gate1585(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate1586(.a(s_148), .O(gate32inter3));
  inv1  gate1587(.a(s_149), .O(gate32inter4));
  nand2 gate1588(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate1589(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate1590(.a(G12), .O(gate32inter7));
  inv1  gate1591(.a(G16), .O(gate32inter8));
  nand2 gate1592(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate1593(.a(s_149), .b(gate32inter3), .O(gate32inter10));
  nor2  gate1594(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate1595(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate1596(.a(gate32inter12), .b(gate32inter1), .O(G335));
nand2 gate33( .a(G17), .b(G21), .O(G338) );
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );

  xor2  gate1065(.a(G23), .b(G19), .O(gate37inter0));
  nand2 gate1066(.a(gate37inter0), .b(s_74), .O(gate37inter1));
  and2  gate1067(.a(G23), .b(G19), .O(gate37inter2));
  inv1  gate1068(.a(s_74), .O(gate37inter3));
  inv1  gate1069(.a(s_75), .O(gate37inter4));
  nand2 gate1070(.a(gate37inter4), .b(gate37inter3), .O(gate37inter5));
  nor2  gate1071(.a(gate37inter5), .b(gate37inter2), .O(gate37inter6));
  inv1  gate1072(.a(G19), .O(gate37inter7));
  inv1  gate1073(.a(G23), .O(gate37inter8));
  nand2 gate1074(.a(gate37inter8), .b(gate37inter7), .O(gate37inter9));
  nand2 gate1075(.a(s_75), .b(gate37inter3), .O(gate37inter10));
  nor2  gate1076(.a(gate37inter10), .b(gate37inter9), .O(gate37inter11));
  nor2  gate1077(.a(gate37inter11), .b(gate37inter6), .O(gate37inter12));
  nand2 gate1078(.a(gate37inter12), .b(gate37inter1), .O(G350));

  xor2  gate1625(.a(G31), .b(G27), .O(gate38inter0));
  nand2 gate1626(.a(gate38inter0), .b(s_154), .O(gate38inter1));
  and2  gate1627(.a(G31), .b(G27), .O(gate38inter2));
  inv1  gate1628(.a(s_154), .O(gate38inter3));
  inv1  gate1629(.a(s_155), .O(gate38inter4));
  nand2 gate1630(.a(gate38inter4), .b(gate38inter3), .O(gate38inter5));
  nor2  gate1631(.a(gate38inter5), .b(gate38inter2), .O(gate38inter6));
  inv1  gate1632(.a(G27), .O(gate38inter7));
  inv1  gate1633(.a(G31), .O(gate38inter8));
  nand2 gate1634(.a(gate38inter8), .b(gate38inter7), .O(gate38inter9));
  nand2 gate1635(.a(s_155), .b(gate38inter3), .O(gate38inter10));
  nor2  gate1636(.a(gate38inter10), .b(gate38inter9), .O(gate38inter11));
  nor2  gate1637(.a(gate38inter11), .b(gate38inter6), .O(gate38inter12));
  nand2 gate1638(.a(gate38inter12), .b(gate38inter1), .O(G353));
nand2 gate39( .a(G20), .b(G24), .O(G356) );

  xor2  gate911(.a(G32), .b(G28), .O(gate40inter0));
  nand2 gate912(.a(gate40inter0), .b(s_52), .O(gate40inter1));
  and2  gate913(.a(G32), .b(G28), .O(gate40inter2));
  inv1  gate914(.a(s_52), .O(gate40inter3));
  inv1  gate915(.a(s_53), .O(gate40inter4));
  nand2 gate916(.a(gate40inter4), .b(gate40inter3), .O(gate40inter5));
  nor2  gate917(.a(gate40inter5), .b(gate40inter2), .O(gate40inter6));
  inv1  gate918(.a(G28), .O(gate40inter7));
  inv1  gate919(.a(G32), .O(gate40inter8));
  nand2 gate920(.a(gate40inter8), .b(gate40inter7), .O(gate40inter9));
  nand2 gate921(.a(s_53), .b(gate40inter3), .O(gate40inter10));
  nor2  gate922(.a(gate40inter10), .b(gate40inter9), .O(gate40inter11));
  nor2  gate923(.a(gate40inter11), .b(gate40inter6), .O(gate40inter12));
  nand2 gate924(.a(gate40inter12), .b(gate40inter1), .O(G359));
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );
nand2 gate43( .a(G3), .b(G269), .O(G364) );
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );

  xor2  gate813(.a(G272), .b(G6), .O(gate46inter0));
  nand2 gate814(.a(gate46inter0), .b(s_38), .O(gate46inter1));
  and2  gate815(.a(G272), .b(G6), .O(gate46inter2));
  inv1  gate816(.a(s_38), .O(gate46inter3));
  inv1  gate817(.a(s_39), .O(gate46inter4));
  nand2 gate818(.a(gate46inter4), .b(gate46inter3), .O(gate46inter5));
  nor2  gate819(.a(gate46inter5), .b(gate46inter2), .O(gate46inter6));
  inv1  gate820(.a(G6), .O(gate46inter7));
  inv1  gate821(.a(G272), .O(gate46inter8));
  nand2 gate822(.a(gate46inter8), .b(gate46inter7), .O(gate46inter9));
  nand2 gate823(.a(s_39), .b(gate46inter3), .O(gate46inter10));
  nor2  gate824(.a(gate46inter10), .b(gate46inter9), .O(gate46inter11));
  nor2  gate825(.a(gate46inter11), .b(gate46inter6), .O(gate46inter12));
  nand2 gate826(.a(gate46inter12), .b(gate46inter1), .O(G367));
nand2 gate47( .a(G7), .b(G275), .O(G368) );
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );

  xor2  gate1331(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate1332(.a(gate53inter0), .b(s_112), .O(gate53inter1));
  and2  gate1333(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate1334(.a(s_112), .O(gate53inter3));
  inv1  gate1335(.a(s_113), .O(gate53inter4));
  nand2 gate1336(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate1337(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate1338(.a(G13), .O(gate53inter7));
  inv1  gate1339(.a(G284), .O(gate53inter8));
  nand2 gate1340(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate1341(.a(s_113), .b(gate53inter3), .O(gate53inter10));
  nor2  gate1342(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate1343(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate1344(.a(gate53inter12), .b(gate53inter1), .O(G374));
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );

  xor2  gate771(.a(G290), .b(G17), .O(gate57inter0));
  nand2 gate772(.a(gate57inter0), .b(s_32), .O(gate57inter1));
  and2  gate773(.a(G290), .b(G17), .O(gate57inter2));
  inv1  gate774(.a(s_32), .O(gate57inter3));
  inv1  gate775(.a(s_33), .O(gate57inter4));
  nand2 gate776(.a(gate57inter4), .b(gate57inter3), .O(gate57inter5));
  nor2  gate777(.a(gate57inter5), .b(gate57inter2), .O(gate57inter6));
  inv1  gate778(.a(G17), .O(gate57inter7));
  inv1  gate779(.a(G290), .O(gate57inter8));
  nand2 gate780(.a(gate57inter8), .b(gate57inter7), .O(gate57inter9));
  nand2 gate781(.a(s_33), .b(gate57inter3), .O(gate57inter10));
  nor2  gate782(.a(gate57inter10), .b(gate57inter9), .O(gate57inter11));
  nor2  gate783(.a(gate57inter11), .b(gate57inter6), .O(gate57inter12));
  nand2 gate784(.a(gate57inter12), .b(gate57inter1), .O(G378));
nand2 gate58( .a(G18), .b(G290), .O(G379) );
nand2 gate59( .a(G19), .b(G293), .O(G380) );
nand2 gate60( .a(G20), .b(G293), .O(G381) );

  xor2  gate1527(.a(G296), .b(G21), .O(gate61inter0));
  nand2 gate1528(.a(gate61inter0), .b(s_140), .O(gate61inter1));
  and2  gate1529(.a(G296), .b(G21), .O(gate61inter2));
  inv1  gate1530(.a(s_140), .O(gate61inter3));
  inv1  gate1531(.a(s_141), .O(gate61inter4));
  nand2 gate1532(.a(gate61inter4), .b(gate61inter3), .O(gate61inter5));
  nor2  gate1533(.a(gate61inter5), .b(gate61inter2), .O(gate61inter6));
  inv1  gate1534(.a(G21), .O(gate61inter7));
  inv1  gate1535(.a(G296), .O(gate61inter8));
  nand2 gate1536(.a(gate61inter8), .b(gate61inter7), .O(gate61inter9));
  nand2 gate1537(.a(s_141), .b(gate61inter3), .O(gate61inter10));
  nor2  gate1538(.a(gate61inter10), .b(gate61inter9), .O(gate61inter11));
  nor2  gate1539(.a(gate61inter11), .b(gate61inter6), .O(gate61inter12));
  nand2 gate1540(.a(gate61inter12), .b(gate61inter1), .O(G382));

  xor2  gate1429(.a(G296), .b(G22), .O(gate62inter0));
  nand2 gate1430(.a(gate62inter0), .b(s_126), .O(gate62inter1));
  and2  gate1431(.a(G296), .b(G22), .O(gate62inter2));
  inv1  gate1432(.a(s_126), .O(gate62inter3));
  inv1  gate1433(.a(s_127), .O(gate62inter4));
  nand2 gate1434(.a(gate62inter4), .b(gate62inter3), .O(gate62inter5));
  nor2  gate1435(.a(gate62inter5), .b(gate62inter2), .O(gate62inter6));
  inv1  gate1436(.a(G22), .O(gate62inter7));
  inv1  gate1437(.a(G296), .O(gate62inter8));
  nand2 gate1438(.a(gate62inter8), .b(gate62inter7), .O(gate62inter9));
  nand2 gate1439(.a(s_127), .b(gate62inter3), .O(gate62inter10));
  nor2  gate1440(.a(gate62inter10), .b(gate62inter9), .O(gate62inter11));
  nor2  gate1441(.a(gate62inter11), .b(gate62inter6), .O(gate62inter12));
  nand2 gate1442(.a(gate62inter12), .b(gate62inter1), .O(G383));
nand2 gate63( .a(G23), .b(G299), .O(G384) );
nand2 gate64( .a(G24), .b(G299), .O(G385) );

  xor2  gate701(.a(G302), .b(G25), .O(gate65inter0));
  nand2 gate702(.a(gate65inter0), .b(s_22), .O(gate65inter1));
  and2  gate703(.a(G302), .b(G25), .O(gate65inter2));
  inv1  gate704(.a(s_22), .O(gate65inter3));
  inv1  gate705(.a(s_23), .O(gate65inter4));
  nand2 gate706(.a(gate65inter4), .b(gate65inter3), .O(gate65inter5));
  nor2  gate707(.a(gate65inter5), .b(gate65inter2), .O(gate65inter6));
  inv1  gate708(.a(G25), .O(gate65inter7));
  inv1  gate709(.a(G302), .O(gate65inter8));
  nand2 gate710(.a(gate65inter8), .b(gate65inter7), .O(gate65inter9));
  nand2 gate711(.a(s_23), .b(gate65inter3), .O(gate65inter10));
  nor2  gate712(.a(gate65inter10), .b(gate65inter9), .O(gate65inter11));
  nor2  gate713(.a(gate65inter11), .b(gate65inter6), .O(gate65inter12));
  nand2 gate714(.a(gate65inter12), .b(gate65inter1), .O(G386));

  xor2  gate883(.a(G302), .b(G26), .O(gate66inter0));
  nand2 gate884(.a(gate66inter0), .b(s_48), .O(gate66inter1));
  and2  gate885(.a(G302), .b(G26), .O(gate66inter2));
  inv1  gate886(.a(s_48), .O(gate66inter3));
  inv1  gate887(.a(s_49), .O(gate66inter4));
  nand2 gate888(.a(gate66inter4), .b(gate66inter3), .O(gate66inter5));
  nor2  gate889(.a(gate66inter5), .b(gate66inter2), .O(gate66inter6));
  inv1  gate890(.a(G26), .O(gate66inter7));
  inv1  gate891(.a(G302), .O(gate66inter8));
  nand2 gate892(.a(gate66inter8), .b(gate66inter7), .O(gate66inter9));
  nand2 gate893(.a(s_49), .b(gate66inter3), .O(gate66inter10));
  nor2  gate894(.a(gate66inter10), .b(gate66inter9), .O(gate66inter11));
  nor2  gate895(.a(gate66inter11), .b(gate66inter6), .O(gate66inter12));
  nand2 gate896(.a(gate66inter12), .b(gate66inter1), .O(G387));
nand2 gate67( .a(G27), .b(G305), .O(G388) );
nand2 gate68( .a(G28), .b(G305), .O(G389) );
nand2 gate69( .a(G29), .b(G308), .O(G390) );
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate673(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate674(.a(gate71inter0), .b(s_18), .O(gate71inter1));
  and2  gate675(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate676(.a(s_18), .O(gate71inter3));
  inv1  gate677(.a(s_19), .O(gate71inter4));
  nand2 gate678(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate679(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate680(.a(G31), .O(gate71inter7));
  inv1  gate681(.a(G311), .O(gate71inter8));
  nand2 gate682(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate683(.a(s_19), .b(gate71inter3), .O(gate71inter10));
  nor2  gate684(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate685(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate686(.a(gate71inter12), .b(gate71inter1), .O(G392));
nand2 gate72( .a(G32), .b(G311), .O(G393) );
nand2 gate73( .a(G1), .b(G314), .O(G394) );
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );
nand2 gate76( .a(G13), .b(G317), .O(G397) );

  xor2  gate645(.a(G320), .b(G2), .O(gate77inter0));
  nand2 gate646(.a(gate77inter0), .b(s_14), .O(gate77inter1));
  and2  gate647(.a(G320), .b(G2), .O(gate77inter2));
  inv1  gate648(.a(s_14), .O(gate77inter3));
  inv1  gate649(.a(s_15), .O(gate77inter4));
  nand2 gate650(.a(gate77inter4), .b(gate77inter3), .O(gate77inter5));
  nor2  gate651(.a(gate77inter5), .b(gate77inter2), .O(gate77inter6));
  inv1  gate652(.a(G2), .O(gate77inter7));
  inv1  gate653(.a(G320), .O(gate77inter8));
  nand2 gate654(.a(gate77inter8), .b(gate77inter7), .O(gate77inter9));
  nand2 gate655(.a(s_15), .b(gate77inter3), .O(gate77inter10));
  nor2  gate656(.a(gate77inter10), .b(gate77inter9), .O(gate77inter11));
  nor2  gate657(.a(gate77inter11), .b(gate77inter6), .O(gate77inter12));
  nand2 gate658(.a(gate77inter12), .b(gate77inter1), .O(G398));
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );

  xor2  gate967(.a(G326), .b(G3), .O(gate81inter0));
  nand2 gate968(.a(gate81inter0), .b(s_60), .O(gate81inter1));
  and2  gate969(.a(G326), .b(G3), .O(gate81inter2));
  inv1  gate970(.a(s_60), .O(gate81inter3));
  inv1  gate971(.a(s_61), .O(gate81inter4));
  nand2 gate972(.a(gate81inter4), .b(gate81inter3), .O(gate81inter5));
  nor2  gate973(.a(gate81inter5), .b(gate81inter2), .O(gate81inter6));
  inv1  gate974(.a(G3), .O(gate81inter7));
  inv1  gate975(.a(G326), .O(gate81inter8));
  nand2 gate976(.a(gate81inter8), .b(gate81inter7), .O(gate81inter9));
  nand2 gate977(.a(s_61), .b(gate81inter3), .O(gate81inter10));
  nor2  gate978(.a(gate81inter10), .b(gate81inter9), .O(gate81inter11));
  nor2  gate979(.a(gate81inter11), .b(gate81inter6), .O(gate81inter12));
  nand2 gate980(.a(gate81inter12), .b(gate81inter1), .O(G402));
nand2 gate82( .a(G7), .b(G326), .O(G403) );
nand2 gate83( .a(G11), .b(G329), .O(G404) );

  xor2  gate757(.a(G329), .b(G15), .O(gate84inter0));
  nand2 gate758(.a(gate84inter0), .b(s_30), .O(gate84inter1));
  and2  gate759(.a(G329), .b(G15), .O(gate84inter2));
  inv1  gate760(.a(s_30), .O(gate84inter3));
  inv1  gate761(.a(s_31), .O(gate84inter4));
  nand2 gate762(.a(gate84inter4), .b(gate84inter3), .O(gate84inter5));
  nor2  gate763(.a(gate84inter5), .b(gate84inter2), .O(gate84inter6));
  inv1  gate764(.a(G15), .O(gate84inter7));
  inv1  gate765(.a(G329), .O(gate84inter8));
  nand2 gate766(.a(gate84inter8), .b(gate84inter7), .O(gate84inter9));
  nand2 gate767(.a(s_31), .b(gate84inter3), .O(gate84inter10));
  nor2  gate768(.a(gate84inter10), .b(gate84inter9), .O(gate84inter11));
  nor2  gate769(.a(gate84inter11), .b(gate84inter6), .O(gate84inter12));
  nand2 gate770(.a(gate84inter12), .b(gate84inter1), .O(G405));
nand2 gate85( .a(G4), .b(G332), .O(G406) );
nand2 gate86( .a(G8), .b(G332), .O(G407) );
nand2 gate87( .a(G12), .b(G335), .O(G408) );
nand2 gate88( .a(G16), .b(G335), .O(G409) );

  xor2  gate1345(.a(G338), .b(G17), .O(gate89inter0));
  nand2 gate1346(.a(gate89inter0), .b(s_114), .O(gate89inter1));
  and2  gate1347(.a(G338), .b(G17), .O(gate89inter2));
  inv1  gate1348(.a(s_114), .O(gate89inter3));
  inv1  gate1349(.a(s_115), .O(gate89inter4));
  nand2 gate1350(.a(gate89inter4), .b(gate89inter3), .O(gate89inter5));
  nor2  gate1351(.a(gate89inter5), .b(gate89inter2), .O(gate89inter6));
  inv1  gate1352(.a(G17), .O(gate89inter7));
  inv1  gate1353(.a(G338), .O(gate89inter8));
  nand2 gate1354(.a(gate89inter8), .b(gate89inter7), .O(gate89inter9));
  nand2 gate1355(.a(s_115), .b(gate89inter3), .O(gate89inter10));
  nor2  gate1356(.a(gate89inter10), .b(gate89inter9), .O(gate89inter11));
  nor2  gate1357(.a(gate89inter11), .b(gate89inter6), .O(gate89inter12));
  nand2 gate1358(.a(gate89inter12), .b(gate89inter1), .O(G410));
nand2 gate90( .a(G21), .b(G338), .O(G411) );
nand2 gate91( .a(G25), .b(G341), .O(G412) );
nand2 gate92( .a(G29), .b(G341), .O(G413) );
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );

  xor2  gate897(.a(G353), .b(G27), .O(gate99inter0));
  nand2 gate898(.a(gate99inter0), .b(s_50), .O(gate99inter1));
  and2  gate899(.a(G353), .b(G27), .O(gate99inter2));
  inv1  gate900(.a(s_50), .O(gate99inter3));
  inv1  gate901(.a(s_51), .O(gate99inter4));
  nand2 gate902(.a(gate99inter4), .b(gate99inter3), .O(gate99inter5));
  nor2  gate903(.a(gate99inter5), .b(gate99inter2), .O(gate99inter6));
  inv1  gate904(.a(G27), .O(gate99inter7));
  inv1  gate905(.a(G353), .O(gate99inter8));
  nand2 gate906(.a(gate99inter8), .b(gate99inter7), .O(gate99inter9));
  nand2 gate907(.a(s_51), .b(gate99inter3), .O(gate99inter10));
  nor2  gate908(.a(gate99inter10), .b(gate99inter9), .O(gate99inter11));
  nor2  gate909(.a(gate99inter11), .b(gate99inter6), .O(gate99inter12));
  nand2 gate910(.a(gate99inter12), .b(gate99inter1), .O(G420));
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );

  xor2  gate1009(.a(G359), .b(G28), .O(gate103inter0));
  nand2 gate1010(.a(gate103inter0), .b(s_66), .O(gate103inter1));
  and2  gate1011(.a(G359), .b(G28), .O(gate103inter2));
  inv1  gate1012(.a(s_66), .O(gate103inter3));
  inv1  gate1013(.a(s_67), .O(gate103inter4));
  nand2 gate1014(.a(gate103inter4), .b(gate103inter3), .O(gate103inter5));
  nor2  gate1015(.a(gate103inter5), .b(gate103inter2), .O(gate103inter6));
  inv1  gate1016(.a(G28), .O(gate103inter7));
  inv1  gate1017(.a(G359), .O(gate103inter8));
  nand2 gate1018(.a(gate103inter8), .b(gate103inter7), .O(gate103inter9));
  nand2 gate1019(.a(s_67), .b(gate103inter3), .O(gate103inter10));
  nor2  gate1020(.a(gate103inter10), .b(gate103inter9), .O(gate103inter11));
  nor2  gate1021(.a(gate103inter11), .b(gate103inter6), .O(gate103inter12));
  nand2 gate1022(.a(gate103inter12), .b(gate103inter1), .O(G424));
nand2 gate104( .a(G32), .b(G359), .O(G425) );
nand2 gate105( .a(G362), .b(G363), .O(G426) );
nand2 gate106( .a(G364), .b(G365), .O(G429) );
nand2 gate107( .a(G366), .b(G367), .O(G432) );
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate1079(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate1080(.a(gate116inter0), .b(s_76), .O(gate116inter1));
  and2  gate1081(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate1082(.a(s_76), .O(gate116inter3));
  inv1  gate1083(.a(s_77), .O(gate116inter4));
  nand2 gate1084(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate1085(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate1086(.a(G384), .O(gate116inter7));
  inv1  gate1087(.a(G385), .O(gate116inter8));
  nand2 gate1088(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate1089(.a(s_77), .b(gate116inter3), .O(gate116inter10));
  nor2  gate1090(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate1091(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate1092(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );

  xor2  gate1499(.a(G403), .b(G402), .O(gate125inter0));
  nand2 gate1500(.a(gate125inter0), .b(s_136), .O(gate125inter1));
  and2  gate1501(.a(G403), .b(G402), .O(gate125inter2));
  inv1  gate1502(.a(s_136), .O(gate125inter3));
  inv1  gate1503(.a(s_137), .O(gate125inter4));
  nand2 gate1504(.a(gate125inter4), .b(gate125inter3), .O(gate125inter5));
  nor2  gate1505(.a(gate125inter5), .b(gate125inter2), .O(gate125inter6));
  inv1  gate1506(.a(G402), .O(gate125inter7));
  inv1  gate1507(.a(G403), .O(gate125inter8));
  nand2 gate1508(.a(gate125inter8), .b(gate125inter7), .O(gate125inter9));
  nand2 gate1509(.a(s_137), .b(gate125inter3), .O(gate125inter10));
  nor2  gate1510(.a(gate125inter10), .b(gate125inter9), .O(gate125inter11));
  nor2  gate1511(.a(gate125inter11), .b(gate125inter6), .O(gate125inter12));
  nand2 gate1512(.a(gate125inter12), .b(gate125inter1), .O(G486));
nand2 gate126( .a(G404), .b(G405), .O(G489) );
nand2 gate127( .a(G406), .b(G407), .O(G492) );
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );

  xor2  gate1093(.a(G423), .b(G422), .O(gate135inter0));
  nand2 gate1094(.a(gate135inter0), .b(s_78), .O(gate135inter1));
  and2  gate1095(.a(G423), .b(G422), .O(gate135inter2));
  inv1  gate1096(.a(s_78), .O(gate135inter3));
  inv1  gate1097(.a(s_79), .O(gate135inter4));
  nand2 gate1098(.a(gate135inter4), .b(gate135inter3), .O(gate135inter5));
  nor2  gate1099(.a(gate135inter5), .b(gate135inter2), .O(gate135inter6));
  inv1  gate1100(.a(G422), .O(gate135inter7));
  inv1  gate1101(.a(G423), .O(gate135inter8));
  nand2 gate1102(.a(gate135inter8), .b(gate135inter7), .O(gate135inter9));
  nand2 gate1103(.a(s_79), .b(gate135inter3), .O(gate135inter10));
  nor2  gate1104(.a(gate135inter10), .b(gate135inter9), .O(gate135inter11));
  nor2  gate1105(.a(gate135inter11), .b(gate135inter6), .O(gate135inter12));
  nand2 gate1106(.a(gate135inter12), .b(gate135inter1), .O(G516));
nand2 gate136( .a(G424), .b(G425), .O(G519) );

  xor2  gate827(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate828(.a(gate137inter0), .b(s_40), .O(gate137inter1));
  and2  gate829(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate830(.a(s_40), .O(gate137inter3));
  inv1  gate831(.a(s_41), .O(gate137inter4));
  nand2 gate832(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate833(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate834(.a(G426), .O(gate137inter7));
  inv1  gate835(.a(G429), .O(gate137inter8));
  nand2 gate836(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate837(.a(s_41), .b(gate137inter3), .O(gate137inter10));
  nor2  gate838(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate839(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate840(.a(gate137inter12), .b(gate137inter1), .O(G522));
nand2 gate138( .a(G432), .b(G435), .O(G525) );
nand2 gate139( .a(G438), .b(G441), .O(G528) );
nand2 gate140( .a(G444), .b(G447), .O(G531) );
nand2 gate141( .a(G450), .b(G453), .O(G534) );
nand2 gate142( .a(G456), .b(G459), .O(G537) );
nand2 gate143( .a(G462), .b(G465), .O(G540) );
nand2 gate144( .a(G468), .b(G471), .O(G543) );

  xor2  gate1121(.a(G477), .b(G474), .O(gate145inter0));
  nand2 gate1122(.a(gate145inter0), .b(s_82), .O(gate145inter1));
  and2  gate1123(.a(G477), .b(G474), .O(gate145inter2));
  inv1  gate1124(.a(s_82), .O(gate145inter3));
  inv1  gate1125(.a(s_83), .O(gate145inter4));
  nand2 gate1126(.a(gate145inter4), .b(gate145inter3), .O(gate145inter5));
  nor2  gate1127(.a(gate145inter5), .b(gate145inter2), .O(gate145inter6));
  inv1  gate1128(.a(G474), .O(gate145inter7));
  inv1  gate1129(.a(G477), .O(gate145inter8));
  nand2 gate1130(.a(gate145inter8), .b(gate145inter7), .O(gate145inter9));
  nand2 gate1131(.a(s_83), .b(gate145inter3), .O(gate145inter10));
  nor2  gate1132(.a(gate145inter10), .b(gate145inter9), .O(gate145inter11));
  nor2  gate1133(.a(gate145inter11), .b(gate145inter6), .O(gate145inter12));
  nand2 gate1134(.a(gate145inter12), .b(gate145inter1), .O(G546));
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );

  xor2  gate1639(.a(G495), .b(G492), .O(gate148inter0));
  nand2 gate1640(.a(gate148inter0), .b(s_156), .O(gate148inter1));
  and2  gate1641(.a(G495), .b(G492), .O(gate148inter2));
  inv1  gate1642(.a(s_156), .O(gate148inter3));
  inv1  gate1643(.a(s_157), .O(gate148inter4));
  nand2 gate1644(.a(gate148inter4), .b(gate148inter3), .O(gate148inter5));
  nor2  gate1645(.a(gate148inter5), .b(gate148inter2), .O(gate148inter6));
  inv1  gate1646(.a(G492), .O(gate148inter7));
  inv1  gate1647(.a(G495), .O(gate148inter8));
  nand2 gate1648(.a(gate148inter8), .b(gate148inter7), .O(gate148inter9));
  nand2 gate1649(.a(s_157), .b(gate148inter3), .O(gate148inter10));
  nor2  gate1650(.a(gate148inter10), .b(gate148inter9), .O(gate148inter11));
  nor2  gate1651(.a(gate148inter11), .b(gate148inter6), .O(gate148inter12));
  nand2 gate1652(.a(gate148inter12), .b(gate148inter1), .O(G555));
nand2 gate149( .a(G498), .b(G501), .O(G558) );
nand2 gate150( .a(G504), .b(G507), .O(G561) );
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );
nand2 gate159( .a(G444), .b(G531), .O(G576) );

  xor2  gate1359(.a(G531), .b(G447), .O(gate160inter0));
  nand2 gate1360(.a(gate160inter0), .b(s_116), .O(gate160inter1));
  and2  gate1361(.a(G531), .b(G447), .O(gate160inter2));
  inv1  gate1362(.a(s_116), .O(gate160inter3));
  inv1  gate1363(.a(s_117), .O(gate160inter4));
  nand2 gate1364(.a(gate160inter4), .b(gate160inter3), .O(gate160inter5));
  nor2  gate1365(.a(gate160inter5), .b(gate160inter2), .O(gate160inter6));
  inv1  gate1366(.a(G447), .O(gate160inter7));
  inv1  gate1367(.a(G531), .O(gate160inter8));
  nand2 gate1368(.a(gate160inter8), .b(gate160inter7), .O(gate160inter9));
  nand2 gate1369(.a(s_117), .b(gate160inter3), .O(gate160inter10));
  nor2  gate1370(.a(gate160inter10), .b(gate160inter9), .O(gate160inter11));
  nor2  gate1371(.a(gate160inter11), .b(gate160inter6), .O(gate160inter12));
  nand2 gate1372(.a(gate160inter12), .b(gate160inter1), .O(G577));
nand2 gate161( .a(G450), .b(G534), .O(G578) );

  xor2  gate1597(.a(G534), .b(G453), .O(gate162inter0));
  nand2 gate1598(.a(gate162inter0), .b(s_150), .O(gate162inter1));
  and2  gate1599(.a(G534), .b(G453), .O(gate162inter2));
  inv1  gate1600(.a(s_150), .O(gate162inter3));
  inv1  gate1601(.a(s_151), .O(gate162inter4));
  nand2 gate1602(.a(gate162inter4), .b(gate162inter3), .O(gate162inter5));
  nor2  gate1603(.a(gate162inter5), .b(gate162inter2), .O(gate162inter6));
  inv1  gate1604(.a(G453), .O(gate162inter7));
  inv1  gate1605(.a(G534), .O(gate162inter8));
  nand2 gate1606(.a(gate162inter8), .b(gate162inter7), .O(gate162inter9));
  nand2 gate1607(.a(s_151), .b(gate162inter3), .O(gate162inter10));
  nor2  gate1608(.a(gate162inter10), .b(gate162inter9), .O(gate162inter11));
  nor2  gate1609(.a(gate162inter11), .b(gate162inter6), .O(gate162inter12));
  nand2 gate1610(.a(gate162inter12), .b(gate162inter1), .O(G579));
nand2 gate163( .a(G456), .b(G537), .O(G580) );
nand2 gate164( .a(G459), .b(G537), .O(G581) );

  xor2  gate561(.a(G540), .b(G462), .O(gate165inter0));
  nand2 gate562(.a(gate165inter0), .b(s_2), .O(gate165inter1));
  and2  gate563(.a(G540), .b(G462), .O(gate165inter2));
  inv1  gate564(.a(s_2), .O(gate165inter3));
  inv1  gate565(.a(s_3), .O(gate165inter4));
  nand2 gate566(.a(gate165inter4), .b(gate165inter3), .O(gate165inter5));
  nor2  gate567(.a(gate165inter5), .b(gate165inter2), .O(gate165inter6));
  inv1  gate568(.a(G462), .O(gate165inter7));
  inv1  gate569(.a(G540), .O(gate165inter8));
  nand2 gate570(.a(gate165inter8), .b(gate165inter7), .O(gate165inter9));
  nand2 gate571(.a(s_3), .b(gate165inter3), .O(gate165inter10));
  nor2  gate572(.a(gate165inter10), .b(gate165inter9), .O(gate165inter11));
  nor2  gate573(.a(gate165inter11), .b(gate165inter6), .O(gate165inter12));
  nand2 gate574(.a(gate165inter12), .b(gate165inter1), .O(G582));

  xor2  gate729(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate730(.a(gate166inter0), .b(s_26), .O(gate166inter1));
  and2  gate731(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate732(.a(s_26), .O(gate166inter3));
  inv1  gate733(.a(s_27), .O(gate166inter4));
  nand2 gate734(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate735(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate736(.a(G465), .O(gate166inter7));
  inv1  gate737(.a(G540), .O(gate166inter8));
  nand2 gate738(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate739(.a(s_27), .b(gate166inter3), .O(gate166inter10));
  nor2  gate740(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate741(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate742(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );

  xor2  gate1317(.a(G543), .b(G471), .O(gate168inter0));
  nand2 gate1318(.a(gate168inter0), .b(s_110), .O(gate168inter1));
  and2  gate1319(.a(G543), .b(G471), .O(gate168inter2));
  inv1  gate1320(.a(s_110), .O(gate168inter3));
  inv1  gate1321(.a(s_111), .O(gate168inter4));
  nand2 gate1322(.a(gate168inter4), .b(gate168inter3), .O(gate168inter5));
  nor2  gate1323(.a(gate168inter5), .b(gate168inter2), .O(gate168inter6));
  inv1  gate1324(.a(G471), .O(gate168inter7));
  inv1  gate1325(.a(G543), .O(gate168inter8));
  nand2 gate1326(.a(gate168inter8), .b(gate168inter7), .O(gate168inter9));
  nand2 gate1327(.a(s_111), .b(gate168inter3), .O(gate168inter10));
  nor2  gate1328(.a(gate168inter10), .b(gate168inter9), .O(gate168inter11));
  nor2  gate1329(.a(gate168inter11), .b(gate168inter6), .O(gate168inter12));
  nand2 gate1330(.a(gate168inter12), .b(gate168inter1), .O(G585));
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );

  xor2  gate631(.a(G549), .b(G483), .O(gate172inter0));
  nand2 gate632(.a(gate172inter0), .b(s_12), .O(gate172inter1));
  and2  gate633(.a(G549), .b(G483), .O(gate172inter2));
  inv1  gate634(.a(s_12), .O(gate172inter3));
  inv1  gate635(.a(s_13), .O(gate172inter4));
  nand2 gate636(.a(gate172inter4), .b(gate172inter3), .O(gate172inter5));
  nor2  gate637(.a(gate172inter5), .b(gate172inter2), .O(gate172inter6));
  inv1  gate638(.a(G483), .O(gate172inter7));
  inv1  gate639(.a(G549), .O(gate172inter8));
  nand2 gate640(.a(gate172inter8), .b(gate172inter7), .O(gate172inter9));
  nand2 gate641(.a(s_13), .b(gate172inter3), .O(gate172inter10));
  nor2  gate642(.a(gate172inter10), .b(gate172inter9), .O(gate172inter11));
  nor2  gate643(.a(gate172inter11), .b(gate172inter6), .O(gate172inter12));
  nand2 gate644(.a(gate172inter12), .b(gate172inter1), .O(G589));
nand2 gate173( .a(G486), .b(G552), .O(G590) );

  xor2  gate1779(.a(G552), .b(G489), .O(gate174inter0));
  nand2 gate1780(.a(gate174inter0), .b(s_176), .O(gate174inter1));
  and2  gate1781(.a(G552), .b(G489), .O(gate174inter2));
  inv1  gate1782(.a(s_176), .O(gate174inter3));
  inv1  gate1783(.a(s_177), .O(gate174inter4));
  nand2 gate1784(.a(gate174inter4), .b(gate174inter3), .O(gate174inter5));
  nor2  gate1785(.a(gate174inter5), .b(gate174inter2), .O(gate174inter6));
  inv1  gate1786(.a(G489), .O(gate174inter7));
  inv1  gate1787(.a(G552), .O(gate174inter8));
  nand2 gate1788(.a(gate174inter8), .b(gate174inter7), .O(gate174inter9));
  nand2 gate1789(.a(s_177), .b(gate174inter3), .O(gate174inter10));
  nor2  gate1790(.a(gate174inter10), .b(gate174inter9), .O(gate174inter11));
  nor2  gate1791(.a(gate174inter11), .b(gate174inter6), .O(gate174inter12));
  nand2 gate1792(.a(gate174inter12), .b(gate174inter1), .O(G591));
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );
nand2 gate178( .a(G501), .b(G558), .O(G595) );
nand2 gate179( .a(G504), .b(G561), .O(G596) );
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate1275(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate1276(.a(gate183inter0), .b(s_104), .O(gate183inter1));
  and2  gate1277(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate1278(.a(s_104), .O(gate183inter3));
  inv1  gate1279(.a(s_105), .O(gate183inter4));
  nand2 gate1280(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate1281(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate1282(.a(G516), .O(gate183inter7));
  inv1  gate1283(.a(G567), .O(gate183inter8));
  nand2 gate1284(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate1285(.a(s_105), .b(gate183inter3), .O(gate183inter10));
  nor2  gate1286(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate1287(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate1288(.a(gate183inter12), .b(gate183inter1), .O(G600));

  xor2  gate1247(.a(G567), .b(G519), .O(gate184inter0));
  nand2 gate1248(.a(gate184inter0), .b(s_100), .O(gate184inter1));
  and2  gate1249(.a(G567), .b(G519), .O(gate184inter2));
  inv1  gate1250(.a(s_100), .O(gate184inter3));
  inv1  gate1251(.a(s_101), .O(gate184inter4));
  nand2 gate1252(.a(gate184inter4), .b(gate184inter3), .O(gate184inter5));
  nor2  gate1253(.a(gate184inter5), .b(gate184inter2), .O(gate184inter6));
  inv1  gate1254(.a(G519), .O(gate184inter7));
  inv1  gate1255(.a(G567), .O(gate184inter8));
  nand2 gate1256(.a(gate184inter8), .b(gate184inter7), .O(gate184inter9));
  nand2 gate1257(.a(s_101), .b(gate184inter3), .O(gate184inter10));
  nor2  gate1258(.a(gate184inter10), .b(gate184inter9), .O(gate184inter11));
  nor2  gate1259(.a(gate184inter11), .b(gate184inter6), .O(gate184inter12));
  nand2 gate1260(.a(gate184inter12), .b(gate184inter1), .O(G601));
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );

  xor2  gate1723(.a(G577), .b(G576), .O(gate188inter0));
  nand2 gate1724(.a(gate188inter0), .b(s_168), .O(gate188inter1));
  and2  gate1725(.a(G577), .b(G576), .O(gate188inter2));
  inv1  gate1726(.a(s_168), .O(gate188inter3));
  inv1  gate1727(.a(s_169), .O(gate188inter4));
  nand2 gate1728(.a(gate188inter4), .b(gate188inter3), .O(gate188inter5));
  nor2  gate1729(.a(gate188inter5), .b(gate188inter2), .O(gate188inter6));
  inv1  gate1730(.a(G576), .O(gate188inter7));
  inv1  gate1731(.a(G577), .O(gate188inter8));
  nand2 gate1732(.a(gate188inter8), .b(gate188inter7), .O(gate188inter9));
  nand2 gate1733(.a(s_169), .b(gate188inter3), .O(gate188inter10));
  nor2  gate1734(.a(gate188inter10), .b(gate188inter9), .O(gate188inter11));
  nor2  gate1735(.a(gate188inter11), .b(gate188inter6), .O(gate188inter12));
  nand2 gate1736(.a(gate188inter12), .b(gate188inter1), .O(G617));
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );
nand2 gate193( .a(G586), .b(G587), .O(G642) );
nand2 gate194( .a(G588), .b(G589), .O(G645) );
nand2 gate195( .a(G590), .b(G591), .O(G648) );
nand2 gate196( .a(G592), .b(G593), .O(G651) );

  xor2  gate617(.a(G595), .b(G594), .O(gate197inter0));
  nand2 gate618(.a(gate197inter0), .b(s_10), .O(gate197inter1));
  and2  gate619(.a(G595), .b(G594), .O(gate197inter2));
  inv1  gate620(.a(s_10), .O(gate197inter3));
  inv1  gate621(.a(s_11), .O(gate197inter4));
  nand2 gate622(.a(gate197inter4), .b(gate197inter3), .O(gate197inter5));
  nor2  gate623(.a(gate197inter5), .b(gate197inter2), .O(gate197inter6));
  inv1  gate624(.a(G594), .O(gate197inter7));
  inv1  gate625(.a(G595), .O(gate197inter8));
  nand2 gate626(.a(gate197inter8), .b(gate197inter7), .O(gate197inter9));
  nand2 gate627(.a(s_11), .b(gate197inter3), .O(gate197inter10));
  nor2  gate628(.a(gate197inter10), .b(gate197inter9), .O(gate197inter11));
  nor2  gate629(.a(gate197inter11), .b(gate197inter6), .O(gate197inter12));
  nand2 gate630(.a(gate197inter12), .b(gate197inter1), .O(G654));

  xor2  gate1569(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate1570(.a(gate198inter0), .b(s_146), .O(gate198inter1));
  and2  gate1571(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate1572(.a(s_146), .O(gate198inter3));
  inv1  gate1573(.a(s_147), .O(gate198inter4));
  nand2 gate1574(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate1575(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate1576(.a(G596), .O(gate198inter7));
  inv1  gate1577(.a(G597), .O(gate198inter8));
  nand2 gate1578(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate1579(.a(s_147), .b(gate198inter3), .O(gate198inter10));
  nor2  gate1580(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate1581(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate1582(.a(gate198inter12), .b(gate198inter1), .O(G657));

  xor2  gate1471(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate1472(.a(gate199inter0), .b(s_132), .O(gate199inter1));
  and2  gate1473(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate1474(.a(s_132), .O(gate199inter3));
  inv1  gate1475(.a(s_133), .O(gate199inter4));
  nand2 gate1476(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate1477(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate1478(.a(G598), .O(gate199inter7));
  inv1  gate1479(.a(G599), .O(gate199inter8));
  nand2 gate1480(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate1481(.a(s_133), .b(gate199inter3), .O(gate199inter10));
  nor2  gate1482(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate1483(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate1484(.a(gate199inter12), .b(gate199inter1), .O(G660));
nand2 gate200( .a(G600), .b(G601), .O(G663) );
nand2 gate201( .a(G602), .b(G607), .O(G666) );
nand2 gate202( .a(G612), .b(G617), .O(G669) );

  xor2  gate1163(.a(G612), .b(G602), .O(gate203inter0));
  nand2 gate1164(.a(gate203inter0), .b(s_88), .O(gate203inter1));
  and2  gate1165(.a(G612), .b(G602), .O(gate203inter2));
  inv1  gate1166(.a(s_88), .O(gate203inter3));
  inv1  gate1167(.a(s_89), .O(gate203inter4));
  nand2 gate1168(.a(gate203inter4), .b(gate203inter3), .O(gate203inter5));
  nor2  gate1169(.a(gate203inter5), .b(gate203inter2), .O(gate203inter6));
  inv1  gate1170(.a(G602), .O(gate203inter7));
  inv1  gate1171(.a(G612), .O(gate203inter8));
  nand2 gate1172(.a(gate203inter8), .b(gate203inter7), .O(gate203inter9));
  nand2 gate1173(.a(s_89), .b(gate203inter3), .O(gate203inter10));
  nor2  gate1174(.a(gate203inter10), .b(gate203inter9), .O(gate203inter11));
  nor2  gate1175(.a(gate203inter11), .b(gate203inter6), .O(gate203inter12));
  nand2 gate1176(.a(gate203inter12), .b(gate203inter1), .O(G672));
nand2 gate204( .a(G607), .b(G617), .O(G675) );
nand2 gate205( .a(G622), .b(G627), .O(G678) );
nand2 gate206( .a(G632), .b(G637), .O(G681) );
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );
nand2 gate210( .a(G607), .b(G666), .O(G691) );
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );

  xor2  gate1751(.a(G678), .b(G627), .O(gate218inter0));
  nand2 gate1752(.a(gate218inter0), .b(s_172), .O(gate218inter1));
  and2  gate1753(.a(G678), .b(G627), .O(gate218inter2));
  inv1  gate1754(.a(s_172), .O(gate218inter3));
  inv1  gate1755(.a(s_173), .O(gate218inter4));
  nand2 gate1756(.a(gate218inter4), .b(gate218inter3), .O(gate218inter5));
  nor2  gate1757(.a(gate218inter5), .b(gate218inter2), .O(gate218inter6));
  inv1  gate1758(.a(G627), .O(gate218inter7));
  inv1  gate1759(.a(G678), .O(gate218inter8));
  nand2 gate1760(.a(gate218inter8), .b(gate218inter7), .O(gate218inter9));
  nand2 gate1761(.a(s_173), .b(gate218inter3), .O(gate218inter10));
  nor2  gate1762(.a(gate218inter10), .b(gate218inter9), .O(gate218inter11));
  nor2  gate1763(.a(gate218inter11), .b(gate218inter6), .O(gate218inter12));
  nand2 gate1764(.a(gate218inter12), .b(gate218inter1), .O(G699));

  xor2  gate1667(.a(G681), .b(G632), .O(gate219inter0));
  nand2 gate1668(.a(gate219inter0), .b(s_160), .O(gate219inter1));
  and2  gate1669(.a(G681), .b(G632), .O(gate219inter2));
  inv1  gate1670(.a(s_160), .O(gate219inter3));
  inv1  gate1671(.a(s_161), .O(gate219inter4));
  nand2 gate1672(.a(gate219inter4), .b(gate219inter3), .O(gate219inter5));
  nor2  gate1673(.a(gate219inter5), .b(gate219inter2), .O(gate219inter6));
  inv1  gate1674(.a(G632), .O(gate219inter7));
  inv1  gate1675(.a(G681), .O(gate219inter8));
  nand2 gate1676(.a(gate219inter8), .b(gate219inter7), .O(gate219inter9));
  nand2 gate1677(.a(s_161), .b(gate219inter3), .O(gate219inter10));
  nor2  gate1678(.a(gate219inter10), .b(gate219inter9), .O(gate219inter11));
  nor2  gate1679(.a(gate219inter11), .b(gate219inter6), .O(gate219inter12));
  nand2 gate1680(.a(gate219inter12), .b(gate219inter1), .O(G700));
nand2 gate220( .a(G637), .b(G681), .O(G701) );

  xor2  gate1219(.a(G684), .b(G622), .O(gate221inter0));
  nand2 gate1220(.a(gate221inter0), .b(s_96), .O(gate221inter1));
  and2  gate1221(.a(G684), .b(G622), .O(gate221inter2));
  inv1  gate1222(.a(s_96), .O(gate221inter3));
  inv1  gate1223(.a(s_97), .O(gate221inter4));
  nand2 gate1224(.a(gate221inter4), .b(gate221inter3), .O(gate221inter5));
  nor2  gate1225(.a(gate221inter5), .b(gate221inter2), .O(gate221inter6));
  inv1  gate1226(.a(G622), .O(gate221inter7));
  inv1  gate1227(.a(G684), .O(gate221inter8));
  nand2 gate1228(.a(gate221inter8), .b(gate221inter7), .O(gate221inter9));
  nand2 gate1229(.a(s_97), .b(gate221inter3), .O(gate221inter10));
  nor2  gate1230(.a(gate221inter10), .b(gate221inter9), .O(gate221inter11));
  nor2  gate1231(.a(gate221inter11), .b(gate221inter6), .O(gate221inter12));
  nand2 gate1232(.a(gate221inter12), .b(gate221inter1), .O(G702));
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );
nand2 gate224( .a(G637), .b(G687), .O(G705) );
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate925(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate926(.a(gate227inter0), .b(s_54), .O(gate227inter1));
  and2  gate927(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate928(.a(s_54), .O(gate227inter3));
  inv1  gate929(.a(s_55), .O(gate227inter4));
  nand2 gate930(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate931(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate932(.a(G694), .O(gate227inter7));
  inv1  gate933(.a(G695), .O(gate227inter8));
  nand2 gate934(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate935(.a(s_55), .b(gate227inter3), .O(gate227inter10));
  nor2  gate936(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate937(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate938(.a(gate227inter12), .b(gate227inter1), .O(G712));
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );
nand2 gate231( .a(G702), .b(G703), .O(G724) );
nand2 gate232( .a(G704), .b(G705), .O(G727) );
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );
nand2 gate236( .a(G251), .b(G727), .O(G739) );
nand2 gate237( .a(G254), .b(G706), .O(G742) );
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );
nand2 gate240( .a(G263), .b(G715), .O(G751) );
nand2 gate241( .a(G242), .b(G730), .O(G754) );
nand2 gate242( .a(G718), .b(G730), .O(G755) );
nand2 gate243( .a(G245), .b(G733), .O(G756) );
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );
nand2 gate247( .a(G251), .b(G739), .O(G760) );
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );

  xor2  gate1443(.a(G745), .b(G257), .O(gate251inter0));
  nand2 gate1444(.a(gate251inter0), .b(s_128), .O(gate251inter1));
  and2  gate1445(.a(G745), .b(G257), .O(gate251inter2));
  inv1  gate1446(.a(s_128), .O(gate251inter3));
  inv1  gate1447(.a(s_129), .O(gate251inter4));
  nand2 gate1448(.a(gate251inter4), .b(gate251inter3), .O(gate251inter5));
  nor2  gate1449(.a(gate251inter5), .b(gate251inter2), .O(gate251inter6));
  inv1  gate1450(.a(G257), .O(gate251inter7));
  inv1  gate1451(.a(G745), .O(gate251inter8));
  nand2 gate1452(.a(gate251inter8), .b(gate251inter7), .O(gate251inter9));
  nand2 gate1453(.a(s_129), .b(gate251inter3), .O(gate251inter10));
  nor2  gate1454(.a(gate251inter10), .b(gate251inter9), .O(gate251inter11));
  nor2  gate1455(.a(gate251inter11), .b(gate251inter6), .O(gate251inter12));
  nand2 gate1456(.a(gate251inter12), .b(gate251inter1), .O(G764));

  xor2  gate687(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate688(.a(gate252inter0), .b(s_20), .O(gate252inter1));
  and2  gate689(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate690(.a(s_20), .O(gate252inter3));
  inv1  gate691(.a(s_21), .O(gate252inter4));
  nand2 gate692(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate693(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate694(.a(G709), .O(gate252inter7));
  inv1  gate695(.a(G745), .O(gate252inter8));
  nand2 gate696(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate697(.a(s_21), .b(gate252inter3), .O(gate252inter10));
  nor2  gate698(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate699(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate700(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );

  xor2  gate1177(.a(G757), .b(G756), .O(gate258inter0));
  nand2 gate1178(.a(gate258inter0), .b(s_90), .O(gate258inter1));
  and2  gate1179(.a(G757), .b(G756), .O(gate258inter2));
  inv1  gate1180(.a(s_90), .O(gate258inter3));
  inv1  gate1181(.a(s_91), .O(gate258inter4));
  nand2 gate1182(.a(gate258inter4), .b(gate258inter3), .O(gate258inter5));
  nor2  gate1183(.a(gate258inter5), .b(gate258inter2), .O(gate258inter6));
  inv1  gate1184(.a(G756), .O(gate258inter7));
  inv1  gate1185(.a(G757), .O(gate258inter8));
  nand2 gate1186(.a(gate258inter8), .b(gate258inter7), .O(gate258inter9));
  nand2 gate1187(.a(s_91), .b(gate258inter3), .O(gate258inter10));
  nor2  gate1188(.a(gate258inter10), .b(gate258inter9), .O(gate258inter11));
  nor2  gate1189(.a(gate258inter11), .b(gate258inter6), .O(gate258inter12));
  nand2 gate1190(.a(gate258inter12), .b(gate258inter1), .O(G773));
nand2 gate259( .a(G758), .b(G759), .O(G776) );
nand2 gate260( .a(G760), .b(G761), .O(G779) );
nand2 gate261( .a(G762), .b(G763), .O(G782) );

  xor2  gate1555(.a(G765), .b(G764), .O(gate262inter0));
  nand2 gate1556(.a(gate262inter0), .b(s_144), .O(gate262inter1));
  and2  gate1557(.a(G765), .b(G764), .O(gate262inter2));
  inv1  gate1558(.a(s_144), .O(gate262inter3));
  inv1  gate1559(.a(s_145), .O(gate262inter4));
  nand2 gate1560(.a(gate262inter4), .b(gate262inter3), .O(gate262inter5));
  nor2  gate1561(.a(gate262inter5), .b(gate262inter2), .O(gate262inter6));
  inv1  gate1562(.a(G764), .O(gate262inter7));
  inv1  gate1563(.a(G765), .O(gate262inter8));
  nand2 gate1564(.a(gate262inter8), .b(gate262inter7), .O(gate262inter9));
  nand2 gate1565(.a(s_145), .b(gate262inter3), .O(gate262inter10));
  nor2  gate1566(.a(gate262inter10), .b(gate262inter9), .O(gate262inter11));
  nor2  gate1567(.a(gate262inter11), .b(gate262inter6), .O(gate262inter12));
  nand2 gate1568(.a(gate262inter12), .b(gate262inter1), .O(G785));

  xor2  gate1149(.a(G767), .b(G766), .O(gate263inter0));
  nand2 gate1150(.a(gate263inter0), .b(s_86), .O(gate263inter1));
  and2  gate1151(.a(G767), .b(G766), .O(gate263inter2));
  inv1  gate1152(.a(s_86), .O(gate263inter3));
  inv1  gate1153(.a(s_87), .O(gate263inter4));
  nand2 gate1154(.a(gate263inter4), .b(gate263inter3), .O(gate263inter5));
  nor2  gate1155(.a(gate263inter5), .b(gate263inter2), .O(gate263inter6));
  inv1  gate1156(.a(G766), .O(gate263inter7));
  inv1  gate1157(.a(G767), .O(gate263inter8));
  nand2 gate1158(.a(gate263inter8), .b(gate263inter7), .O(gate263inter9));
  nand2 gate1159(.a(s_87), .b(gate263inter3), .O(gate263inter10));
  nor2  gate1160(.a(gate263inter10), .b(gate263inter9), .O(gate263inter11));
  nor2  gate1161(.a(gate263inter11), .b(gate263inter6), .O(gate263inter12));
  nand2 gate1162(.a(gate263inter12), .b(gate263inter1), .O(G788));
nand2 gate264( .a(G768), .b(G769), .O(G791) );

  xor2  gate603(.a(G770), .b(G642), .O(gate265inter0));
  nand2 gate604(.a(gate265inter0), .b(s_8), .O(gate265inter1));
  and2  gate605(.a(G770), .b(G642), .O(gate265inter2));
  inv1  gate606(.a(s_8), .O(gate265inter3));
  inv1  gate607(.a(s_9), .O(gate265inter4));
  nand2 gate608(.a(gate265inter4), .b(gate265inter3), .O(gate265inter5));
  nor2  gate609(.a(gate265inter5), .b(gate265inter2), .O(gate265inter6));
  inv1  gate610(.a(G642), .O(gate265inter7));
  inv1  gate611(.a(G770), .O(gate265inter8));
  nand2 gate612(.a(gate265inter8), .b(gate265inter7), .O(gate265inter9));
  nand2 gate613(.a(s_9), .b(gate265inter3), .O(gate265inter10));
  nor2  gate614(.a(gate265inter10), .b(gate265inter9), .O(gate265inter11));
  nor2  gate615(.a(gate265inter11), .b(gate265inter6), .O(gate265inter12));
  nand2 gate616(.a(gate265inter12), .b(gate265inter1), .O(G794));
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );
nand2 gate268( .a(G651), .b(G779), .O(G803) );
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );
nand2 gate272( .a(G663), .b(G791), .O(G815) );

  xor2  gate1387(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate1388(.a(gate273inter0), .b(s_120), .O(gate273inter1));
  and2  gate1389(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate1390(.a(s_120), .O(gate273inter3));
  inv1  gate1391(.a(s_121), .O(gate273inter4));
  nand2 gate1392(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate1393(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate1394(.a(G642), .O(gate273inter7));
  inv1  gate1395(.a(G794), .O(gate273inter8));
  nand2 gate1396(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate1397(.a(s_121), .b(gate273inter3), .O(gate273inter10));
  nor2  gate1398(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate1399(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate1400(.a(gate273inter12), .b(gate273inter1), .O(G818));

  xor2  gate1793(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate1794(.a(gate274inter0), .b(s_178), .O(gate274inter1));
  and2  gate1795(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate1796(.a(s_178), .O(gate274inter3));
  inv1  gate1797(.a(s_179), .O(gate274inter4));
  nand2 gate1798(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate1799(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate1800(.a(G770), .O(gate274inter7));
  inv1  gate1801(.a(G794), .O(gate274inter8));
  nand2 gate1802(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate1803(.a(s_179), .b(gate274inter3), .O(gate274inter10));
  nor2  gate1804(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate1805(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate1806(.a(gate274inter12), .b(gate274inter1), .O(G819));
nand2 gate275( .a(G645), .b(G797), .O(G820) );
nand2 gate276( .a(G773), .b(G797), .O(G821) );

  xor2  gate953(.a(G800), .b(G648), .O(gate277inter0));
  nand2 gate954(.a(gate277inter0), .b(s_58), .O(gate277inter1));
  and2  gate955(.a(G800), .b(G648), .O(gate277inter2));
  inv1  gate956(.a(s_58), .O(gate277inter3));
  inv1  gate957(.a(s_59), .O(gate277inter4));
  nand2 gate958(.a(gate277inter4), .b(gate277inter3), .O(gate277inter5));
  nor2  gate959(.a(gate277inter5), .b(gate277inter2), .O(gate277inter6));
  inv1  gate960(.a(G648), .O(gate277inter7));
  inv1  gate961(.a(G800), .O(gate277inter8));
  nand2 gate962(.a(gate277inter8), .b(gate277inter7), .O(gate277inter9));
  nand2 gate963(.a(s_59), .b(gate277inter3), .O(gate277inter10));
  nor2  gate964(.a(gate277inter10), .b(gate277inter9), .O(gate277inter11));
  nor2  gate965(.a(gate277inter11), .b(gate277inter6), .O(gate277inter12));
  nand2 gate966(.a(gate277inter12), .b(gate277inter1), .O(G822));
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate1415(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate1416(.a(gate279inter0), .b(s_124), .O(gate279inter1));
  and2  gate1417(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate1418(.a(s_124), .O(gate279inter3));
  inv1  gate1419(.a(s_125), .O(gate279inter4));
  nand2 gate1420(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate1421(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate1422(.a(G651), .O(gate279inter7));
  inv1  gate1423(.a(G803), .O(gate279inter8));
  nand2 gate1424(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate1425(.a(s_125), .b(gate279inter3), .O(gate279inter10));
  nor2  gate1426(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate1427(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate1428(.a(gate279inter12), .b(gate279inter1), .O(G824));
nand2 gate280( .a(G779), .b(G803), .O(G825) );

  xor2  gate1541(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate1542(.a(gate281inter0), .b(s_142), .O(gate281inter1));
  and2  gate1543(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate1544(.a(s_142), .O(gate281inter3));
  inv1  gate1545(.a(s_143), .O(gate281inter4));
  nand2 gate1546(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate1547(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate1548(.a(G654), .O(gate281inter7));
  inv1  gate1549(.a(G806), .O(gate281inter8));
  nand2 gate1550(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate1551(.a(s_143), .b(gate281inter3), .O(gate281inter10));
  nor2  gate1552(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate1553(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate1554(.a(gate281inter12), .b(gate281inter1), .O(G826));
nand2 gate282( .a(G782), .b(G806), .O(G827) );
nand2 gate283( .a(G657), .b(G809), .O(G828) );

  xor2  gate995(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate996(.a(gate284inter0), .b(s_64), .O(gate284inter1));
  and2  gate997(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate998(.a(s_64), .O(gate284inter3));
  inv1  gate999(.a(s_65), .O(gate284inter4));
  nand2 gate1000(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate1001(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate1002(.a(G785), .O(gate284inter7));
  inv1  gate1003(.a(G809), .O(gate284inter8));
  nand2 gate1004(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate1005(.a(s_65), .b(gate284inter3), .O(gate284inter10));
  nor2  gate1006(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate1007(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate1008(.a(gate284inter12), .b(gate284inter1), .O(G829));

  xor2  gate1303(.a(G812), .b(G660), .O(gate285inter0));
  nand2 gate1304(.a(gate285inter0), .b(s_108), .O(gate285inter1));
  and2  gate1305(.a(G812), .b(G660), .O(gate285inter2));
  inv1  gate1306(.a(s_108), .O(gate285inter3));
  inv1  gate1307(.a(s_109), .O(gate285inter4));
  nand2 gate1308(.a(gate285inter4), .b(gate285inter3), .O(gate285inter5));
  nor2  gate1309(.a(gate285inter5), .b(gate285inter2), .O(gate285inter6));
  inv1  gate1310(.a(G660), .O(gate285inter7));
  inv1  gate1311(.a(G812), .O(gate285inter8));
  nand2 gate1312(.a(gate285inter8), .b(gate285inter7), .O(gate285inter9));
  nand2 gate1313(.a(s_109), .b(gate285inter3), .O(gate285inter10));
  nor2  gate1314(.a(gate285inter10), .b(gate285inter9), .O(gate285inter11));
  nor2  gate1315(.a(gate285inter11), .b(gate285inter6), .O(gate285inter12));
  nand2 gate1316(.a(gate285inter12), .b(gate285inter1), .O(G830));
nand2 gate286( .a(G788), .b(G812), .O(G831) );
nand2 gate287( .a(G663), .b(G815), .O(G832) );
nand2 gate288( .a(G791), .b(G815), .O(G833) );
nand2 gate289( .a(G818), .b(G819), .O(G834) );

  xor2  gate1261(.a(G821), .b(G820), .O(gate290inter0));
  nand2 gate1262(.a(gate290inter0), .b(s_102), .O(gate290inter1));
  and2  gate1263(.a(G821), .b(G820), .O(gate290inter2));
  inv1  gate1264(.a(s_102), .O(gate290inter3));
  inv1  gate1265(.a(s_103), .O(gate290inter4));
  nand2 gate1266(.a(gate290inter4), .b(gate290inter3), .O(gate290inter5));
  nor2  gate1267(.a(gate290inter5), .b(gate290inter2), .O(gate290inter6));
  inv1  gate1268(.a(G820), .O(gate290inter7));
  inv1  gate1269(.a(G821), .O(gate290inter8));
  nand2 gate1270(.a(gate290inter8), .b(gate290inter7), .O(gate290inter9));
  nand2 gate1271(.a(s_103), .b(gate290inter3), .O(gate290inter10));
  nor2  gate1272(.a(gate290inter10), .b(gate290inter9), .O(gate290inter11));
  nor2  gate1273(.a(gate290inter11), .b(gate290inter6), .O(gate290inter12));
  nand2 gate1274(.a(gate290inter12), .b(gate290inter1), .O(G847));
nand2 gate291( .a(G822), .b(G823), .O(G860) );

  xor2  gate547(.a(G825), .b(G824), .O(gate292inter0));
  nand2 gate548(.a(gate292inter0), .b(s_0), .O(gate292inter1));
  and2  gate549(.a(G825), .b(G824), .O(gate292inter2));
  inv1  gate550(.a(s_0), .O(gate292inter3));
  inv1  gate551(.a(s_1), .O(gate292inter4));
  nand2 gate552(.a(gate292inter4), .b(gate292inter3), .O(gate292inter5));
  nor2  gate553(.a(gate292inter5), .b(gate292inter2), .O(gate292inter6));
  inv1  gate554(.a(G824), .O(gate292inter7));
  inv1  gate555(.a(G825), .O(gate292inter8));
  nand2 gate556(.a(gate292inter8), .b(gate292inter7), .O(gate292inter9));
  nand2 gate557(.a(s_1), .b(gate292inter3), .O(gate292inter10));
  nor2  gate558(.a(gate292inter10), .b(gate292inter9), .O(gate292inter11));
  nor2  gate559(.a(gate292inter11), .b(gate292inter6), .O(gate292inter12));
  nand2 gate560(.a(gate292inter12), .b(gate292inter1), .O(G873));

  xor2  gate1457(.a(G829), .b(G828), .O(gate293inter0));
  nand2 gate1458(.a(gate293inter0), .b(s_130), .O(gate293inter1));
  and2  gate1459(.a(G829), .b(G828), .O(gate293inter2));
  inv1  gate1460(.a(s_130), .O(gate293inter3));
  inv1  gate1461(.a(s_131), .O(gate293inter4));
  nand2 gate1462(.a(gate293inter4), .b(gate293inter3), .O(gate293inter5));
  nor2  gate1463(.a(gate293inter5), .b(gate293inter2), .O(gate293inter6));
  inv1  gate1464(.a(G828), .O(gate293inter7));
  inv1  gate1465(.a(G829), .O(gate293inter8));
  nand2 gate1466(.a(gate293inter8), .b(gate293inter7), .O(gate293inter9));
  nand2 gate1467(.a(s_131), .b(gate293inter3), .O(gate293inter10));
  nor2  gate1468(.a(gate293inter10), .b(gate293inter9), .O(gate293inter11));
  nor2  gate1469(.a(gate293inter11), .b(gate293inter6), .O(gate293inter12));
  nand2 gate1470(.a(gate293inter12), .b(gate293inter1), .O(G886));
nand2 gate294( .a(G832), .b(G833), .O(G899) );
nand2 gate295( .a(G830), .b(G831), .O(G912) );

  xor2  gate589(.a(G827), .b(G826), .O(gate296inter0));
  nand2 gate590(.a(gate296inter0), .b(s_6), .O(gate296inter1));
  and2  gate591(.a(G827), .b(G826), .O(gate296inter2));
  inv1  gate592(.a(s_6), .O(gate296inter3));
  inv1  gate593(.a(s_7), .O(gate296inter4));
  nand2 gate594(.a(gate296inter4), .b(gate296inter3), .O(gate296inter5));
  nor2  gate595(.a(gate296inter5), .b(gate296inter2), .O(gate296inter6));
  inv1  gate596(.a(G826), .O(gate296inter7));
  inv1  gate597(.a(G827), .O(gate296inter8));
  nand2 gate598(.a(gate296inter8), .b(gate296inter7), .O(gate296inter9));
  nand2 gate599(.a(s_7), .b(gate296inter3), .O(gate296inter10));
  nor2  gate600(.a(gate296inter10), .b(gate296inter9), .O(gate296inter11));
  nor2  gate601(.a(gate296inter11), .b(gate296inter6), .O(gate296inter12));
  nand2 gate602(.a(gate296inter12), .b(gate296inter1), .O(G925));
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );
nand2 gate387( .a(G1), .b(G1036), .O(G1132) );
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );

  xor2  gate659(.a(G1045), .b(G4), .O(gate390inter0));
  nand2 gate660(.a(gate390inter0), .b(s_16), .O(gate390inter1));
  and2  gate661(.a(G1045), .b(G4), .O(gate390inter2));
  inv1  gate662(.a(s_16), .O(gate390inter3));
  inv1  gate663(.a(s_17), .O(gate390inter4));
  nand2 gate664(.a(gate390inter4), .b(gate390inter3), .O(gate390inter5));
  nor2  gate665(.a(gate390inter5), .b(gate390inter2), .O(gate390inter6));
  inv1  gate666(.a(G4), .O(gate390inter7));
  inv1  gate667(.a(G1045), .O(gate390inter8));
  nand2 gate668(.a(gate390inter8), .b(gate390inter7), .O(gate390inter9));
  nand2 gate669(.a(s_17), .b(gate390inter3), .O(gate390inter10));
  nor2  gate670(.a(gate390inter10), .b(gate390inter9), .O(gate390inter11));
  nor2  gate671(.a(gate390inter11), .b(gate390inter6), .O(gate390inter12));
  nand2 gate672(.a(gate390inter12), .b(gate390inter1), .O(G1141));

  xor2  gate1373(.a(G1048), .b(G5), .O(gate391inter0));
  nand2 gate1374(.a(gate391inter0), .b(s_118), .O(gate391inter1));
  and2  gate1375(.a(G1048), .b(G5), .O(gate391inter2));
  inv1  gate1376(.a(s_118), .O(gate391inter3));
  inv1  gate1377(.a(s_119), .O(gate391inter4));
  nand2 gate1378(.a(gate391inter4), .b(gate391inter3), .O(gate391inter5));
  nor2  gate1379(.a(gate391inter5), .b(gate391inter2), .O(gate391inter6));
  inv1  gate1380(.a(G5), .O(gate391inter7));
  inv1  gate1381(.a(G1048), .O(gate391inter8));
  nand2 gate1382(.a(gate391inter8), .b(gate391inter7), .O(gate391inter9));
  nand2 gate1383(.a(s_119), .b(gate391inter3), .O(gate391inter10));
  nor2  gate1384(.a(gate391inter10), .b(gate391inter9), .O(gate391inter11));
  nor2  gate1385(.a(gate391inter11), .b(gate391inter6), .O(gate391inter12));
  nand2 gate1386(.a(gate391inter12), .b(gate391inter1), .O(G1144));
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );
nand2 gate393( .a(G7), .b(G1054), .O(G1150) );
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );

  xor2  gate1653(.a(G1075), .b(G14), .O(gate400inter0));
  nand2 gate1654(.a(gate400inter0), .b(s_158), .O(gate400inter1));
  and2  gate1655(.a(G1075), .b(G14), .O(gate400inter2));
  inv1  gate1656(.a(s_158), .O(gate400inter3));
  inv1  gate1657(.a(s_159), .O(gate400inter4));
  nand2 gate1658(.a(gate400inter4), .b(gate400inter3), .O(gate400inter5));
  nor2  gate1659(.a(gate400inter5), .b(gate400inter2), .O(gate400inter6));
  inv1  gate1660(.a(G14), .O(gate400inter7));
  inv1  gate1661(.a(G1075), .O(gate400inter8));
  nand2 gate1662(.a(gate400inter8), .b(gate400inter7), .O(gate400inter9));
  nand2 gate1663(.a(s_159), .b(gate400inter3), .O(gate400inter10));
  nor2  gate1664(.a(gate400inter10), .b(gate400inter9), .O(gate400inter11));
  nor2  gate1665(.a(gate400inter11), .b(gate400inter6), .O(gate400inter12));
  nand2 gate1666(.a(gate400inter12), .b(gate400inter1), .O(G1171));
nand2 gate401( .a(G15), .b(G1078), .O(G1174) );
nand2 gate402( .a(G16), .b(G1081), .O(G1177) );

  xor2  gate1513(.a(G1084), .b(G17), .O(gate403inter0));
  nand2 gate1514(.a(gate403inter0), .b(s_138), .O(gate403inter1));
  and2  gate1515(.a(G1084), .b(G17), .O(gate403inter2));
  inv1  gate1516(.a(s_138), .O(gate403inter3));
  inv1  gate1517(.a(s_139), .O(gate403inter4));
  nand2 gate1518(.a(gate403inter4), .b(gate403inter3), .O(gate403inter5));
  nor2  gate1519(.a(gate403inter5), .b(gate403inter2), .O(gate403inter6));
  inv1  gate1520(.a(G17), .O(gate403inter7));
  inv1  gate1521(.a(G1084), .O(gate403inter8));
  nand2 gate1522(.a(gate403inter8), .b(gate403inter7), .O(gate403inter9));
  nand2 gate1523(.a(s_139), .b(gate403inter3), .O(gate403inter10));
  nor2  gate1524(.a(gate403inter10), .b(gate403inter9), .O(gate403inter11));
  nor2  gate1525(.a(gate403inter11), .b(gate403inter6), .O(gate403inter12));
  nand2 gate1526(.a(gate403inter12), .b(gate403inter1), .O(G1180));
nand2 gate404( .a(G18), .b(G1087), .O(G1183) );
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );

  xor2  gate575(.a(G1096), .b(G21), .O(gate407inter0));
  nand2 gate576(.a(gate407inter0), .b(s_4), .O(gate407inter1));
  and2  gate577(.a(G1096), .b(G21), .O(gate407inter2));
  inv1  gate578(.a(s_4), .O(gate407inter3));
  inv1  gate579(.a(s_5), .O(gate407inter4));
  nand2 gate580(.a(gate407inter4), .b(gate407inter3), .O(gate407inter5));
  nor2  gate581(.a(gate407inter5), .b(gate407inter2), .O(gate407inter6));
  inv1  gate582(.a(G21), .O(gate407inter7));
  inv1  gate583(.a(G1096), .O(gate407inter8));
  nand2 gate584(.a(gate407inter8), .b(gate407inter7), .O(gate407inter9));
  nand2 gate585(.a(s_5), .b(gate407inter3), .O(gate407inter10));
  nor2  gate586(.a(gate407inter10), .b(gate407inter9), .O(gate407inter11));
  nor2  gate587(.a(gate407inter11), .b(gate407inter6), .O(gate407inter12));
  nand2 gate588(.a(gate407inter12), .b(gate407inter1), .O(G1192));

  xor2  gate1037(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate1038(.a(gate408inter0), .b(s_70), .O(gate408inter1));
  and2  gate1039(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate1040(.a(s_70), .O(gate408inter3));
  inv1  gate1041(.a(s_71), .O(gate408inter4));
  nand2 gate1042(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate1043(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate1044(.a(G22), .O(gate408inter7));
  inv1  gate1045(.a(G1099), .O(gate408inter8));
  nand2 gate1046(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate1047(.a(s_71), .b(gate408inter3), .O(gate408inter10));
  nor2  gate1048(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate1049(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate1050(.a(gate408inter12), .b(gate408inter1), .O(G1195));
nand2 gate409( .a(G23), .b(G1102), .O(G1198) );
nand2 gate410( .a(G24), .b(G1105), .O(G1201) );
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );
nand2 gate412( .a(G26), .b(G1111), .O(G1207) );
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );
nand2 gate415( .a(G29), .b(G1120), .O(G1216) );
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );
nand2 gate417( .a(G31), .b(G1126), .O(G1222) );

  xor2  gate1611(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate1612(.a(gate418inter0), .b(s_152), .O(gate418inter1));
  and2  gate1613(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate1614(.a(s_152), .O(gate418inter3));
  inv1  gate1615(.a(s_153), .O(gate418inter4));
  nand2 gate1616(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate1617(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate1618(.a(G32), .O(gate418inter7));
  inv1  gate1619(.a(G1129), .O(gate418inter8));
  nand2 gate1620(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate1621(.a(s_153), .b(gate418inter3), .O(gate418inter10));
  nor2  gate1622(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate1623(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate1624(.a(gate418inter12), .b(gate418inter1), .O(G1225));
nand2 gate419( .a(G1), .b(G1132), .O(G1228) );
nand2 gate420( .a(G1036), .b(G1132), .O(G1229) );
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );

  xor2  gate1485(.a(G1135), .b(G1039), .O(gate422inter0));
  nand2 gate1486(.a(gate422inter0), .b(s_134), .O(gate422inter1));
  and2  gate1487(.a(G1135), .b(G1039), .O(gate422inter2));
  inv1  gate1488(.a(s_134), .O(gate422inter3));
  inv1  gate1489(.a(s_135), .O(gate422inter4));
  nand2 gate1490(.a(gate422inter4), .b(gate422inter3), .O(gate422inter5));
  nor2  gate1491(.a(gate422inter5), .b(gate422inter2), .O(gate422inter6));
  inv1  gate1492(.a(G1039), .O(gate422inter7));
  inv1  gate1493(.a(G1135), .O(gate422inter8));
  nand2 gate1494(.a(gate422inter8), .b(gate422inter7), .O(gate422inter9));
  nand2 gate1495(.a(s_135), .b(gate422inter3), .O(gate422inter10));
  nor2  gate1496(.a(gate422inter10), .b(gate422inter9), .O(gate422inter11));
  nor2  gate1497(.a(gate422inter11), .b(gate422inter6), .O(gate422inter12));
  nand2 gate1498(.a(gate422inter12), .b(gate422inter1), .O(G1231));
nand2 gate423( .a(G3), .b(G1138), .O(G1232) );

  xor2  gate841(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate842(.a(gate424inter0), .b(s_42), .O(gate424inter1));
  and2  gate843(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate844(.a(s_42), .O(gate424inter3));
  inv1  gate845(.a(s_43), .O(gate424inter4));
  nand2 gate846(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate847(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate848(.a(G1042), .O(gate424inter7));
  inv1  gate849(.a(G1138), .O(gate424inter8));
  nand2 gate850(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate851(.a(s_43), .b(gate424inter3), .O(gate424inter10));
  nor2  gate852(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate853(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate854(.a(gate424inter12), .b(gate424inter1), .O(G1233));
nand2 gate425( .a(G4), .b(G1141), .O(G1234) );
nand2 gate426( .a(G1045), .b(G1141), .O(G1235) );
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );
nand2 gate433( .a(G8), .b(G1153), .O(G1242) );
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );

  xor2  gate1051(.a(G1156), .b(G9), .O(gate435inter0));
  nand2 gate1052(.a(gate435inter0), .b(s_72), .O(gate435inter1));
  and2  gate1053(.a(G1156), .b(G9), .O(gate435inter2));
  inv1  gate1054(.a(s_72), .O(gate435inter3));
  inv1  gate1055(.a(s_73), .O(gate435inter4));
  nand2 gate1056(.a(gate435inter4), .b(gate435inter3), .O(gate435inter5));
  nor2  gate1057(.a(gate435inter5), .b(gate435inter2), .O(gate435inter6));
  inv1  gate1058(.a(G9), .O(gate435inter7));
  inv1  gate1059(.a(G1156), .O(gate435inter8));
  nand2 gate1060(.a(gate435inter8), .b(gate435inter7), .O(gate435inter9));
  nand2 gate1061(.a(s_73), .b(gate435inter3), .O(gate435inter10));
  nor2  gate1062(.a(gate435inter10), .b(gate435inter9), .O(gate435inter11));
  nor2  gate1063(.a(gate435inter11), .b(gate435inter6), .O(gate435inter12));
  nand2 gate1064(.a(gate435inter12), .b(gate435inter1), .O(G1244));
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );

  xor2  gate1023(.a(G1162), .b(G11), .O(gate439inter0));
  nand2 gate1024(.a(gate439inter0), .b(s_68), .O(gate439inter1));
  and2  gate1025(.a(G1162), .b(G11), .O(gate439inter2));
  inv1  gate1026(.a(s_68), .O(gate439inter3));
  inv1  gate1027(.a(s_69), .O(gate439inter4));
  nand2 gate1028(.a(gate439inter4), .b(gate439inter3), .O(gate439inter5));
  nor2  gate1029(.a(gate439inter5), .b(gate439inter2), .O(gate439inter6));
  inv1  gate1030(.a(G11), .O(gate439inter7));
  inv1  gate1031(.a(G1162), .O(gate439inter8));
  nand2 gate1032(.a(gate439inter8), .b(gate439inter7), .O(gate439inter9));
  nand2 gate1033(.a(s_69), .b(gate439inter3), .O(gate439inter10));
  nor2  gate1034(.a(gate439inter10), .b(gate439inter9), .O(gate439inter11));
  nor2  gate1035(.a(gate439inter11), .b(gate439inter6), .O(gate439inter12));
  nand2 gate1036(.a(gate439inter12), .b(gate439inter1), .O(G1248));
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );

  xor2  gate1289(.a(G1165), .b(G12), .O(gate441inter0));
  nand2 gate1290(.a(gate441inter0), .b(s_106), .O(gate441inter1));
  and2  gate1291(.a(G1165), .b(G12), .O(gate441inter2));
  inv1  gate1292(.a(s_106), .O(gate441inter3));
  inv1  gate1293(.a(s_107), .O(gate441inter4));
  nand2 gate1294(.a(gate441inter4), .b(gate441inter3), .O(gate441inter5));
  nor2  gate1295(.a(gate441inter5), .b(gate441inter2), .O(gate441inter6));
  inv1  gate1296(.a(G12), .O(gate441inter7));
  inv1  gate1297(.a(G1165), .O(gate441inter8));
  nand2 gate1298(.a(gate441inter8), .b(gate441inter7), .O(gate441inter9));
  nand2 gate1299(.a(s_107), .b(gate441inter3), .O(gate441inter10));
  nor2  gate1300(.a(gate441inter10), .b(gate441inter9), .O(gate441inter11));
  nor2  gate1301(.a(gate441inter11), .b(gate441inter6), .O(gate441inter12));
  nand2 gate1302(.a(gate441inter12), .b(gate441inter1), .O(G1250));

  xor2  gate1695(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate1696(.a(gate442inter0), .b(s_164), .O(gate442inter1));
  and2  gate1697(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate1698(.a(s_164), .O(gate442inter3));
  inv1  gate1699(.a(s_165), .O(gate442inter4));
  nand2 gate1700(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate1701(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate1702(.a(G1069), .O(gate442inter7));
  inv1  gate1703(.a(G1165), .O(gate442inter8));
  nand2 gate1704(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate1705(.a(s_165), .b(gate442inter3), .O(gate442inter10));
  nor2  gate1706(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate1707(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate1708(.a(gate442inter12), .b(gate442inter1), .O(G1251));

  xor2  gate1681(.a(G1168), .b(G13), .O(gate443inter0));
  nand2 gate1682(.a(gate443inter0), .b(s_162), .O(gate443inter1));
  and2  gate1683(.a(G1168), .b(G13), .O(gate443inter2));
  inv1  gate1684(.a(s_162), .O(gate443inter3));
  inv1  gate1685(.a(s_163), .O(gate443inter4));
  nand2 gate1686(.a(gate443inter4), .b(gate443inter3), .O(gate443inter5));
  nor2  gate1687(.a(gate443inter5), .b(gate443inter2), .O(gate443inter6));
  inv1  gate1688(.a(G13), .O(gate443inter7));
  inv1  gate1689(.a(G1168), .O(gate443inter8));
  nand2 gate1690(.a(gate443inter8), .b(gate443inter7), .O(gate443inter9));
  nand2 gate1691(.a(s_163), .b(gate443inter3), .O(gate443inter10));
  nor2  gate1692(.a(gate443inter10), .b(gate443inter9), .O(gate443inter11));
  nor2  gate1693(.a(gate443inter11), .b(gate443inter6), .O(gate443inter12));
  nand2 gate1694(.a(gate443inter12), .b(gate443inter1), .O(G1252));
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );

  xor2  gate715(.a(G1171), .b(G1075), .O(gate446inter0));
  nand2 gate716(.a(gate446inter0), .b(s_24), .O(gate446inter1));
  and2  gate717(.a(G1171), .b(G1075), .O(gate446inter2));
  inv1  gate718(.a(s_24), .O(gate446inter3));
  inv1  gate719(.a(s_25), .O(gate446inter4));
  nand2 gate720(.a(gate446inter4), .b(gate446inter3), .O(gate446inter5));
  nor2  gate721(.a(gate446inter5), .b(gate446inter2), .O(gate446inter6));
  inv1  gate722(.a(G1075), .O(gate446inter7));
  inv1  gate723(.a(G1171), .O(gate446inter8));
  nand2 gate724(.a(gate446inter8), .b(gate446inter7), .O(gate446inter9));
  nand2 gate725(.a(s_25), .b(gate446inter3), .O(gate446inter10));
  nor2  gate726(.a(gate446inter10), .b(gate446inter9), .O(gate446inter11));
  nor2  gate727(.a(gate446inter11), .b(gate446inter6), .O(gate446inter12));
  nand2 gate728(.a(gate446inter12), .b(gate446inter1), .O(G1255));
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );
nand2 gate449( .a(G16), .b(G1177), .O(G1258) );
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );

  xor2  gate1709(.a(G1183), .b(G18), .O(gate453inter0));
  nand2 gate1710(.a(gate453inter0), .b(s_166), .O(gate453inter1));
  and2  gate1711(.a(G1183), .b(G18), .O(gate453inter2));
  inv1  gate1712(.a(s_166), .O(gate453inter3));
  inv1  gate1713(.a(s_167), .O(gate453inter4));
  nand2 gate1714(.a(gate453inter4), .b(gate453inter3), .O(gate453inter5));
  nor2  gate1715(.a(gate453inter5), .b(gate453inter2), .O(gate453inter6));
  inv1  gate1716(.a(G18), .O(gate453inter7));
  inv1  gate1717(.a(G1183), .O(gate453inter8));
  nand2 gate1718(.a(gate453inter8), .b(gate453inter7), .O(gate453inter9));
  nand2 gate1719(.a(s_167), .b(gate453inter3), .O(gate453inter10));
  nor2  gate1720(.a(gate453inter10), .b(gate453inter9), .O(gate453inter11));
  nor2  gate1721(.a(gate453inter11), .b(gate453inter6), .O(gate453inter12));
  nand2 gate1722(.a(gate453inter12), .b(gate453inter1), .O(G1262));
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );
nand2 gate455( .a(G19), .b(G1186), .O(G1264) );
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );
nand2 gate459( .a(G21), .b(G1192), .O(G1268) );
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );
nand2 gate461( .a(G22), .b(G1195), .O(G1270) );
nand2 gate462( .a(G1099), .b(G1195), .O(G1271) );

  xor2  gate785(.a(G1198), .b(G23), .O(gate463inter0));
  nand2 gate786(.a(gate463inter0), .b(s_34), .O(gate463inter1));
  and2  gate787(.a(G1198), .b(G23), .O(gate463inter2));
  inv1  gate788(.a(s_34), .O(gate463inter3));
  inv1  gate789(.a(s_35), .O(gate463inter4));
  nand2 gate790(.a(gate463inter4), .b(gate463inter3), .O(gate463inter5));
  nor2  gate791(.a(gate463inter5), .b(gate463inter2), .O(gate463inter6));
  inv1  gate792(.a(G23), .O(gate463inter7));
  inv1  gate793(.a(G1198), .O(gate463inter8));
  nand2 gate794(.a(gate463inter8), .b(gate463inter7), .O(gate463inter9));
  nand2 gate795(.a(s_35), .b(gate463inter3), .O(gate463inter10));
  nor2  gate796(.a(gate463inter10), .b(gate463inter9), .O(gate463inter11));
  nor2  gate797(.a(gate463inter11), .b(gate463inter6), .O(gate463inter12));
  nand2 gate798(.a(gate463inter12), .b(gate463inter1), .O(G1272));

  xor2  gate1233(.a(G1198), .b(G1102), .O(gate464inter0));
  nand2 gate1234(.a(gate464inter0), .b(s_98), .O(gate464inter1));
  and2  gate1235(.a(G1198), .b(G1102), .O(gate464inter2));
  inv1  gate1236(.a(s_98), .O(gate464inter3));
  inv1  gate1237(.a(s_99), .O(gate464inter4));
  nand2 gate1238(.a(gate464inter4), .b(gate464inter3), .O(gate464inter5));
  nor2  gate1239(.a(gate464inter5), .b(gate464inter2), .O(gate464inter6));
  inv1  gate1240(.a(G1102), .O(gate464inter7));
  inv1  gate1241(.a(G1198), .O(gate464inter8));
  nand2 gate1242(.a(gate464inter8), .b(gate464inter7), .O(gate464inter9));
  nand2 gate1243(.a(s_99), .b(gate464inter3), .O(gate464inter10));
  nor2  gate1244(.a(gate464inter10), .b(gate464inter9), .O(gate464inter11));
  nor2  gate1245(.a(gate464inter11), .b(gate464inter6), .O(gate464inter12));
  nand2 gate1246(.a(gate464inter12), .b(gate464inter1), .O(G1273));
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate743(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate744(.a(gate466inter0), .b(s_28), .O(gate466inter1));
  and2  gate745(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate746(.a(s_28), .O(gate466inter3));
  inv1  gate747(.a(s_29), .O(gate466inter4));
  nand2 gate748(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate749(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate750(.a(G1105), .O(gate466inter7));
  inv1  gate751(.a(G1201), .O(gate466inter8));
  nand2 gate752(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate753(.a(s_29), .b(gate466inter3), .O(gate466inter10));
  nor2  gate754(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate755(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate756(.a(gate466inter12), .b(gate466inter1), .O(G1275));
nand2 gate467( .a(G25), .b(G1204), .O(G1276) );
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );
nand2 gate471( .a(G27), .b(G1210), .O(G1280) );
nand2 gate472( .a(G1114), .b(G1210), .O(G1281) );
nand2 gate473( .a(G28), .b(G1213), .O(G1282) );
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );
nand2 gate475( .a(G29), .b(G1216), .O(G1284) );
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );
nand2 gate477( .a(G30), .b(G1219), .O(G1286) );

  xor2  gate1807(.a(G1219), .b(G1123), .O(gate478inter0));
  nand2 gate1808(.a(gate478inter0), .b(s_180), .O(gate478inter1));
  and2  gate1809(.a(G1219), .b(G1123), .O(gate478inter2));
  inv1  gate1810(.a(s_180), .O(gate478inter3));
  inv1  gate1811(.a(s_181), .O(gate478inter4));
  nand2 gate1812(.a(gate478inter4), .b(gate478inter3), .O(gate478inter5));
  nor2  gate1813(.a(gate478inter5), .b(gate478inter2), .O(gate478inter6));
  inv1  gate1814(.a(G1123), .O(gate478inter7));
  inv1  gate1815(.a(G1219), .O(gate478inter8));
  nand2 gate1816(.a(gate478inter8), .b(gate478inter7), .O(gate478inter9));
  nand2 gate1817(.a(s_181), .b(gate478inter3), .O(gate478inter10));
  nor2  gate1818(.a(gate478inter10), .b(gate478inter9), .O(gate478inter11));
  nor2  gate1819(.a(gate478inter11), .b(gate478inter6), .O(gate478inter12));
  nand2 gate1820(.a(gate478inter12), .b(gate478inter1), .O(G1287));
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate1135(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate1136(.a(gate480inter0), .b(s_84), .O(gate480inter1));
  and2  gate1137(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate1138(.a(s_84), .O(gate480inter3));
  inv1  gate1139(.a(s_85), .O(gate480inter4));
  nand2 gate1140(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate1141(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate1142(.a(G1126), .O(gate480inter7));
  inv1  gate1143(.a(G1222), .O(gate480inter8));
  nand2 gate1144(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate1145(.a(s_85), .b(gate480inter3), .O(gate480inter10));
  nor2  gate1146(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate1147(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate1148(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );
nand2 gate482( .a(G1129), .b(G1225), .O(G1291) );
nand2 gate483( .a(G1228), .b(G1229), .O(G1292) );
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );

  xor2  gate981(.a(G1233), .b(G1232), .O(gate485inter0));
  nand2 gate982(.a(gate485inter0), .b(s_62), .O(gate485inter1));
  and2  gate983(.a(G1233), .b(G1232), .O(gate485inter2));
  inv1  gate984(.a(s_62), .O(gate485inter3));
  inv1  gate985(.a(s_63), .O(gate485inter4));
  nand2 gate986(.a(gate485inter4), .b(gate485inter3), .O(gate485inter5));
  nor2  gate987(.a(gate485inter5), .b(gate485inter2), .O(gate485inter6));
  inv1  gate988(.a(G1232), .O(gate485inter7));
  inv1  gate989(.a(G1233), .O(gate485inter8));
  nand2 gate990(.a(gate485inter8), .b(gate485inter7), .O(gate485inter9));
  nand2 gate991(.a(s_63), .b(gate485inter3), .O(gate485inter10));
  nor2  gate992(.a(gate485inter10), .b(gate485inter9), .O(gate485inter11));
  nor2  gate993(.a(gate485inter11), .b(gate485inter6), .O(gate485inter12));
  nand2 gate994(.a(gate485inter12), .b(gate485inter1), .O(G1294));

  xor2  gate939(.a(G1235), .b(G1234), .O(gate486inter0));
  nand2 gate940(.a(gate486inter0), .b(s_56), .O(gate486inter1));
  and2  gate941(.a(G1235), .b(G1234), .O(gate486inter2));
  inv1  gate942(.a(s_56), .O(gate486inter3));
  inv1  gate943(.a(s_57), .O(gate486inter4));
  nand2 gate944(.a(gate486inter4), .b(gate486inter3), .O(gate486inter5));
  nor2  gate945(.a(gate486inter5), .b(gate486inter2), .O(gate486inter6));
  inv1  gate946(.a(G1234), .O(gate486inter7));
  inv1  gate947(.a(G1235), .O(gate486inter8));
  nand2 gate948(.a(gate486inter8), .b(gate486inter7), .O(gate486inter9));
  nand2 gate949(.a(s_57), .b(gate486inter3), .O(gate486inter10));
  nor2  gate950(.a(gate486inter10), .b(gate486inter9), .O(gate486inter11));
  nor2  gate951(.a(gate486inter11), .b(gate486inter6), .O(gate486inter12));
  nand2 gate952(.a(gate486inter12), .b(gate486inter1), .O(G1295));
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );
nand2 gate490( .a(G1242), .b(G1243), .O(G1299) );
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );

  xor2  gate799(.a(G1247), .b(G1246), .O(gate492inter0));
  nand2 gate800(.a(gate492inter0), .b(s_36), .O(gate492inter1));
  and2  gate801(.a(G1247), .b(G1246), .O(gate492inter2));
  inv1  gate802(.a(s_36), .O(gate492inter3));
  inv1  gate803(.a(s_37), .O(gate492inter4));
  nand2 gate804(.a(gate492inter4), .b(gate492inter3), .O(gate492inter5));
  nor2  gate805(.a(gate492inter5), .b(gate492inter2), .O(gate492inter6));
  inv1  gate806(.a(G1246), .O(gate492inter7));
  inv1  gate807(.a(G1247), .O(gate492inter8));
  nand2 gate808(.a(gate492inter8), .b(gate492inter7), .O(gate492inter9));
  nand2 gate809(.a(s_37), .b(gate492inter3), .O(gate492inter10));
  nor2  gate810(.a(gate492inter10), .b(gate492inter9), .O(gate492inter11));
  nor2  gate811(.a(gate492inter11), .b(gate492inter6), .O(gate492inter12));
  nand2 gate812(.a(gate492inter12), .b(gate492inter1), .O(G1301));
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );

  xor2  gate855(.a(G1255), .b(G1254), .O(gate496inter0));
  nand2 gate856(.a(gate496inter0), .b(s_44), .O(gate496inter1));
  and2  gate857(.a(G1255), .b(G1254), .O(gate496inter2));
  inv1  gate858(.a(s_44), .O(gate496inter3));
  inv1  gate859(.a(s_45), .O(gate496inter4));
  nand2 gate860(.a(gate496inter4), .b(gate496inter3), .O(gate496inter5));
  nor2  gate861(.a(gate496inter5), .b(gate496inter2), .O(gate496inter6));
  inv1  gate862(.a(G1254), .O(gate496inter7));
  inv1  gate863(.a(G1255), .O(gate496inter8));
  nand2 gate864(.a(gate496inter8), .b(gate496inter7), .O(gate496inter9));
  nand2 gate865(.a(s_45), .b(gate496inter3), .O(gate496inter10));
  nor2  gate866(.a(gate496inter10), .b(gate496inter9), .O(gate496inter11));
  nor2  gate867(.a(gate496inter11), .b(gate496inter6), .O(gate496inter12));
  nand2 gate868(.a(gate496inter12), .b(gate496inter1), .O(G1305));
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );
nand2 gate501( .a(G1264), .b(G1265), .O(G1310) );
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );

  xor2  gate1107(.a(G1271), .b(G1270), .O(gate504inter0));
  nand2 gate1108(.a(gate504inter0), .b(s_80), .O(gate504inter1));
  and2  gate1109(.a(G1271), .b(G1270), .O(gate504inter2));
  inv1  gate1110(.a(s_80), .O(gate504inter3));
  inv1  gate1111(.a(s_81), .O(gate504inter4));
  nand2 gate1112(.a(gate504inter4), .b(gate504inter3), .O(gate504inter5));
  nor2  gate1113(.a(gate504inter5), .b(gate504inter2), .O(gate504inter6));
  inv1  gate1114(.a(G1270), .O(gate504inter7));
  inv1  gate1115(.a(G1271), .O(gate504inter8));
  nand2 gate1116(.a(gate504inter8), .b(gate504inter7), .O(gate504inter9));
  nand2 gate1117(.a(s_81), .b(gate504inter3), .O(gate504inter10));
  nor2  gate1118(.a(gate504inter10), .b(gate504inter9), .O(gate504inter11));
  nor2  gate1119(.a(gate504inter11), .b(gate504inter6), .O(gate504inter12));
  nand2 gate1120(.a(gate504inter12), .b(gate504inter1), .O(G1313));
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );
nand2 gate508( .a(G1278), .b(G1279), .O(G1317) );
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );

  xor2  gate1765(.a(G1283), .b(G1282), .O(gate510inter0));
  nand2 gate1766(.a(gate510inter0), .b(s_174), .O(gate510inter1));
  and2  gate1767(.a(G1283), .b(G1282), .O(gate510inter2));
  inv1  gate1768(.a(s_174), .O(gate510inter3));
  inv1  gate1769(.a(s_175), .O(gate510inter4));
  nand2 gate1770(.a(gate510inter4), .b(gate510inter3), .O(gate510inter5));
  nor2  gate1771(.a(gate510inter5), .b(gate510inter2), .O(gate510inter6));
  inv1  gate1772(.a(G1282), .O(gate510inter7));
  inv1  gate1773(.a(G1283), .O(gate510inter8));
  nand2 gate1774(.a(gate510inter8), .b(gate510inter7), .O(gate510inter9));
  nand2 gate1775(.a(s_175), .b(gate510inter3), .O(gate510inter10));
  nor2  gate1776(.a(gate510inter10), .b(gate510inter9), .O(gate510inter11));
  nor2  gate1777(.a(gate510inter11), .b(gate510inter6), .O(gate510inter12));
  nand2 gate1778(.a(gate510inter12), .b(gate510inter1), .O(G1319));

  xor2  gate1401(.a(G1285), .b(G1284), .O(gate511inter0));
  nand2 gate1402(.a(gate511inter0), .b(s_122), .O(gate511inter1));
  and2  gate1403(.a(G1285), .b(G1284), .O(gate511inter2));
  inv1  gate1404(.a(s_122), .O(gate511inter3));
  inv1  gate1405(.a(s_123), .O(gate511inter4));
  nand2 gate1406(.a(gate511inter4), .b(gate511inter3), .O(gate511inter5));
  nor2  gate1407(.a(gate511inter5), .b(gate511inter2), .O(gate511inter6));
  inv1  gate1408(.a(G1284), .O(gate511inter7));
  inv1  gate1409(.a(G1285), .O(gate511inter8));
  nand2 gate1410(.a(gate511inter8), .b(gate511inter7), .O(gate511inter9));
  nand2 gate1411(.a(s_123), .b(gate511inter3), .O(gate511inter10));
  nor2  gate1412(.a(gate511inter10), .b(gate511inter9), .O(gate511inter11));
  nor2  gate1413(.a(gate511inter11), .b(gate511inter6), .O(gate511inter12));
  nand2 gate1414(.a(gate511inter12), .b(gate511inter1), .O(G1320));
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );
nand2 gate514( .a(G1290), .b(G1291), .O(G1323) );
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule