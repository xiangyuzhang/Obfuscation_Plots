module c1355 (G1, G10, G11, G12, G13, G1324, G1325, G1326, G1327, G1328, G1329, G1330, 
  G1331, G1332, G1333, G1334, G1335, G1336, G1337, G1338, G1339, G1340, G1341, G1342, 
  G1343, G1344, G1345, G1346, G1347, G1348, G1349, G1350, G1351, G1352, G1353, G1354, 
  G1355, G14, G15, G16, G17, G18, G19, G2, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G3, 
  G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G4, G40, G41, G5, G6, G7, G8, G9);
input G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, 
  G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, 
  G40, G41;
  input s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9, s_10, s_11, s_12, s_13, s_14, s_15, s_16, s_17, s_18, s_19, s_20, s_21, s_22, s_23, s_24, s_25, s_26, s_27, s_28, s_29, s_30, s_31, s_32, s_33, s_34, s_35, s_36, s_37, s_38, s_39, s_40, s_41, s_42, s_43, s_44, s_45, s_46, s_47, s_48, s_49, s_50, s_51, s_52, s_53, s_54, s_55, s_56, s_57, s_58, s_59, s_60, s_61, s_62, s_63, s_64, s_65, s_66, s_67, s_68, s_69, s_70, s_71, s_72, s_73, s_74, s_75, s_76, s_77, s_78, s_79, s_80, s_81, s_82, s_83, s_84, s_85, s_86, s_87, s_88, s_89, s_90, s_91, s_92, s_93, s_94, s_95, s_96, s_97, s_98, s_99, s_100, s_101, s_102, s_103, s_104, s_105, s_106, s_107, s_108, s_109, s_110, s_111, s_112, s_113, s_114, s_115, s_116, s_117, s_118, s_119, s_120, s_121, s_122, s_123, s_124, s_125, s_126, s_127, s_128, s_129, s_130, s_131, s_132, s_133, s_134, s_135, s_136, s_137, s_138, s_139, s_140, s_141, s_142, s_143, s_144, s_145, s_146, s_147, s_148, s_149, s_150, s_151, s_152, s_153, s_154, s_155, s_156, s_157, s_158, s_159, s_160, s_161, s_162, s_163, s_164, s_165, s_166, s_167, s_168, s_169, s_170, s_171, s_172, s_173, s_174, s_175, s_176, s_177, s_178, s_179, s_180, s_181, s_182, s_183, s_184, s_185, s_186, s_187, s_188, s_189, s_190, s_191, s_192, s_193, s_194, s_195, s_196, s_197, s_198, s_199, s_200, s_201, s_202, s_203, s_204, s_205, s_206, s_207, s_208, s_209, s_210, s_211, s_212, s_213, s_214, s_215, s_216, s_217, s_218, s_219, s_220, s_221, s_222, s_223, s_224, s_225, s_226, s_227, s_228, s_229, s_230, s_231, s_232, s_233, s_234, s_235, s_236, s_237, s_238, s_239, s_240, s_241, s_242, s_243, s_244, s_245, s_246, s_247, s_248, s_249, s_250, s_251;
output G1324, G1325, G1326, G1327, G1328, G1329, G1330, G1331, G1332, G1333, G1334, G1335, 
  G1336, G1337, G1338, G1339, G1340, G1341, G1342, G1343, G1344, G1345, G1346, G1347, 
  G1348, G1349, G1350, G1351, G1352, G1353, G1354, G1355;
  wire G242, G245, G248, G251, G254, G257, G260, G263, G266, G269, G272, G275, G278, G281, 
    G284, G287, G290, G293, G296, G299, G302, G305, G308, G311, G314, G317, G320, G323, G326, 
    G329, G332, G335, G338, G341, G344, G347, G350, G353, G356, G359, G362, G363, G364, G365, 
    G366, G367, G368, G369, G370, G371, G372, G373, G374, G375, G376, G377, G378, G379, G380, 
    G381, G382, G383, G384, G385, G386, G387, G388, G389, G390, G391, G392, G393, G394, G395, 
    G396, G397, G398, G399, G400, G401, G402, G403, G404, G405, G406, G407, G408, G409, G410, 
    G411, G412, G413, G414, G415, G416, G417, G418, G419, G420, G421, G422, G423, G424, G425, 
    G426, G429, G432, G435, G438, G441, G444, G447, G450, G453, G456, G459, G462, G465, G468, 
    G471, G474, G477, G480, G483, G486, G489, G492, G495, G498, G501, G504, G507, G510, G513, 
    G516, G519, G522, G525, G528, G531, G534, G537, G540, G543, G546, G549, G552, G555, G558, 
    G561, G564, G567, G570, G571, G572, G573, G574, G575, G576, G577, G578, G579, G580, G581, 
    G582, G583, G584, G585, G586, G587, G588, G589, G590, G591, G592, G593, G594, G595, G596, 
    G597, G598, G599, G600, G601, G602, G607, G612, G617, G622, G627, G632, G637, G642, G645, 
    G648, G651, G654, G657, G660, G663, G666, G669, G672, G675, G678, G681, G684, G687, G690, 
    G691, G692, G693, G694, G695, G696, G697, G698, G699, G700, G701, G702, G703, G704, G705, 
    G706, G709, G712, G715, G718, G721, G724, G727, G730, G733, G736, G739, G742, G745, G748, 
    G751, G754, G755, G756, G757, G758, G759, G760, G761, G762, G763, G764, G765, G766, G767, 
    G768, G769, G770, G773, G776, G779, G782, G785, G788, G791, G794, G797, G800, G803, G806, 
    G809, G812, G815, G818, G819, G820, G821, G822, G823, G824, G825, G826, G827, G828, G829, 
    G830, G831, G832, G833, G834, G847, G860, G873, G886, G899, G912, G925, G938, G939, G940, 
    G941, G942, G943, G944, G945, G946, G947, G948, G949, G950, G951, G952, G953, G954, G955, 
    G956, G957, G958, G959, G960, G961, G962, G963, G964, G965, G966, G967, G968, G969, G970, 
    G971, G972, G973, G974, G975, G976, G977, G978, G979, G980, G981, G982, G983, G984, G985, 
    G986, G991, G996, G1001, G1006, G1011, G1016, G1021, G1026, G1031, G1036, G1039, G1042, 
    G1045, G1048, G1051, G1054, G1057, G1060, G1063, G1066, G1069, G1072, G1075, G1078, 
    G1081, G1084, G1087, G1090, G1093, G1096, G1099, G1102, G1105, G1108, G1111, G1114, 
    G1117, G1120, G1123, G1126, G1129, G1132, G1135, G1138, G1141, G1144, G1147, G1150, 
    G1153, G1156, G1159, G1162, G1165, G1168, G1171, G1174, G1177, G1180, G1183, G1186, 
    G1189, G1192, G1195, G1198, G1201, G1204, G1207, G1210, G1213, G1216, G1219, G1222, 
    G1225, G1228, G1229, G1230, G1231, G1232, G1233, G1234, G1235, G1236, G1237, G1238, 
    G1239, G1240, G1241, G1242, G1243, G1244, G1245, G1246, G1247, G1248, G1249, G1250, 
    G1251, G1252, G1253, G1254, G1255, G1256, G1257, G1258, G1259, G1260, G1261, G1262, 
    G1263, G1264, G1265, G1266, G1267, G1268, G1269, G1270, G1271, G1272, G1273, G1274, 
    G1275, G1276, G1277, G1278, G1279, G1280, G1281, G1282, G1283, G1284, G1285, G1286, 
    G1287, G1288, G1289, G1290, G1291, G1292, G1293, G1294, G1295, G1296, G1297, G1298, 
    G1299, G1300, G1301, G1302, G1303, G1304, G1305, G1306, G1307, G1308, G1309, G1310, 
    G1311, G1312, G1313, G1314, G1315, G1316, G1317, G1318, G1319, G1320, G1321, G1322, 
    G1323, gate508inter0, gate508inter1, gate508inter2, gate508inter3, gate508inter4, gate508inter5, gate508inter6, gate508inter7, gate508inter8, gate508inter9, gate508inter10, gate508inter11, gate508inter12, gate116inter0, gate116inter1, gate116inter2, gate116inter3, gate116inter4, gate116inter5, gate116inter6, gate116inter7, gate116inter8, gate116inter9, gate116inter10, gate116inter11, gate116inter12, gate59inter0, gate59inter1, gate59inter2, gate59inter3, gate59inter4, gate59inter5, gate59inter6, gate59inter7, gate59inter8, gate59inter9, gate59inter10, gate59inter11, gate59inter12, gate419inter0, gate419inter1, gate419inter2, gate419inter3, gate419inter4, gate419inter5, gate419inter6, gate419inter7, gate419inter8, gate419inter9, gate419inter10, gate419inter11, gate419inter12, gate159inter0, gate159inter1, gate159inter2, gate159inter3, gate159inter4, gate159inter5, gate159inter6, gate159inter7, gate159inter8, gate159inter9, gate159inter10, gate159inter11, gate159inter12, gate86inter0, gate86inter1, gate86inter2, gate86inter3, gate86inter4, gate86inter5, gate86inter6, gate86inter7, gate86inter8, gate86inter9, gate86inter10, gate86inter11, gate86inter12, gate200inter0, gate200inter1, gate200inter2, gate200inter3, gate200inter4, gate200inter5, gate200inter6, gate200inter7, gate200inter8, gate200inter9, gate200inter10, gate200inter11, gate200inter12, gate16inter0, gate16inter1, gate16inter2, gate16inter3, gate16inter4, gate16inter5, gate16inter6, gate16inter7, gate16inter8, gate16inter9, gate16inter10, gate16inter11, gate16inter12, gate409inter0, gate409inter1, gate409inter2, gate409inter3, gate409inter4, gate409inter5, gate409inter6, gate409inter7, gate409inter8, gate409inter9, gate409inter10, gate409inter11, gate409inter12, gate83inter0, gate83inter1, gate83inter2, gate83inter3, gate83inter4, gate83inter5, gate83inter6, gate83inter7, gate83inter8, gate83inter9, gate83inter10, gate83inter11, gate83inter12, gate105inter0, gate105inter1, gate105inter2, gate105inter3, gate105inter4, gate105inter5, gate105inter6, gate105inter7, gate105inter8, gate105inter9, gate105inter10, gate105inter11, gate105inter12, gate472inter0, gate472inter1, gate472inter2, gate472inter3, gate472inter4, gate472inter5, gate472inter6, gate472inter7, gate472inter8, gate472inter9, gate472inter10, gate472inter11, gate472inter12, gate295inter0, gate295inter1, gate295inter2, gate295inter3, gate295inter4, gate295inter5, gate295inter6, gate295inter7, gate295inter8, gate295inter9, gate295inter10, gate295inter11, gate295inter12, gate418inter0, gate418inter1, gate418inter2, gate418inter3, gate418inter4, gate418inter5, gate418inter6, gate418inter7, gate418inter8, gate418inter9, gate418inter10, gate418inter11, gate418inter12, gate237inter0, gate237inter1, gate237inter2, gate237inter3, gate237inter4, gate237inter5, gate237inter6, gate237inter7, gate237inter8, gate237inter9, gate237inter10, gate237inter11, gate237inter12, gate71inter0, gate71inter1, gate71inter2, gate71inter3, gate71inter4, gate71inter5, gate71inter6, gate71inter7, gate71inter8, gate71inter9, gate71inter10, gate71inter11, gate71inter12, gate287inter0, gate287inter1, gate287inter2, gate287inter3, gate287inter4, gate287inter5, gate287inter6, gate287inter7, gate287inter8, gate287inter9, gate287inter10, gate287inter11, gate287inter12, gate210inter0, gate210inter1, gate210inter2, gate210inter3, gate210inter4, gate210inter5, gate210inter6, gate210inter7, gate210inter8, gate210inter9, gate210inter10, gate210inter11, gate210inter12, gate17inter0, gate17inter1, gate17inter2, gate17inter3, gate17inter4, gate17inter5, gate17inter6, gate17inter7, gate17inter8, gate17inter9, gate17inter10, gate17inter11, gate17inter12, gate466inter0, gate466inter1, gate466inter2, gate466inter3, gate466inter4, gate466inter5, gate466inter6, gate466inter7, gate466inter8, gate466inter9, gate466inter10, gate466inter11, gate466inter12, gate202inter0, gate202inter1, gate202inter2, gate202inter3, gate202inter4, gate202inter5, gate202inter6, gate202inter7, gate202inter8, gate202inter9, gate202inter10, gate202inter11, gate202inter12, gate21inter0, gate21inter1, gate21inter2, gate21inter3, gate21inter4, gate21inter5, gate21inter6, gate21inter7, gate21inter8, gate21inter9, gate21inter10, gate21inter11, gate21inter12, gate106inter0, gate106inter1, gate106inter2, gate106inter3, gate106inter4, gate106inter5, gate106inter6, gate106inter7, gate106inter8, gate106inter9, gate106inter10, gate106inter11, gate106inter12, gate273inter0, gate273inter1, gate273inter2, gate273inter3, gate273inter4, gate273inter5, gate273inter6, gate273inter7, gate273inter8, gate273inter9, gate273inter10, gate273inter11, gate273inter12, gate475inter0, gate475inter1, gate475inter2, gate475inter3, gate475inter4, gate475inter5, gate475inter6, gate475inter7, gate475inter8, gate475inter9, gate475inter10, gate475inter11, gate475inter12, gate442inter0, gate442inter1, gate442inter2, gate442inter3, gate442inter4, gate442inter5, gate442inter6, gate442inter7, gate442inter8, gate442inter9, gate442inter10, gate442inter11, gate442inter12, gate425inter0, gate425inter1, gate425inter2, gate425inter3, gate425inter4, gate425inter5, gate425inter6, gate425inter7, gate425inter8, gate425inter9, gate425inter10, gate425inter11, gate425inter12, gate136inter0, gate136inter1, gate136inter2, gate136inter3, gate136inter4, gate136inter5, gate136inter6, gate136inter7, gate136inter8, gate136inter9, gate136inter10, gate136inter11, gate136inter12, gate9inter0, gate9inter1, gate9inter2, gate9inter3, gate9inter4, gate9inter5, gate9inter6, gate9inter7, gate9inter8, gate9inter9, gate9inter10, gate9inter11, gate9inter12, gate166inter0, gate166inter1, gate166inter2, gate166inter3, gate166inter4, gate166inter5, gate166inter6, gate166inter7, gate166inter8, gate166inter9, gate166inter10, gate166inter11, gate166inter12, gate275inter0, gate275inter1, gate275inter2, gate275inter3, gate275inter4, gate275inter5, gate275inter6, gate275inter7, gate275inter8, gate275inter9, gate275inter10, gate275inter11, gate275inter12, gate179inter0, gate179inter1, gate179inter2, gate179inter3, gate179inter4, gate179inter5, gate179inter6, gate179inter7, gate179inter8, gate179inter9, gate179inter10, gate179inter11, gate179inter12, gate281inter0, gate281inter1, gate281inter2, gate281inter3, gate281inter4, gate281inter5, gate281inter6, gate281inter7, gate281inter8, gate281inter9, gate281inter10, gate281inter11, gate281inter12, gate13inter0, gate13inter1, gate13inter2, gate13inter3, gate13inter4, gate13inter5, gate13inter6, gate13inter7, gate13inter8, gate13inter9, gate13inter10, gate13inter11, gate13inter12, gate426inter0, gate426inter1, gate426inter2, gate426inter3, gate426inter4, gate426inter5, gate426inter6, gate426inter7, gate426inter8, gate426inter9, gate426inter10, gate426inter11, gate426inter12, gate260inter0, gate260inter1, gate260inter2, gate260inter3, gate260inter4, gate260inter5, gate260inter6, gate260inter7, gate260inter8, gate260inter9, gate260inter10, gate260inter11, gate260inter12, gate43inter0, gate43inter1, gate43inter2, gate43inter3, gate43inter4, gate43inter5, gate43inter6, gate43inter7, gate43inter8, gate43inter9, gate43inter10, gate43inter11, gate43inter12, gate514inter0, gate514inter1, gate514inter2, gate514inter3, gate514inter4, gate514inter5, gate514inter6, gate514inter7, gate514inter8, gate514inter9, gate514inter10, gate514inter11, gate514inter12, gate268inter0, gate268inter1, gate268inter2, gate268inter3, gate268inter4, gate268inter5, gate268inter6, gate268inter7, gate268inter8, gate268inter9, gate268inter10, gate268inter11, gate268inter12, gate471inter0, gate471inter1, gate471inter2, gate471inter3, gate471inter4, gate471inter5, gate471inter6, gate471inter7, gate471inter8, gate471inter9, gate471inter10, gate471inter11, gate471inter12, gate53inter0, gate53inter1, gate53inter2, gate53inter3, gate53inter4, gate53inter5, gate53inter6, gate53inter7, gate53inter8, gate53inter9, gate53inter10, gate53inter11, gate53inter12, gate231inter0, gate231inter1, gate231inter2, gate231inter3, gate231inter4, gate231inter5, gate231inter6, gate231inter7, gate231inter8, gate231inter9, gate231inter10, gate231inter11, gate231inter12, gate401inter0, gate401inter1, gate401inter2, gate401inter3, gate401inter4, gate401inter5, gate401inter6, gate401inter7, gate401inter8, gate401inter9, gate401inter10, gate401inter11, gate401inter12, gate417inter0, gate417inter1, gate417inter2, gate417inter3, gate417inter4, gate417inter5, gate417inter6, gate417inter7, gate417inter8, gate417inter9, gate417inter10, gate417inter11, gate417inter12, gate224inter0, gate224inter1, gate224inter2, gate224inter3, gate224inter4, gate224inter5, gate224inter6, gate224inter7, gate224inter8, gate224inter9, gate224inter10, gate224inter11, gate224inter12, gate32inter0, gate32inter1, gate32inter2, gate32inter3, gate32inter4, gate32inter5, gate32inter6, gate32inter7, gate32inter8, gate32inter9, gate32inter10, gate32inter11, gate32inter12, gate227inter0, gate227inter1, gate227inter2, gate227inter3, gate227inter4, gate227inter5, gate227inter6, gate227inter7, gate227inter8, gate227inter9, gate227inter10, gate227inter11, gate227inter12, gate206inter0, gate206inter1, gate206inter2, gate206inter3, gate206inter4, gate206inter5, gate206inter6, gate206inter7, gate206inter8, gate206inter9, gate206inter10, gate206inter11, gate206inter12, gate58inter0, gate58inter1, gate58inter2, gate58inter3, gate58inter4, gate58inter5, gate58inter6, gate58inter7, gate58inter8, gate58inter9, gate58inter10, gate58inter11, gate58inter12, gate27inter0, gate27inter1, gate27inter2, gate27inter3, gate27inter4, gate27inter5, gate27inter6, gate27inter7, gate27inter8, gate27inter9, gate27inter10, gate27inter11, gate27inter12, gate288inter0, gate288inter1, gate288inter2, gate288inter3, gate288inter4, gate288inter5, gate288inter6, gate288inter7, gate288inter8, gate288inter9, gate288inter10, gate288inter11, gate288inter12, gate473inter0, gate473inter1, gate473inter2, gate473inter3, gate473inter4, gate473inter5, gate473inter6, gate473inter7, gate473inter8, gate473inter9, gate473inter10, gate473inter11, gate473inter12, gate173inter0, gate173inter1, gate173inter2, gate173inter3, gate173inter4, gate173inter5, gate173inter6, gate173inter7, gate173inter8, gate173inter9, gate173inter10, gate173inter11, gate173inter12, gate142inter0, gate142inter1, gate142inter2, gate142inter3, gate142inter4, gate142inter5, gate142inter6, gate142inter7, gate142inter8, gate142inter9, gate142inter10, gate142inter11, gate142inter12, gate220inter0, gate220inter1, gate220inter2, gate220inter3, gate220inter4, gate220inter5, gate220inter6, gate220inter7, gate220inter8, gate220inter9, gate220inter10, gate220inter11, gate220inter12, gate272inter0, gate272inter1, gate272inter2, gate272inter3, gate272inter4, gate272inter5, gate272inter6, gate272inter7, gate272inter8, gate272inter9, gate272inter10, gate272inter11, gate272inter12, gate72inter0, gate72inter1, gate72inter2, gate72inter3, gate72inter4, gate72inter5, gate72inter6, gate72inter7, gate72inter8, gate72inter9, gate72inter10, gate72inter11, gate72inter12, gate276inter0, gate276inter1, gate276inter2, gate276inter3, gate276inter4, gate276inter5, gate276inter6, gate276inter7, gate276inter8, gate276inter9, gate276inter10, gate276inter11, gate276inter12, gate240inter0, gate240inter1, gate240inter2, gate240inter3, gate240inter4, gate240inter5, gate240inter6, gate240inter7, gate240inter8, gate240inter9, gate240inter10, gate240inter11, gate240inter12, gate69inter0, gate69inter1, gate69inter2, gate69inter3, gate69inter4, gate69inter5, gate69inter6, gate69inter7, gate69inter8, gate69inter9, gate69inter10, gate69inter11, gate69inter12, gate462inter0, gate462inter1, gate462inter2, gate462inter3, gate462inter4, gate462inter5, gate462inter6, gate462inter7, gate462inter8, gate462inter9, gate462inter10, gate462inter11, gate462inter12, gate73inter0, gate73inter1, gate73inter2, gate73inter3, gate73inter4, gate73inter5, gate73inter6, gate73inter7, gate73inter8, gate73inter9, gate73inter10, gate73inter11, gate73inter12, gate410inter0, gate410inter1, gate410inter2, gate410inter3, gate410inter4, gate410inter5, gate410inter6, gate410inter7, gate410inter8, gate410inter9, gate410inter10, gate410inter11, gate410inter12, gate433inter0, gate433inter1, gate433inter2, gate433inter3, gate433inter4, gate433inter5, gate433inter6, gate433inter7, gate433inter8, gate433inter9, gate433inter10, gate433inter11, gate433inter12, gate31inter0, gate31inter1, gate31inter2, gate31inter3, gate31inter4, gate31inter5, gate31inter6, gate31inter7, gate31inter8, gate31inter9, gate31inter10, gate31inter11, gate31inter12, gate393inter0, gate393inter1, gate393inter2, gate393inter3, gate393inter4, gate393inter5, gate393inter6, gate393inter7, gate393inter8, gate393inter9, gate393inter10, gate393inter11, gate393inter12, gate144inter0, gate144inter1, gate144inter2, gate144inter3, gate144inter4, gate144inter5, gate144inter6, gate144inter7, gate144inter8, gate144inter9, gate144inter10, gate144inter11, gate144inter12, gate449inter0, gate449inter1, gate449inter2, gate449inter3, gate449inter4, gate449inter5, gate449inter6, gate449inter7, gate449inter8, gate449inter9, gate449inter10, gate449inter11, gate449inter12, gate47inter0, gate47inter1, gate47inter2, gate47inter3, gate47inter4, gate47inter5, gate47inter6, gate47inter7, gate47inter8, gate47inter9, gate47inter10, gate47inter11, gate47inter12, gate91inter0, gate91inter1, gate91inter2, gate91inter3, gate91inter4, gate91inter5, gate91inter6, gate91inter7, gate91inter8, gate91inter9, gate91inter10, gate91inter11, gate91inter12, gate76inter0, gate76inter1, gate76inter2, gate76inter3, gate76inter4, gate76inter5, gate76inter6, gate76inter7, gate76inter8, gate76inter9, gate76inter10, gate76inter11, gate76inter12, gate282inter0, gate282inter1, gate282inter2, gate282inter3, gate282inter4, gate282inter5, gate282inter6, gate282inter7, gate282inter8, gate282inter9, gate282inter10, gate282inter11, gate282inter12, gate423inter0, gate423inter1, gate423inter2, gate423inter3, gate423inter4, gate423inter5, gate423inter6, gate423inter7, gate423inter8, gate423inter9, gate423inter10, gate423inter11, gate423inter12, gate501inter0, gate501inter1, gate501inter2, gate501inter3, gate501inter4, gate501inter5, gate501inter6, gate501inter7, gate501inter8, gate501inter9, gate501inter10, gate501inter11, gate501inter12, gate243inter0, gate243inter1, gate243inter2, gate243inter3, gate243inter4, gate243inter5, gate243inter6, gate243inter7, gate243inter8, gate243inter9, gate243inter10, gate243inter11, gate243inter12, gate195inter0, gate195inter1, gate195inter2, gate195inter3, gate195inter4, gate195inter5, gate195inter6, gate195inter7, gate195inter8, gate195inter9, gate195inter10, gate195inter11, gate195inter12, gate236inter0, gate236inter1, gate236inter2, gate236inter3, gate236inter4, gate236inter5, gate236inter6, gate236inter7, gate236inter8, gate236inter9, gate236inter10, gate236inter11, gate236inter12, gate33inter0, gate33inter1, gate33inter2, gate33inter3, gate33inter4, gate33inter5, gate33inter6, gate33inter7, gate33inter8, gate33inter9, gate33inter10, gate33inter11, gate33inter12, gate477inter0, gate477inter1, gate477inter2, gate477inter3, gate477inter4, gate477inter5, gate477inter6, gate477inter7, gate477inter8, gate477inter9, gate477inter10, gate477inter11, gate477inter12, gate150inter0, gate150inter1, gate150inter2, gate150inter3, gate150inter4, gate150inter5, gate150inter6, gate150inter7, gate150inter8, gate150inter9, gate150inter10, gate150inter11, gate150inter12, gate87inter0, gate87inter1, gate87inter2, gate87inter3, gate87inter4, gate87inter5, gate87inter6, gate87inter7, gate87inter8, gate87inter9, gate87inter10, gate87inter11, gate87inter12, gate490inter0, gate490inter1, gate490inter2, gate490inter3, gate490inter4, gate490inter5, gate490inter6, gate490inter7, gate490inter8, gate490inter9, gate490inter10, gate490inter11, gate490inter12, gate482inter0, gate482inter1, gate482inter2, gate482inter3, gate482inter4, gate482inter5, gate482inter6, gate482inter7, gate482inter8, gate482inter9, gate482inter10, gate482inter11, gate482inter12, gate291inter0, gate291inter1, gate291inter2, gate291inter3, gate291inter4, gate291inter5, gate291inter6, gate291inter7, gate291inter8, gate291inter9, gate291inter10, gate291inter11, gate291inter12, gate137inter0, gate137inter1, gate137inter2, gate137inter3, gate137inter4, gate137inter5, gate137inter6, gate137inter7, gate137inter8, gate137inter9, gate137inter10, gate137inter11, gate137inter12, gate459inter0, gate459inter1, gate459inter2, gate459inter3, gate459inter4, gate459inter5, gate459inter6, gate459inter7, gate459inter8, gate459inter9, gate459inter10, gate459inter11, gate459inter12, gate247inter0, gate247inter1, gate247inter2, gate247inter3, gate247inter4, gate247inter5, gate247inter6, gate247inter7, gate247inter8, gate247inter9, gate247inter10, gate247inter11, gate247inter12, gate252inter0, gate252inter1, gate252inter2, gate252inter3, gate252inter4, gate252inter5, gate252inter6, gate252inter7, gate252inter8, gate252inter9, gate252inter10, gate252inter11, gate252inter12, gate198inter0, gate198inter1, gate198inter2, gate198inter3, gate198inter4, gate198inter5, gate198inter6, gate198inter7, gate198inter8, gate198inter9, gate198inter10, gate198inter11, gate198inter12, gate67inter0, gate67inter1, gate67inter2, gate67inter3, gate67inter4, gate67inter5, gate67inter6, gate67inter7, gate67inter8, gate67inter9, gate67inter10, gate67inter11, gate67inter12, gate415inter0, gate415inter1, gate415inter2, gate415inter3, gate415inter4, gate415inter5, gate415inter6, gate415inter7, gate415inter8, gate415inter9, gate415inter10, gate415inter11, gate415inter12, gate261inter0, gate261inter1, gate261inter2, gate261inter3, gate261inter4, gate261inter5, gate261inter6, gate261inter7, gate261inter8, gate261inter9, gate261inter10, gate261inter11, gate261inter12, gate178inter0, gate178inter1, gate178inter2, gate178inter3, gate178inter4, gate178inter5, gate178inter6, gate178inter7, gate178inter8, gate178inter9, gate178inter10, gate178inter11, gate178inter12, gate420inter0, gate420inter1, gate420inter2, gate420inter3, gate420inter4, gate420inter5, gate420inter6, gate420inter7, gate420inter8, gate420inter9, gate420inter10, gate420inter11, gate420inter12, gate138inter0, gate138inter1, gate138inter2, gate138inter3, gate138inter4, gate138inter5, gate138inter6, gate138inter7, gate138inter8, gate138inter9, gate138inter10, gate138inter11, gate138inter12, gate461inter0, gate461inter1, gate461inter2, gate461inter3, gate461inter4, gate461inter5, gate461inter6, gate461inter7, gate461inter8, gate461inter9, gate461inter10, gate461inter11, gate461inter12, gate63inter0, gate63inter1, gate63inter2, gate63inter3, gate63inter4, gate63inter5, gate63inter6, gate63inter7, gate63inter8, gate63inter9, gate63inter10, gate63inter11, gate63inter12, gate483inter0, gate483inter1, gate483inter2, gate483inter3, gate483inter4, gate483inter5, gate483inter6, gate483inter7, gate483inter8, gate483inter9, gate483inter10, gate483inter11, gate483inter12, gate242inter0, gate242inter1, gate242inter2, gate242inter3, gate242inter4, gate242inter5, gate242inter6, gate242inter7, gate242inter8, gate242inter9, gate242inter10, gate242inter11, gate242inter12, gate455inter0, gate455inter1, gate455inter2, gate455inter3, gate455inter4, gate455inter5, gate455inter6, gate455inter7, gate455inter8, gate455inter9, gate455inter10, gate455inter11, gate455inter12, gate279inter0, gate279inter1, gate279inter2, gate279inter3, gate279inter4, gate279inter5, gate279inter6, gate279inter7, gate279inter8, gate279inter9, gate279inter10, gate279inter11, gate279inter12, gate107inter0, gate107inter1, gate107inter2, gate107inter3, gate107inter4, gate107inter5, gate107inter6, gate107inter7, gate107inter8, gate107inter9, gate107inter10, gate107inter11, gate107inter12, gate232inter0, gate232inter1, gate232inter2, gate232inter3, gate232inter4, gate232inter5, gate232inter6, gate232inter7, gate232inter8, gate232inter9, gate232inter10, gate232inter11, gate232inter12, gate424inter0, gate424inter1, gate424inter2, gate424inter3, gate424inter4, gate424inter5, gate424inter6, gate424inter7, gate424inter8, gate424inter9, gate424inter10, gate424inter11, gate424inter12, gate284inter0, gate284inter1, gate284inter2, gate284inter3, gate284inter4, gate284inter5, gate284inter6, gate284inter7, gate284inter8, gate284inter9, gate284inter10, gate284inter11, gate284inter12, gate164inter0, gate164inter1, gate164inter2, gate164inter3, gate164inter4, gate164inter5, gate164inter6, gate164inter7, gate164inter8, gate164inter9, gate164inter10, gate164inter11, gate164inter12, gate387inter0, gate387inter1, gate387inter2, gate387inter3, gate387inter4, gate387inter5, gate387inter6, gate387inter7, gate387inter8, gate387inter9, gate387inter10, gate387inter11, gate387inter12, gate274inter0, gate274inter1, gate274inter2, gate274inter3, gate274inter4, gate274inter5, gate274inter6, gate274inter7, gate274inter8, gate274inter9, gate274inter10, gate274inter11, gate274inter12, gate408inter0, gate408inter1, gate408inter2, gate408inter3, gate408inter4, gate408inter5, gate408inter6, gate408inter7, gate408inter8, gate408inter9, gate408inter10, gate408inter11, gate408inter12, gate404inter0, gate404inter1, gate404inter2, gate404inter3, gate404inter4, gate404inter5, gate404inter6, gate404inter7, gate404inter8, gate404inter9, gate404inter10, gate404inter11, gate404inter12, gate402inter0, gate402inter1, gate402inter2, gate402inter3, gate402inter4, gate402inter5, gate402inter6, gate402inter7, gate402inter8, gate402inter9, gate402inter10, gate402inter11, gate402inter12, gate183inter0, gate183inter1, gate183inter2, gate183inter3, gate183inter4, gate183inter5, gate183inter6, gate183inter7, gate183inter8, gate183inter9, gate183inter10, gate183inter11, gate183inter12, gate412inter0, gate412inter1, gate412inter2, gate412inter3, gate412inter4, gate412inter5, gate412inter6, gate412inter7, gate412inter8, gate412inter9, gate412inter10, gate412inter11, gate412inter12, gate467inter0, gate467inter1, gate467inter2, gate467inter3, gate467inter4, gate467inter5, gate467inter6, gate467inter7, gate467inter8, gate467inter9, gate467inter10, gate467inter11, gate467inter12, gate85inter0, gate85inter1, gate85inter2, gate85inter3, gate85inter4, gate85inter5, gate85inter6, gate85inter7, gate85inter8, gate85inter9, gate85inter10, gate85inter11, gate85inter12, gate127inter0, gate127inter1, gate127inter2, gate127inter3, gate127inter4, gate127inter5, gate127inter6, gate127inter7, gate127inter8, gate127inter9, gate127inter10, gate127inter11, gate127inter12, gate10inter0, gate10inter1, gate10inter2, gate10inter3, gate10inter4, gate10inter5, gate10inter6, gate10inter7, gate10inter8, gate10inter9, gate10inter10, gate10inter11, gate10inter12, gate480inter0, gate480inter1, gate480inter2, gate480inter3, gate480inter4, gate480inter5, gate480inter6, gate480inter7, gate480inter8, gate480inter9, gate480inter10, gate480inter11, gate480inter12, gate280inter0, gate280inter1, gate280inter2, gate280inter3, gate280inter4, gate280inter5, gate280inter6, gate280inter7, gate280inter8, gate280inter9, gate280inter10, gate280inter11, gate280inter12, gate140inter0, gate140inter1, gate140inter2, gate140inter3, gate140inter4, gate140inter5, gate140inter6, gate140inter7, gate140inter8, gate140inter9, gate140inter10, gate140inter11, gate140inter12, gate199inter0, gate199inter1, gate199inter2, gate199inter3, gate199inter4, gate199inter5, gate199inter6, gate199inter7, gate199inter8, gate199inter9, gate199inter10, gate199inter11, gate199inter12, gate193inter0, gate193inter1, gate193inter2, gate193inter3, gate193inter4, gate193inter5, gate193inter6, gate193inter7, gate193inter8, gate193inter9, gate193inter10, gate193inter11, gate193inter12, gate29inter0, gate29inter1, gate29inter2, gate29inter3, gate29inter4, gate29inter5, gate29inter6, gate29inter7, gate29inter8, gate29inter9, gate29inter10, gate29inter11, gate29inter12, gate19inter0, gate19inter1, gate19inter2, gate19inter3, gate19inter4, gate19inter5, gate19inter6, gate19inter7, gate19inter8, gate19inter9, gate19inter10, gate19inter11, gate19inter12, gate92inter0, gate92inter1, gate92inter2, gate92inter3, gate92inter4, gate92inter5, gate92inter6, gate92inter7, gate92inter8, gate92inter9, gate92inter10, gate92inter11, gate92inter12, gate205inter0, gate205inter1, gate205inter2, gate205inter3, gate205inter4, gate205inter5, gate205inter6, gate205inter7, gate205inter8, gate205inter9, gate205inter10, gate205inter11, gate205inter12;


and2 gate1( .a(G33), .b(G41), .O(G242) );
and2 gate2( .a(G34), .b(G41), .O(G245) );
and2 gate3( .a(G35), .b(G41), .O(G248) );
and2 gate4( .a(G36), .b(G41), .O(G251) );
and2 gate5( .a(G37), .b(G41), .O(G254) );
and2 gate6( .a(G38), .b(G41), .O(G257) );
and2 gate7( .a(G39), .b(G41), .O(G260) );
and2 gate8( .a(G40), .b(G41), .O(G263) );

  xor2  gate939(.a(G2), .b(G1), .O(gate9inter0));
  nand2 gate940(.a(gate9inter0), .b(s_56), .O(gate9inter1));
  and2  gate941(.a(G2), .b(G1), .O(gate9inter2));
  inv1  gate942(.a(s_56), .O(gate9inter3));
  inv1  gate943(.a(s_57), .O(gate9inter4));
  nand2 gate944(.a(gate9inter4), .b(gate9inter3), .O(gate9inter5));
  nor2  gate945(.a(gate9inter5), .b(gate9inter2), .O(gate9inter6));
  inv1  gate946(.a(G1), .O(gate9inter7));
  inv1  gate947(.a(G2), .O(gate9inter8));
  nand2 gate948(.a(gate9inter8), .b(gate9inter7), .O(gate9inter9));
  nand2 gate949(.a(s_57), .b(gate9inter3), .O(gate9inter10));
  nor2  gate950(.a(gate9inter10), .b(gate9inter9), .O(gate9inter11));
  nor2  gate951(.a(gate9inter11), .b(gate9inter6), .O(gate9inter12));
  nand2 gate952(.a(gate9inter12), .b(gate9inter1), .O(G266));

  xor2  gate2171(.a(G4), .b(G3), .O(gate10inter0));
  nand2 gate2172(.a(gate10inter0), .b(s_232), .O(gate10inter1));
  and2  gate2173(.a(G4), .b(G3), .O(gate10inter2));
  inv1  gate2174(.a(s_232), .O(gate10inter3));
  inv1  gate2175(.a(s_233), .O(gate10inter4));
  nand2 gate2176(.a(gate10inter4), .b(gate10inter3), .O(gate10inter5));
  nor2  gate2177(.a(gate10inter5), .b(gate10inter2), .O(gate10inter6));
  inv1  gate2178(.a(G3), .O(gate10inter7));
  inv1  gate2179(.a(G4), .O(gate10inter8));
  nand2 gate2180(.a(gate10inter8), .b(gate10inter7), .O(gate10inter9));
  nand2 gate2181(.a(s_233), .b(gate10inter3), .O(gate10inter10));
  nor2  gate2182(.a(gate10inter10), .b(gate10inter9), .O(gate10inter11));
  nor2  gate2183(.a(gate10inter11), .b(gate10inter6), .O(gate10inter12));
  nand2 gate2184(.a(gate10inter12), .b(gate10inter1), .O(G269));
nand2 gate11( .a(G5), .b(G6), .O(G272) );
nand2 gate12( .a(G7), .b(G8), .O(G275) );

  xor2  gate1009(.a(G10), .b(G9), .O(gate13inter0));
  nand2 gate1010(.a(gate13inter0), .b(s_66), .O(gate13inter1));
  and2  gate1011(.a(G10), .b(G9), .O(gate13inter2));
  inv1  gate1012(.a(s_66), .O(gate13inter3));
  inv1  gate1013(.a(s_67), .O(gate13inter4));
  nand2 gate1014(.a(gate13inter4), .b(gate13inter3), .O(gate13inter5));
  nor2  gate1015(.a(gate13inter5), .b(gate13inter2), .O(gate13inter6));
  inv1  gate1016(.a(G9), .O(gate13inter7));
  inv1  gate1017(.a(G10), .O(gate13inter8));
  nand2 gate1018(.a(gate13inter8), .b(gate13inter7), .O(gate13inter9));
  nand2 gate1019(.a(s_67), .b(gate13inter3), .O(gate13inter10));
  nor2  gate1020(.a(gate13inter10), .b(gate13inter9), .O(gate13inter11));
  nor2  gate1021(.a(gate13inter11), .b(gate13inter6), .O(gate13inter12));
  nand2 gate1022(.a(gate13inter12), .b(gate13inter1), .O(G278));
nand2 gate14( .a(G11), .b(G12), .O(G281) );
nand2 gate15( .a(G13), .b(G14), .O(G284) );

  xor2  gate645(.a(G16), .b(G15), .O(gate16inter0));
  nand2 gate646(.a(gate16inter0), .b(s_14), .O(gate16inter1));
  and2  gate647(.a(G16), .b(G15), .O(gate16inter2));
  inv1  gate648(.a(s_14), .O(gate16inter3));
  inv1  gate649(.a(s_15), .O(gate16inter4));
  nand2 gate650(.a(gate16inter4), .b(gate16inter3), .O(gate16inter5));
  nor2  gate651(.a(gate16inter5), .b(gate16inter2), .O(gate16inter6));
  inv1  gate652(.a(G15), .O(gate16inter7));
  inv1  gate653(.a(G16), .O(gate16inter8));
  nand2 gate654(.a(gate16inter8), .b(gate16inter7), .O(gate16inter9));
  nand2 gate655(.a(s_15), .b(gate16inter3), .O(gate16inter10));
  nor2  gate656(.a(gate16inter10), .b(gate16inter9), .O(gate16inter11));
  nor2  gate657(.a(gate16inter11), .b(gate16inter6), .O(gate16inter12));
  nand2 gate658(.a(gate16inter12), .b(gate16inter1), .O(G287));

  xor2  gate799(.a(G18), .b(G17), .O(gate17inter0));
  nand2 gate800(.a(gate17inter0), .b(s_36), .O(gate17inter1));
  and2  gate801(.a(G18), .b(G17), .O(gate17inter2));
  inv1  gate802(.a(s_36), .O(gate17inter3));
  inv1  gate803(.a(s_37), .O(gate17inter4));
  nand2 gate804(.a(gate17inter4), .b(gate17inter3), .O(gate17inter5));
  nor2  gate805(.a(gate17inter5), .b(gate17inter2), .O(gate17inter6));
  inv1  gate806(.a(G17), .O(gate17inter7));
  inv1  gate807(.a(G18), .O(gate17inter8));
  nand2 gate808(.a(gate17inter8), .b(gate17inter7), .O(gate17inter9));
  nand2 gate809(.a(s_37), .b(gate17inter3), .O(gate17inter10));
  nor2  gate810(.a(gate17inter10), .b(gate17inter9), .O(gate17inter11));
  nor2  gate811(.a(gate17inter11), .b(gate17inter6), .O(gate17inter12));
  nand2 gate812(.a(gate17inter12), .b(gate17inter1), .O(G290));
nand2 gate18( .a(G19), .b(G20), .O(G293) );

  xor2  gate2269(.a(G22), .b(G21), .O(gate19inter0));
  nand2 gate2270(.a(gate19inter0), .b(s_246), .O(gate19inter1));
  and2  gate2271(.a(G22), .b(G21), .O(gate19inter2));
  inv1  gate2272(.a(s_246), .O(gate19inter3));
  inv1  gate2273(.a(s_247), .O(gate19inter4));
  nand2 gate2274(.a(gate19inter4), .b(gate19inter3), .O(gate19inter5));
  nor2  gate2275(.a(gate19inter5), .b(gate19inter2), .O(gate19inter6));
  inv1  gate2276(.a(G21), .O(gate19inter7));
  inv1  gate2277(.a(G22), .O(gate19inter8));
  nand2 gate2278(.a(gate19inter8), .b(gate19inter7), .O(gate19inter9));
  nand2 gate2279(.a(s_247), .b(gate19inter3), .O(gate19inter10));
  nor2  gate2280(.a(gate19inter10), .b(gate19inter9), .O(gate19inter11));
  nor2  gate2281(.a(gate19inter11), .b(gate19inter6), .O(gate19inter12));
  nand2 gate2282(.a(gate19inter12), .b(gate19inter1), .O(G296));
nand2 gate20( .a(G23), .b(G24), .O(G299) );

  xor2  gate841(.a(G26), .b(G25), .O(gate21inter0));
  nand2 gate842(.a(gate21inter0), .b(s_42), .O(gate21inter1));
  and2  gate843(.a(G26), .b(G25), .O(gate21inter2));
  inv1  gate844(.a(s_42), .O(gate21inter3));
  inv1  gate845(.a(s_43), .O(gate21inter4));
  nand2 gate846(.a(gate21inter4), .b(gate21inter3), .O(gate21inter5));
  nor2  gate847(.a(gate21inter5), .b(gate21inter2), .O(gate21inter6));
  inv1  gate848(.a(G25), .O(gate21inter7));
  inv1  gate849(.a(G26), .O(gate21inter8));
  nand2 gate850(.a(gate21inter8), .b(gate21inter7), .O(gate21inter9));
  nand2 gate851(.a(s_43), .b(gate21inter3), .O(gate21inter10));
  nor2  gate852(.a(gate21inter10), .b(gate21inter9), .O(gate21inter11));
  nor2  gate853(.a(gate21inter11), .b(gate21inter6), .O(gate21inter12));
  nand2 gate854(.a(gate21inter12), .b(gate21inter1), .O(G302));
nand2 gate22( .a(G27), .b(G28), .O(G305) );
nand2 gate23( .a(G29), .b(G30), .O(G308) );
nand2 gate24( .a(G31), .b(G32), .O(G311) );
nand2 gate25( .a(G1), .b(G5), .O(G314) );
nand2 gate26( .a(G9), .b(G13), .O(G317) );

  xor2  gate1233(.a(G6), .b(G2), .O(gate27inter0));
  nand2 gate1234(.a(gate27inter0), .b(s_98), .O(gate27inter1));
  and2  gate1235(.a(G6), .b(G2), .O(gate27inter2));
  inv1  gate1236(.a(s_98), .O(gate27inter3));
  inv1  gate1237(.a(s_99), .O(gate27inter4));
  nand2 gate1238(.a(gate27inter4), .b(gate27inter3), .O(gate27inter5));
  nor2  gate1239(.a(gate27inter5), .b(gate27inter2), .O(gate27inter6));
  inv1  gate1240(.a(G2), .O(gate27inter7));
  inv1  gate1241(.a(G6), .O(gate27inter8));
  nand2 gate1242(.a(gate27inter8), .b(gate27inter7), .O(gate27inter9));
  nand2 gate1243(.a(s_99), .b(gate27inter3), .O(gate27inter10));
  nor2  gate1244(.a(gate27inter10), .b(gate27inter9), .O(gate27inter11));
  nor2  gate1245(.a(gate27inter11), .b(gate27inter6), .O(gate27inter12));
  nand2 gate1246(.a(gate27inter12), .b(gate27inter1), .O(G320));
nand2 gate28( .a(G10), .b(G14), .O(G323) );

  xor2  gate2255(.a(G7), .b(G3), .O(gate29inter0));
  nand2 gate2256(.a(gate29inter0), .b(s_244), .O(gate29inter1));
  and2  gate2257(.a(G7), .b(G3), .O(gate29inter2));
  inv1  gate2258(.a(s_244), .O(gate29inter3));
  inv1  gate2259(.a(s_245), .O(gate29inter4));
  nand2 gate2260(.a(gate29inter4), .b(gate29inter3), .O(gate29inter5));
  nor2  gate2261(.a(gate29inter5), .b(gate29inter2), .O(gate29inter6));
  inv1  gate2262(.a(G3), .O(gate29inter7));
  inv1  gate2263(.a(G7), .O(gate29inter8));
  nand2 gate2264(.a(gate29inter8), .b(gate29inter7), .O(gate29inter9));
  nand2 gate2265(.a(s_245), .b(gate29inter3), .O(gate29inter10));
  nor2  gate2266(.a(gate29inter10), .b(gate29inter9), .O(gate29inter11));
  nor2  gate2267(.a(gate29inter11), .b(gate29inter6), .O(gate29inter12));
  nand2 gate2268(.a(gate29inter12), .b(gate29inter1), .O(G326));
nand2 gate30( .a(G11), .b(G15), .O(G329) );

  xor2  gate1443(.a(G8), .b(G4), .O(gate31inter0));
  nand2 gate1444(.a(gate31inter0), .b(s_128), .O(gate31inter1));
  and2  gate1445(.a(G8), .b(G4), .O(gate31inter2));
  inv1  gate1446(.a(s_128), .O(gate31inter3));
  inv1  gate1447(.a(s_129), .O(gate31inter4));
  nand2 gate1448(.a(gate31inter4), .b(gate31inter3), .O(gate31inter5));
  nor2  gate1449(.a(gate31inter5), .b(gate31inter2), .O(gate31inter6));
  inv1  gate1450(.a(G4), .O(gate31inter7));
  inv1  gate1451(.a(G8), .O(gate31inter8));
  nand2 gate1452(.a(gate31inter8), .b(gate31inter7), .O(gate31inter9));
  nand2 gate1453(.a(s_129), .b(gate31inter3), .O(gate31inter10));
  nor2  gate1454(.a(gate31inter10), .b(gate31inter9), .O(gate31inter11));
  nor2  gate1455(.a(gate31inter11), .b(gate31inter6), .O(gate31inter12));
  nand2 gate1456(.a(gate31inter12), .b(gate31inter1), .O(G332));

  xor2  gate1177(.a(G16), .b(G12), .O(gate32inter0));
  nand2 gate1178(.a(gate32inter0), .b(s_90), .O(gate32inter1));
  and2  gate1179(.a(G16), .b(G12), .O(gate32inter2));
  inv1  gate1180(.a(s_90), .O(gate32inter3));
  inv1  gate1181(.a(s_91), .O(gate32inter4));
  nand2 gate1182(.a(gate32inter4), .b(gate32inter3), .O(gate32inter5));
  nor2  gate1183(.a(gate32inter5), .b(gate32inter2), .O(gate32inter6));
  inv1  gate1184(.a(G12), .O(gate32inter7));
  inv1  gate1185(.a(G16), .O(gate32inter8));
  nand2 gate1186(.a(gate32inter8), .b(gate32inter7), .O(gate32inter9));
  nand2 gate1187(.a(s_91), .b(gate32inter3), .O(gate32inter10));
  nor2  gate1188(.a(gate32inter10), .b(gate32inter9), .O(gate32inter11));
  nor2  gate1189(.a(gate32inter11), .b(gate32inter6), .O(gate32inter12));
  nand2 gate1190(.a(gate32inter12), .b(gate32inter1), .O(G335));

  xor2  gate1625(.a(G21), .b(G17), .O(gate33inter0));
  nand2 gate1626(.a(gate33inter0), .b(s_154), .O(gate33inter1));
  and2  gate1627(.a(G21), .b(G17), .O(gate33inter2));
  inv1  gate1628(.a(s_154), .O(gate33inter3));
  inv1  gate1629(.a(s_155), .O(gate33inter4));
  nand2 gate1630(.a(gate33inter4), .b(gate33inter3), .O(gate33inter5));
  nor2  gate1631(.a(gate33inter5), .b(gate33inter2), .O(gate33inter6));
  inv1  gate1632(.a(G17), .O(gate33inter7));
  inv1  gate1633(.a(G21), .O(gate33inter8));
  nand2 gate1634(.a(gate33inter8), .b(gate33inter7), .O(gate33inter9));
  nand2 gate1635(.a(s_155), .b(gate33inter3), .O(gate33inter10));
  nor2  gate1636(.a(gate33inter10), .b(gate33inter9), .O(gate33inter11));
  nor2  gate1637(.a(gate33inter11), .b(gate33inter6), .O(gate33inter12));
  nand2 gate1638(.a(gate33inter12), .b(gate33inter1), .O(G338));
nand2 gate34( .a(G25), .b(G29), .O(G341) );
nand2 gate35( .a(G18), .b(G22), .O(G344) );
nand2 gate36( .a(G26), .b(G30), .O(G347) );
nand2 gate37( .a(G19), .b(G23), .O(G350) );
nand2 gate38( .a(G27), .b(G31), .O(G353) );
nand2 gate39( .a(G20), .b(G24), .O(G356) );
nand2 gate40( .a(G28), .b(G32), .O(G359) );
nand2 gate41( .a(G1), .b(G266), .O(G362) );
nand2 gate42( .a(G2), .b(G266), .O(G363) );

  xor2  gate1051(.a(G269), .b(G3), .O(gate43inter0));
  nand2 gate1052(.a(gate43inter0), .b(s_72), .O(gate43inter1));
  and2  gate1053(.a(G269), .b(G3), .O(gate43inter2));
  inv1  gate1054(.a(s_72), .O(gate43inter3));
  inv1  gate1055(.a(s_73), .O(gate43inter4));
  nand2 gate1056(.a(gate43inter4), .b(gate43inter3), .O(gate43inter5));
  nor2  gate1057(.a(gate43inter5), .b(gate43inter2), .O(gate43inter6));
  inv1  gate1058(.a(G3), .O(gate43inter7));
  inv1  gate1059(.a(G269), .O(gate43inter8));
  nand2 gate1060(.a(gate43inter8), .b(gate43inter7), .O(gate43inter9));
  nand2 gate1061(.a(s_73), .b(gate43inter3), .O(gate43inter10));
  nor2  gate1062(.a(gate43inter10), .b(gate43inter9), .O(gate43inter11));
  nor2  gate1063(.a(gate43inter11), .b(gate43inter6), .O(gate43inter12));
  nand2 gate1064(.a(gate43inter12), .b(gate43inter1), .O(G364));
nand2 gate44( .a(G4), .b(G269), .O(G365) );
nand2 gate45( .a(G5), .b(G272), .O(G366) );
nand2 gate46( .a(G6), .b(G272), .O(G367) );

  xor2  gate1499(.a(G275), .b(G7), .O(gate47inter0));
  nand2 gate1500(.a(gate47inter0), .b(s_136), .O(gate47inter1));
  and2  gate1501(.a(G275), .b(G7), .O(gate47inter2));
  inv1  gate1502(.a(s_136), .O(gate47inter3));
  inv1  gate1503(.a(s_137), .O(gate47inter4));
  nand2 gate1504(.a(gate47inter4), .b(gate47inter3), .O(gate47inter5));
  nor2  gate1505(.a(gate47inter5), .b(gate47inter2), .O(gate47inter6));
  inv1  gate1506(.a(G7), .O(gate47inter7));
  inv1  gate1507(.a(G275), .O(gate47inter8));
  nand2 gate1508(.a(gate47inter8), .b(gate47inter7), .O(gate47inter9));
  nand2 gate1509(.a(s_137), .b(gate47inter3), .O(gate47inter10));
  nor2  gate1510(.a(gate47inter10), .b(gate47inter9), .O(gate47inter11));
  nor2  gate1511(.a(gate47inter11), .b(gate47inter6), .O(gate47inter12));
  nand2 gate1512(.a(gate47inter12), .b(gate47inter1), .O(G368));
nand2 gate48( .a(G8), .b(G275), .O(G369) );
nand2 gate49( .a(G9), .b(G278), .O(G370) );
nand2 gate50( .a(G10), .b(G278), .O(G371) );
nand2 gate51( .a(G11), .b(G281), .O(G372) );
nand2 gate52( .a(G12), .b(G281), .O(G373) );

  xor2  gate1107(.a(G284), .b(G13), .O(gate53inter0));
  nand2 gate1108(.a(gate53inter0), .b(s_80), .O(gate53inter1));
  and2  gate1109(.a(G284), .b(G13), .O(gate53inter2));
  inv1  gate1110(.a(s_80), .O(gate53inter3));
  inv1  gate1111(.a(s_81), .O(gate53inter4));
  nand2 gate1112(.a(gate53inter4), .b(gate53inter3), .O(gate53inter5));
  nor2  gate1113(.a(gate53inter5), .b(gate53inter2), .O(gate53inter6));
  inv1  gate1114(.a(G13), .O(gate53inter7));
  inv1  gate1115(.a(G284), .O(gate53inter8));
  nand2 gate1116(.a(gate53inter8), .b(gate53inter7), .O(gate53inter9));
  nand2 gate1117(.a(s_81), .b(gate53inter3), .O(gate53inter10));
  nor2  gate1118(.a(gate53inter10), .b(gate53inter9), .O(gate53inter11));
  nor2  gate1119(.a(gate53inter11), .b(gate53inter6), .O(gate53inter12));
  nand2 gate1120(.a(gate53inter12), .b(gate53inter1), .O(G374));
nand2 gate54( .a(G14), .b(G284), .O(G375) );
nand2 gate55( .a(G15), .b(G287), .O(G376) );
nand2 gate56( .a(G16), .b(G287), .O(G377) );
nand2 gate57( .a(G17), .b(G290), .O(G378) );

  xor2  gate1219(.a(G290), .b(G18), .O(gate58inter0));
  nand2 gate1220(.a(gate58inter0), .b(s_96), .O(gate58inter1));
  and2  gate1221(.a(G290), .b(G18), .O(gate58inter2));
  inv1  gate1222(.a(s_96), .O(gate58inter3));
  inv1  gate1223(.a(s_97), .O(gate58inter4));
  nand2 gate1224(.a(gate58inter4), .b(gate58inter3), .O(gate58inter5));
  nor2  gate1225(.a(gate58inter5), .b(gate58inter2), .O(gate58inter6));
  inv1  gate1226(.a(G18), .O(gate58inter7));
  inv1  gate1227(.a(G290), .O(gate58inter8));
  nand2 gate1228(.a(gate58inter8), .b(gate58inter7), .O(gate58inter9));
  nand2 gate1229(.a(s_97), .b(gate58inter3), .O(gate58inter10));
  nor2  gate1230(.a(gate58inter10), .b(gate58inter9), .O(gate58inter11));
  nor2  gate1231(.a(gate58inter11), .b(gate58inter6), .O(gate58inter12));
  nand2 gate1232(.a(gate58inter12), .b(gate58inter1), .O(G379));

  xor2  gate575(.a(G293), .b(G19), .O(gate59inter0));
  nand2 gate576(.a(gate59inter0), .b(s_4), .O(gate59inter1));
  and2  gate577(.a(G293), .b(G19), .O(gate59inter2));
  inv1  gate578(.a(s_4), .O(gate59inter3));
  inv1  gate579(.a(s_5), .O(gate59inter4));
  nand2 gate580(.a(gate59inter4), .b(gate59inter3), .O(gate59inter5));
  nor2  gate581(.a(gate59inter5), .b(gate59inter2), .O(gate59inter6));
  inv1  gate582(.a(G19), .O(gate59inter7));
  inv1  gate583(.a(G293), .O(gate59inter8));
  nand2 gate584(.a(gate59inter8), .b(gate59inter7), .O(gate59inter9));
  nand2 gate585(.a(s_5), .b(gate59inter3), .O(gate59inter10));
  nor2  gate586(.a(gate59inter10), .b(gate59inter9), .O(gate59inter11));
  nor2  gate587(.a(gate59inter11), .b(gate59inter6), .O(gate59inter12));
  nand2 gate588(.a(gate59inter12), .b(gate59inter1), .O(G380));
nand2 gate60( .a(G20), .b(G293), .O(G381) );
nand2 gate61( .a(G21), .b(G296), .O(G382) );
nand2 gate62( .a(G22), .b(G296), .O(G383) );

  xor2  gate1891(.a(G299), .b(G23), .O(gate63inter0));
  nand2 gate1892(.a(gate63inter0), .b(s_192), .O(gate63inter1));
  and2  gate1893(.a(G299), .b(G23), .O(gate63inter2));
  inv1  gate1894(.a(s_192), .O(gate63inter3));
  inv1  gate1895(.a(s_193), .O(gate63inter4));
  nand2 gate1896(.a(gate63inter4), .b(gate63inter3), .O(gate63inter5));
  nor2  gate1897(.a(gate63inter5), .b(gate63inter2), .O(gate63inter6));
  inv1  gate1898(.a(G23), .O(gate63inter7));
  inv1  gate1899(.a(G299), .O(gate63inter8));
  nand2 gate1900(.a(gate63inter8), .b(gate63inter7), .O(gate63inter9));
  nand2 gate1901(.a(s_193), .b(gate63inter3), .O(gate63inter10));
  nor2  gate1902(.a(gate63inter10), .b(gate63inter9), .O(gate63inter11));
  nor2  gate1903(.a(gate63inter11), .b(gate63inter6), .O(gate63inter12));
  nand2 gate1904(.a(gate63inter12), .b(gate63inter1), .O(G384));
nand2 gate64( .a(G24), .b(G299), .O(G385) );
nand2 gate65( .a(G25), .b(G302), .O(G386) );
nand2 gate66( .a(G26), .b(G302), .O(G387) );

  xor2  gate1793(.a(G305), .b(G27), .O(gate67inter0));
  nand2 gate1794(.a(gate67inter0), .b(s_178), .O(gate67inter1));
  and2  gate1795(.a(G305), .b(G27), .O(gate67inter2));
  inv1  gate1796(.a(s_178), .O(gate67inter3));
  inv1  gate1797(.a(s_179), .O(gate67inter4));
  nand2 gate1798(.a(gate67inter4), .b(gate67inter3), .O(gate67inter5));
  nor2  gate1799(.a(gate67inter5), .b(gate67inter2), .O(gate67inter6));
  inv1  gate1800(.a(G27), .O(gate67inter7));
  inv1  gate1801(.a(G305), .O(gate67inter8));
  nand2 gate1802(.a(gate67inter8), .b(gate67inter7), .O(gate67inter9));
  nand2 gate1803(.a(s_179), .b(gate67inter3), .O(gate67inter10));
  nor2  gate1804(.a(gate67inter10), .b(gate67inter9), .O(gate67inter11));
  nor2  gate1805(.a(gate67inter11), .b(gate67inter6), .O(gate67inter12));
  nand2 gate1806(.a(gate67inter12), .b(gate67inter1), .O(G388));
nand2 gate68( .a(G28), .b(G305), .O(G389) );

  xor2  gate1373(.a(G308), .b(G29), .O(gate69inter0));
  nand2 gate1374(.a(gate69inter0), .b(s_118), .O(gate69inter1));
  and2  gate1375(.a(G308), .b(G29), .O(gate69inter2));
  inv1  gate1376(.a(s_118), .O(gate69inter3));
  inv1  gate1377(.a(s_119), .O(gate69inter4));
  nand2 gate1378(.a(gate69inter4), .b(gate69inter3), .O(gate69inter5));
  nor2  gate1379(.a(gate69inter5), .b(gate69inter2), .O(gate69inter6));
  inv1  gate1380(.a(G29), .O(gate69inter7));
  inv1  gate1381(.a(G308), .O(gate69inter8));
  nand2 gate1382(.a(gate69inter8), .b(gate69inter7), .O(gate69inter9));
  nand2 gate1383(.a(s_119), .b(gate69inter3), .O(gate69inter10));
  nor2  gate1384(.a(gate69inter10), .b(gate69inter9), .O(gate69inter11));
  nor2  gate1385(.a(gate69inter11), .b(gate69inter6), .O(gate69inter12));
  nand2 gate1386(.a(gate69inter12), .b(gate69inter1), .O(G390));
nand2 gate70( .a(G30), .b(G308), .O(G391) );

  xor2  gate757(.a(G311), .b(G31), .O(gate71inter0));
  nand2 gate758(.a(gate71inter0), .b(s_30), .O(gate71inter1));
  and2  gate759(.a(G311), .b(G31), .O(gate71inter2));
  inv1  gate760(.a(s_30), .O(gate71inter3));
  inv1  gate761(.a(s_31), .O(gate71inter4));
  nand2 gate762(.a(gate71inter4), .b(gate71inter3), .O(gate71inter5));
  nor2  gate763(.a(gate71inter5), .b(gate71inter2), .O(gate71inter6));
  inv1  gate764(.a(G31), .O(gate71inter7));
  inv1  gate765(.a(G311), .O(gate71inter8));
  nand2 gate766(.a(gate71inter8), .b(gate71inter7), .O(gate71inter9));
  nand2 gate767(.a(s_31), .b(gate71inter3), .O(gate71inter10));
  nor2  gate768(.a(gate71inter10), .b(gate71inter9), .O(gate71inter11));
  nor2  gate769(.a(gate71inter11), .b(gate71inter6), .O(gate71inter12));
  nand2 gate770(.a(gate71inter12), .b(gate71inter1), .O(G392));

  xor2  gate1331(.a(G311), .b(G32), .O(gate72inter0));
  nand2 gate1332(.a(gate72inter0), .b(s_112), .O(gate72inter1));
  and2  gate1333(.a(G311), .b(G32), .O(gate72inter2));
  inv1  gate1334(.a(s_112), .O(gate72inter3));
  inv1  gate1335(.a(s_113), .O(gate72inter4));
  nand2 gate1336(.a(gate72inter4), .b(gate72inter3), .O(gate72inter5));
  nor2  gate1337(.a(gate72inter5), .b(gate72inter2), .O(gate72inter6));
  inv1  gate1338(.a(G32), .O(gate72inter7));
  inv1  gate1339(.a(G311), .O(gate72inter8));
  nand2 gate1340(.a(gate72inter8), .b(gate72inter7), .O(gate72inter9));
  nand2 gate1341(.a(s_113), .b(gate72inter3), .O(gate72inter10));
  nor2  gate1342(.a(gate72inter10), .b(gate72inter9), .O(gate72inter11));
  nor2  gate1343(.a(gate72inter11), .b(gate72inter6), .O(gate72inter12));
  nand2 gate1344(.a(gate72inter12), .b(gate72inter1), .O(G393));

  xor2  gate1401(.a(G314), .b(G1), .O(gate73inter0));
  nand2 gate1402(.a(gate73inter0), .b(s_122), .O(gate73inter1));
  and2  gate1403(.a(G314), .b(G1), .O(gate73inter2));
  inv1  gate1404(.a(s_122), .O(gate73inter3));
  inv1  gate1405(.a(s_123), .O(gate73inter4));
  nand2 gate1406(.a(gate73inter4), .b(gate73inter3), .O(gate73inter5));
  nor2  gate1407(.a(gate73inter5), .b(gate73inter2), .O(gate73inter6));
  inv1  gate1408(.a(G1), .O(gate73inter7));
  inv1  gate1409(.a(G314), .O(gate73inter8));
  nand2 gate1410(.a(gate73inter8), .b(gate73inter7), .O(gate73inter9));
  nand2 gate1411(.a(s_123), .b(gate73inter3), .O(gate73inter10));
  nor2  gate1412(.a(gate73inter10), .b(gate73inter9), .O(gate73inter11));
  nor2  gate1413(.a(gate73inter11), .b(gate73inter6), .O(gate73inter12));
  nand2 gate1414(.a(gate73inter12), .b(gate73inter1), .O(G394));
nand2 gate74( .a(G5), .b(G314), .O(G395) );
nand2 gate75( .a(G9), .b(G317), .O(G396) );

  xor2  gate1527(.a(G317), .b(G13), .O(gate76inter0));
  nand2 gate1528(.a(gate76inter0), .b(s_140), .O(gate76inter1));
  and2  gate1529(.a(G317), .b(G13), .O(gate76inter2));
  inv1  gate1530(.a(s_140), .O(gate76inter3));
  inv1  gate1531(.a(s_141), .O(gate76inter4));
  nand2 gate1532(.a(gate76inter4), .b(gate76inter3), .O(gate76inter5));
  nor2  gate1533(.a(gate76inter5), .b(gate76inter2), .O(gate76inter6));
  inv1  gate1534(.a(G13), .O(gate76inter7));
  inv1  gate1535(.a(G317), .O(gate76inter8));
  nand2 gate1536(.a(gate76inter8), .b(gate76inter7), .O(gate76inter9));
  nand2 gate1537(.a(s_141), .b(gate76inter3), .O(gate76inter10));
  nor2  gate1538(.a(gate76inter10), .b(gate76inter9), .O(gate76inter11));
  nor2  gate1539(.a(gate76inter11), .b(gate76inter6), .O(gate76inter12));
  nand2 gate1540(.a(gate76inter12), .b(gate76inter1), .O(G397));
nand2 gate77( .a(G2), .b(G320), .O(G398) );
nand2 gate78( .a(G6), .b(G320), .O(G399) );
nand2 gate79( .a(G10), .b(G323), .O(G400) );
nand2 gate80( .a(G14), .b(G323), .O(G401) );
nand2 gate81( .a(G3), .b(G326), .O(G402) );
nand2 gate82( .a(G7), .b(G326), .O(G403) );

  xor2  gate673(.a(G329), .b(G11), .O(gate83inter0));
  nand2 gate674(.a(gate83inter0), .b(s_18), .O(gate83inter1));
  and2  gate675(.a(G329), .b(G11), .O(gate83inter2));
  inv1  gate676(.a(s_18), .O(gate83inter3));
  inv1  gate677(.a(s_19), .O(gate83inter4));
  nand2 gate678(.a(gate83inter4), .b(gate83inter3), .O(gate83inter5));
  nor2  gate679(.a(gate83inter5), .b(gate83inter2), .O(gate83inter6));
  inv1  gate680(.a(G11), .O(gate83inter7));
  inv1  gate681(.a(G329), .O(gate83inter8));
  nand2 gate682(.a(gate83inter8), .b(gate83inter7), .O(gate83inter9));
  nand2 gate683(.a(s_19), .b(gate83inter3), .O(gate83inter10));
  nor2  gate684(.a(gate83inter10), .b(gate83inter9), .O(gate83inter11));
  nor2  gate685(.a(gate83inter11), .b(gate83inter6), .O(gate83inter12));
  nand2 gate686(.a(gate83inter12), .b(gate83inter1), .O(G404));
nand2 gate84( .a(G15), .b(G329), .O(G405) );

  xor2  gate2143(.a(G332), .b(G4), .O(gate85inter0));
  nand2 gate2144(.a(gate85inter0), .b(s_228), .O(gate85inter1));
  and2  gate2145(.a(G332), .b(G4), .O(gate85inter2));
  inv1  gate2146(.a(s_228), .O(gate85inter3));
  inv1  gate2147(.a(s_229), .O(gate85inter4));
  nand2 gate2148(.a(gate85inter4), .b(gate85inter3), .O(gate85inter5));
  nor2  gate2149(.a(gate85inter5), .b(gate85inter2), .O(gate85inter6));
  inv1  gate2150(.a(G4), .O(gate85inter7));
  inv1  gate2151(.a(G332), .O(gate85inter8));
  nand2 gate2152(.a(gate85inter8), .b(gate85inter7), .O(gate85inter9));
  nand2 gate2153(.a(s_229), .b(gate85inter3), .O(gate85inter10));
  nor2  gate2154(.a(gate85inter10), .b(gate85inter9), .O(gate85inter11));
  nor2  gate2155(.a(gate85inter11), .b(gate85inter6), .O(gate85inter12));
  nand2 gate2156(.a(gate85inter12), .b(gate85inter1), .O(G406));

  xor2  gate617(.a(G332), .b(G8), .O(gate86inter0));
  nand2 gate618(.a(gate86inter0), .b(s_10), .O(gate86inter1));
  and2  gate619(.a(G332), .b(G8), .O(gate86inter2));
  inv1  gate620(.a(s_10), .O(gate86inter3));
  inv1  gate621(.a(s_11), .O(gate86inter4));
  nand2 gate622(.a(gate86inter4), .b(gate86inter3), .O(gate86inter5));
  nor2  gate623(.a(gate86inter5), .b(gate86inter2), .O(gate86inter6));
  inv1  gate624(.a(G8), .O(gate86inter7));
  inv1  gate625(.a(G332), .O(gate86inter8));
  nand2 gate626(.a(gate86inter8), .b(gate86inter7), .O(gate86inter9));
  nand2 gate627(.a(s_11), .b(gate86inter3), .O(gate86inter10));
  nor2  gate628(.a(gate86inter10), .b(gate86inter9), .O(gate86inter11));
  nor2  gate629(.a(gate86inter11), .b(gate86inter6), .O(gate86inter12));
  nand2 gate630(.a(gate86inter12), .b(gate86inter1), .O(G407));

  xor2  gate1667(.a(G335), .b(G12), .O(gate87inter0));
  nand2 gate1668(.a(gate87inter0), .b(s_160), .O(gate87inter1));
  and2  gate1669(.a(G335), .b(G12), .O(gate87inter2));
  inv1  gate1670(.a(s_160), .O(gate87inter3));
  inv1  gate1671(.a(s_161), .O(gate87inter4));
  nand2 gate1672(.a(gate87inter4), .b(gate87inter3), .O(gate87inter5));
  nor2  gate1673(.a(gate87inter5), .b(gate87inter2), .O(gate87inter6));
  inv1  gate1674(.a(G12), .O(gate87inter7));
  inv1  gate1675(.a(G335), .O(gate87inter8));
  nand2 gate1676(.a(gate87inter8), .b(gate87inter7), .O(gate87inter9));
  nand2 gate1677(.a(s_161), .b(gate87inter3), .O(gate87inter10));
  nor2  gate1678(.a(gate87inter10), .b(gate87inter9), .O(gate87inter11));
  nor2  gate1679(.a(gate87inter11), .b(gate87inter6), .O(gate87inter12));
  nand2 gate1680(.a(gate87inter12), .b(gate87inter1), .O(G408));
nand2 gate88( .a(G16), .b(G335), .O(G409) );
nand2 gate89( .a(G17), .b(G338), .O(G410) );
nand2 gate90( .a(G21), .b(G338), .O(G411) );

  xor2  gate1513(.a(G341), .b(G25), .O(gate91inter0));
  nand2 gate1514(.a(gate91inter0), .b(s_138), .O(gate91inter1));
  and2  gate1515(.a(G341), .b(G25), .O(gate91inter2));
  inv1  gate1516(.a(s_138), .O(gate91inter3));
  inv1  gate1517(.a(s_139), .O(gate91inter4));
  nand2 gate1518(.a(gate91inter4), .b(gate91inter3), .O(gate91inter5));
  nor2  gate1519(.a(gate91inter5), .b(gate91inter2), .O(gate91inter6));
  inv1  gate1520(.a(G25), .O(gate91inter7));
  inv1  gate1521(.a(G341), .O(gate91inter8));
  nand2 gate1522(.a(gate91inter8), .b(gate91inter7), .O(gate91inter9));
  nand2 gate1523(.a(s_139), .b(gate91inter3), .O(gate91inter10));
  nor2  gate1524(.a(gate91inter10), .b(gate91inter9), .O(gate91inter11));
  nor2  gate1525(.a(gate91inter11), .b(gate91inter6), .O(gate91inter12));
  nand2 gate1526(.a(gate91inter12), .b(gate91inter1), .O(G412));

  xor2  gate2283(.a(G341), .b(G29), .O(gate92inter0));
  nand2 gate2284(.a(gate92inter0), .b(s_248), .O(gate92inter1));
  and2  gate2285(.a(G341), .b(G29), .O(gate92inter2));
  inv1  gate2286(.a(s_248), .O(gate92inter3));
  inv1  gate2287(.a(s_249), .O(gate92inter4));
  nand2 gate2288(.a(gate92inter4), .b(gate92inter3), .O(gate92inter5));
  nor2  gate2289(.a(gate92inter5), .b(gate92inter2), .O(gate92inter6));
  inv1  gate2290(.a(G29), .O(gate92inter7));
  inv1  gate2291(.a(G341), .O(gate92inter8));
  nand2 gate2292(.a(gate92inter8), .b(gate92inter7), .O(gate92inter9));
  nand2 gate2293(.a(s_249), .b(gate92inter3), .O(gate92inter10));
  nor2  gate2294(.a(gate92inter10), .b(gate92inter9), .O(gate92inter11));
  nor2  gate2295(.a(gate92inter11), .b(gate92inter6), .O(gate92inter12));
  nand2 gate2296(.a(gate92inter12), .b(gate92inter1), .O(G413));
nand2 gate93( .a(G18), .b(G344), .O(G414) );
nand2 gate94( .a(G22), .b(G344), .O(G415) );
nand2 gate95( .a(G26), .b(G347), .O(G416) );
nand2 gate96( .a(G30), .b(G347), .O(G417) );
nand2 gate97( .a(G19), .b(G350), .O(G418) );
nand2 gate98( .a(G23), .b(G350), .O(G419) );
nand2 gate99( .a(G27), .b(G353), .O(G420) );
nand2 gate100( .a(G31), .b(G353), .O(G421) );
nand2 gate101( .a(G20), .b(G356), .O(G422) );
nand2 gate102( .a(G24), .b(G356), .O(G423) );
nand2 gate103( .a(G28), .b(G359), .O(G424) );
nand2 gate104( .a(G32), .b(G359), .O(G425) );

  xor2  gate687(.a(G363), .b(G362), .O(gate105inter0));
  nand2 gate688(.a(gate105inter0), .b(s_20), .O(gate105inter1));
  and2  gate689(.a(G363), .b(G362), .O(gate105inter2));
  inv1  gate690(.a(s_20), .O(gate105inter3));
  inv1  gate691(.a(s_21), .O(gate105inter4));
  nand2 gate692(.a(gate105inter4), .b(gate105inter3), .O(gate105inter5));
  nor2  gate693(.a(gate105inter5), .b(gate105inter2), .O(gate105inter6));
  inv1  gate694(.a(G362), .O(gate105inter7));
  inv1  gate695(.a(G363), .O(gate105inter8));
  nand2 gate696(.a(gate105inter8), .b(gate105inter7), .O(gate105inter9));
  nand2 gate697(.a(s_21), .b(gate105inter3), .O(gate105inter10));
  nor2  gate698(.a(gate105inter10), .b(gate105inter9), .O(gate105inter11));
  nor2  gate699(.a(gate105inter11), .b(gate105inter6), .O(gate105inter12));
  nand2 gate700(.a(gate105inter12), .b(gate105inter1), .O(G426));

  xor2  gate855(.a(G365), .b(G364), .O(gate106inter0));
  nand2 gate856(.a(gate106inter0), .b(s_44), .O(gate106inter1));
  and2  gate857(.a(G365), .b(G364), .O(gate106inter2));
  inv1  gate858(.a(s_44), .O(gate106inter3));
  inv1  gate859(.a(s_45), .O(gate106inter4));
  nand2 gate860(.a(gate106inter4), .b(gate106inter3), .O(gate106inter5));
  nor2  gate861(.a(gate106inter5), .b(gate106inter2), .O(gate106inter6));
  inv1  gate862(.a(G364), .O(gate106inter7));
  inv1  gate863(.a(G365), .O(gate106inter8));
  nand2 gate864(.a(gate106inter8), .b(gate106inter7), .O(gate106inter9));
  nand2 gate865(.a(s_45), .b(gate106inter3), .O(gate106inter10));
  nor2  gate866(.a(gate106inter10), .b(gate106inter9), .O(gate106inter11));
  nor2  gate867(.a(gate106inter11), .b(gate106inter6), .O(gate106inter12));
  nand2 gate868(.a(gate106inter12), .b(gate106inter1), .O(G429));

  xor2  gate1961(.a(G367), .b(G366), .O(gate107inter0));
  nand2 gate1962(.a(gate107inter0), .b(s_202), .O(gate107inter1));
  and2  gate1963(.a(G367), .b(G366), .O(gate107inter2));
  inv1  gate1964(.a(s_202), .O(gate107inter3));
  inv1  gate1965(.a(s_203), .O(gate107inter4));
  nand2 gate1966(.a(gate107inter4), .b(gate107inter3), .O(gate107inter5));
  nor2  gate1967(.a(gate107inter5), .b(gate107inter2), .O(gate107inter6));
  inv1  gate1968(.a(G366), .O(gate107inter7));
  inv1  gate1969(.a(G367), .O(gate107inter8));
  nand2 gate1970(.a(gate107inter8), .b(gate107inter7), .O(gate107inter9));
  nand2 gate1971(.a(s_203), .b(gate107inter3), .O(gate107inter10));
  nor2  gate1972(.a(gate107inter10), .b(gate107inter9), .O(gate107inter11));
  nor2  gate1973(.a(gate107inter11), .b(gate107inter6), .O(gate107inter12));
  nand2 gate1974(.a(gate107inter12), .b(gate107inter1), .O(G432));
nand2 gate108( .a(G368), .b(G369), .O(G435) );
nand2 gate109( .a(G370), .b(G371), .O(G438) );
nand2 gate110( .a(G372), .b(G373), .O(G441) );
nand2 gate111( .a(G374), .b(G375), .O(G444) );
nand2 gate112( .a(G376), .b(G377), .O(G447) );
nand2 gate113( .a(G378), .b(G379), .O(G450) );
nand2 gate114( .a(G380), .b(G381), .O(G453) );
nand2 gate115( .a(G382), .b(G383), .O(G456) );

  xor2  gate561(.a(G385), .b(G384), .O(gate116inter0));
  nand2 gate562(.a(gate116inter0), .b(s_2), .O(gate116inter1));
  and2  gate563(.a(G385), .b(G384), .O(gate116inter2));
  inv1  gate564(.a(s_2), .O(gate116inter3));
  inv1  gate565(.a(s_3), .O(gate116inter4));
  nand2 gate566(.a(gate116inter4), .b(gate116inter3), .O(gate116inter5));
  nor2  gate567(.a(gate116inter5), .b(gate116inter2), .O(gate116inter6));
  inv1  gate568(.a(G384), .O(gate116inter7));
  inv1  gate569(.a(G385), .O(gate116inter8));
  nand2 gate570(.a(gate116inter8), .b(gate116inter7), .O(gate116inter9));
  nand2 gate571(.a(s_3), .b(gate116inter3), .O(gate116inter10));
  nor2  gate572(.a(gate116inter10), .b(gate116inter9), .O(gate116inter11));
  nor2  gate573(.a(gate116inter11), .b(gate116inter6), .O(gate116inter12));
  nand2 gate574(.a(gate116inter12), .b(gate116inter1), .O(G459));
nand2 gate117( .a(G386), .b(G387), .O(G462) );
nand2 gate118( .a(G388), .b(G389), .O(G465) );
nand2 gate119( .a(G390), .b(G391), .O(G468) );
nand2 gate120( .a(G392), .b(G393), .O(G471) );
nand2 gate121( .a(G394), .b(G395), .O(G474) );
nand2 gate122( .a(G396), .b(G397), .O(G477) );
nand2 gate123( .a(G398), .b(G399), .O(G480) );
nand2 gate124( .a(G400), .b(G401), .O(G483) );
nand2 gate125( .a(G402), .b(G403), .O(G486) );
nand2 gate126( .a(G404), .b(G405), .O(G489) );

  xor2  gate2157(.a(G407), .b(G406), .O(gate127inter0));
  nand2 gate2158(.a(gate127inter0), .b(s_230), .O(gate127inter1));
  and2  gate2159(.a(G407), .b(G406), .O(gate127inter2));
  inv1  gate2160(.a(s_230), .O(gate127inter3));
  inv1  gate2161(.a(s_231), .O(gate127inter4));
  nand2 gate2162(.a(gate127inter4), .b(gate127inter3), .O(gate127inter5));
  nor2  gate2163(.a(gate127inter5), .b(gate127inter2), .O(gate127inter6));
  inv1  gate2164(.a(G406), .O(gate127inter7));
  inv1  gate2165(.a(G407), .O(gate127inter8));
  nand2 gate2166(.a(gate127inter8), .b(gate127inter7), .O(gate127inter9));
  nand2 gate2167(.a(s_231), .b(gate127inter3), .O(gate127inter10));
  nor2  gate2168(.a(gate127inter10), .b(gate127inter9), .O(gate127inter11));
  nor2  gate2169(.a(gate127inter11), .b(gate127inter6), .O(gate127inter12));
  nand2 gate2170(.a(gate127inter12), .b(gate127inter1), .O(G492));
nand2 gate128( .a(G408), .b(G409), .O(G495) );
nand2 gate129( .a(G410), .b(G411), .O(G498) );
nand2 gate130( .a(G412), .b(G413), .O(G501) );
nand2 gate131( .a(G414), .b(G415), .O(G504) );
nand2 gate132( .a(G416), .b(G417), .O(G507) );
nand2 gate133( .a(G418), .b(G419), .O(G510) );
nand2 gate134( .a(G420), .b(G421), .O(G513) );
nand2 gate135( .a(G422), .b(G423), .O(G516) );

  xor2  gate925(.a(G425), .b(G424), .O(gate136inter0));
  nand2 gate926(.a(gate136inter0), .b(s_54), .O(gate136inter1));
  and2  gate927(.a(G425), .b(G424), .O(gate136inter2));
  inv1  gate928(.a(s_54), .O(gate136inter3));
  inv1  gate929(.a(s_55), .O(gate136inter4));
  nand2 gate930(.a(gate136inter4), .b(gate136inter3), .O(gate136inter5));
  nor2  gate931(.a(gate136inter5), .b(gate136inter2), .O(gate136inter6));
  inv1  gate932(.a(G424), .O(gate136inter7));
  inv1  gate933(.a(G425), .O(gate136inter8));
  nand2 gate934(.a(gate136inter8), .b(gate136inter7), .O(gate136inter9));
  nand2 gate935(.a(s_55), .b(gate136inter3), .O(gate136inter10));
  nor2  gate936(.a(gate136inter10), .b(gate136inter9), .O(gate136inter11));
  nor2  gate937(.a(gate136inter11), .b(gate136inter6), .O(gate136inter12));
  nand2 gate938(.a(gate136inter12), .b(gate136inter1), .O(G519));

  xor2  gate1723(.a(G429), .b(G426), .O(gate137inter0));
  nand2 gate1724(.a(gate137inter0), .b(s_168), .O(gate137inter1));
  and2  gate1725(.a(G429), .b(G426), .O(gate137inter2));
  inv1  gate1726(.a(s_168), .O(gate137inter3));
  inv1  gate1727(.a(s_169), .O(gate137inter4));
  nand2 gate1728(.a(gate137inter4), .b(gate137inter3), .O(gate137inter5));
  nor2  gate1729(.a(gate137inter5), .b(gate137inter2), .O(gate137inter6));
  inv1  gate1730(.a(G426), .O(gate137inter7));
  inv1  gate1731(.a(G429), .O(gate137inter8));
  nand2 gate1732(.a(gate137inter8), .b(gate137inter7), .O(gate137inter9));
  nand2 gate1733(.a(s_169), .b(gate137inter3), .O(gate137inter10));
  nor2  gate1734(.a(gate137inter10), .b(gate137inter9), .O(gate137inter11));
  nor2  gate1735(.a(gate137inter11), .b(gate137inter6), .O(gate137inter12));
  nand2 gate1736(.a(gate137inter12), .b(gate137inter1), .O(G522));

  xor2  gate1863(.a(G435), .b(G432), .O(gate138inter0));
  nand2 gate1864(.a(gate138inter0), .b(s_188), .O(gate138inter1));
  and2  gate1865(.a(G435), .b(G432), .O(gate138inter2));
  inv1  gate1866(.a(s_188), .O(gate138inter3));
  inv1  gate1867(.a(s_189), .O(gate138inter4));
  nand2 gate1868(.a(gate138inter4), .b(gate138inter3), .O(gate138inter5));
  nor2  gate1869(.a(gate138inter5), .b(gate138inter2), .O(gate138inter6));
  inv1  gate1870(.a(G432), .O(gate138inter7));
  inv1  gate1871(.a(G435), .O(gate138inter8));
  nand2 gate1872(.a(gate138inter8), .b(gate138inter7), .O(gate138inter9));
  nand2 gate1873(.a(s_189), .b(gate138inter3), .O(gate138inter10));
  nor2  gate1874(.a(gate138inter10), .b(gate138inter9), .O(gate138inter11));
  nor2  gate1875(.a(gate138inter11), .b(gate138inter6), .O(gate138inter12));
  nand2 gate1876(.a(gate138inter12), .b(gate138inter1), .O(G525));
nand2 gate139( .a(G438), .b(G441), .O(G528) );

  xor2  gate2213(.a(G447), .b(G444), .O(gate140inter0));
  nand2 gate2214(.a(gate140inter0), .b(s_238), .O(gate140inter1));
  and2  gate2215(.a(G447), .b(G444), .O(gate140inter2));
  inv1  gate2216(.a(s_238), .O(gate140inter3));
  inv1  gate2217(.a(s_239), .O(gate140inter4));
  nand2 gate2218(.a(gate140inter4), .b(gate140inter3), .O(gate140inter5));
  nor2  gate2219(.a(gate140inter5), .b(gate140inter2), .O(gate140inter6));
  inv1  gate2220(.a(G444), .O(gate140inter7));
  inv1  gate2221(.a(G447), .O(gate140inter8));
  nand2 gate2222(.a(gate140inter8), .b(gate140inter7), .O(gate140inter9));
  nand2 gate2223(.a(s_239), .b(gate140inter3), .O(gate140inter10));
  nor2  gate2224(.a(gate140inter10), .b(gate140inter9), .O(gate140inter11));
  nor2  gate2225(.a(gate140inter11), .b(gate140inter6), .O(gate140inter12));
  nand2 gate2226(.a(gate140inter12), .b(gate140inter1), .O(G531));
nand2 gate141( .a(G450), .b(G453), .O(G534) );

  xor2  gate1289(.a(G459), .b(G456), .O(gate142inter0));
  nand2 gate1290(.a(gate142inter0), .b(s_106), .O(gate142inter1));
  and2  gate1291(.a(G459), .b(G456), .O(gate142inter2));
  inv1  gate1292(.a(s_106), .O(gate142inter3));
  inv1  gate1293(.a(s_107), .O(gate142inter4));
  nand2 gate1294(.a(gate142inter4), .b(gate142inter3), .O(gate142inter5));
  nor2  gate1295(.a(gate142inter5), .b(gate142inter2), .O(gate142inter6));
  inv1  gate1296(.a(G456), .O(gate142inter7));
  inv1  gate1297(.a(G459), .O(gate142inter8));
  nand2 gate1298(.a(gate142inter8), .b(gate142inter7), .O(gate142inter9));
  nand2 gate1299(.a(s_107), .b(gate142inter3), .O(gate142inter10));
  nor2  gate1300(.a(gate142inter10), .b(gate142inter9), .O(gate142inter11));
  nor2  gate1301(.a(gate142inter11), .b(gate142inter6), .O(gate142inter12));
  nand2 gate1302(.a(gate142inter12), .b(gate142inter1), .O(G537));
nand2 gate143( .a(G462), .b(G465), .O(G540) );

  xor2  gate1471(.a(G471), .b(G468), .O(gate144inter0));
  nand2 gate1472(.a(gate144inter0), .b(s_132), .O(gate144inter1));
  and2  gate1473(.a(G471), .b(G468), .O(gate144inter2));
  inv1  gate1474(.a(s_132), .O(gate144inter3));
  inv1  gate1475(.a(s_133), .O(gate144inter4));
  nand2 gate1476(.a(gate144inter4), .b(gate144inter3), .O(gate144inter5));
  nor2  gate1477(.a(gate144inter5), .b(gate144inter2), .O(gate144inter6));
  inv1  gate1478(.a(G468), .O(gate144inter7));
  inv1  gate1479(.a(G471), .O(gate144inter8));
  nand2 gate1480(.a(gate144inter8), .b(gate144inter7), .O(gate144inter9));
  nand2 gate1481(.a(s_133), .b(gate144inter3), .O(gate144inter10));
  nor2  gate1482(.a(gate144inter10), .b(gate144inter9), .O(gate144inter11));
  nor2  gate1483(.a(gate144inter11), .b(gate144inter6), .O(gate144inter12));
  nand2 gate1484(.a(gate144inter12), .b(gate144inter1), .O(G543));
nand2 gate145( .a(G474), .b(G477), .O(G546) );
nand2 gate146( .a(G480), .b(G483), .O(G549) );
nand2 gate147( .a(G486), .b(G489), .O(G552) );
nand2 gate148( .a(G492), .b(G495), .O(G555) );
nand2 gate149( .a(G498), .b(G501), .O(G558) );

  xor2  gate1653(.a(G507), .b(G504), .O(gate150inter0));
  nand2 gate1654(.a(gate150inter0), .b(s_158), .O(gate150inter1));
  and2  gate1655(.a(G507), .b(G504), .O(gate150inter2));
  inv1  gate1656(.a(s_158), .O(gate150inter3));
  inv1  gate1657(.a(s_159), .O(gate150inter4));
  nand2 gate1658(.a(gate150inter4), .b(gate150inter3), .O(gate150inter5));
  nor2  gate1659(.a(gate150inter5), .b(gate150inter2), .O(gate150inter6));
  inv1  gate1660(.a(G504), .O(gate150inter7));
  inv1  gate1661(.a(G507), .O(gate150inter8));
  nand2 gate1662(.a(gate150inter8), .b(gate150inter7), .O(gate150inter9));
  nand2 gate1663(.a(s_159), .b(gate150inter3), .O(gate150inter10));
  nor2  gate1664(.a(gate150inter10), .b(gate150inter9), .O(gate150inter11));
  nor2  gate1665(.a(gate150inter11), .b(gate150inter6), .O(gate150inter12));
  nand2 gate1666(.a(gate150inter12), .b(gate150inter1), .O(G561));
nand2 gate151( .a(G510), .b(G513), .O(G564) );
nand2 gate152( .a(G516), .b(G519), .O(G567) );
nand2 gate153( .a(G426), .b(G522), .O(G570) );
nand2 gate154( .a(G429), .b(G522), .O(G571) );
nand2 gate155( .a(G432), .b(G525), .O(G572) );
nand2 gate156( .a(G435), .b(G525), .O(G573) );
nand2 gate157( .a(G438), .b(G528), .O(G574) );
nand2 gate158( .a(G441), .b(G528), .O(G575) );

  xor2  gate603(.a(G531), .b(G444), .O(gate159inter0));
  nand2 gate604(.a(gate159inter0), .b(s_8), .O(gate159inter1));
  and2  gate605(.a(G531), .b(G444), .O(gate159inter2));
  inv1  gate606(.a(s_8), .O(gate159inter3));
  inv1  gate607(.a(s_9), .O(gate159inter4));
  nand2 gate608(.a(gate159inter4), .b(gate159inter3), .O(gate159inter5));
  nor2  gate609(.a(gate159inter5), .b(gate159inter2), .O(gate159inter6));
  inv1  gate610(.a(G444), .O(gate159inter7));
  inv1  gate611(.a(G531), .O(gate159inter8));
  nand2 gate612(.a(gate159inter8), .b(gate159inter7), .O(gate159inter9));
  nand2 gate613(.a(s_9), .b(gate159inter3), .O(gate159inter10));
  nor2  gate614(.a(gate159inter10), .b(gate159inter9), .O(gate159inter11));
  nor2  gate615(.a(gate159inter11), .b(gate159inter6), .O(gate159inter12));
  nand2 gate616(.a(gate159inter12), .b(gate159inter1), .O(G576));
nand2 gate160( .a(G447), .b(G531), .O(G577) );
nand2 gate161( .a(G450), .b(G534), .O(G578) );
nand2 gate162( .a(G453), .b(G534), .O(G579) );
nand2 gate163( .a(G456), .b(G537), .O(G580) );

  xor2  gate2017(.a(G537), .b(G459), .O(gate164inter0));
  nand2 gate2018(.a(gate164inter0), .b(s_210), .O(gate164inter1));
  and2  gate2019(.a(G537), .b(G459), .O(gate164inter2));
  inv1  gate2020(.a(s_210), .O(gate164inter3));
  inv1  gate2021(.a(s_211), .O(gate164inter4));
  nand2 gate2022(.a(gate164inter4), .b(gate164inter3), .O(gate164inter5));
  nor2  gate2023(.a(gate164inter5), .b(gate164inter2), .O(gate164inter6));
  inv1  gate2024(.a(G459), .O(gate164inter7));
  inv1  gate2025(.a(G537), .O(gate164inter8));
  nand2 gate2026(.a(gate164inter8), .b(gate164inter7), .O(gate164inter9));
  nand2 gate2027(.a(s_211), .b(gate164inter3), .O(gate164inter10));
  nor2  gate2028(.a(gate164inter10), .b(gate164inter9), .O(gate164inter11));
  nor2  gate2029(.a(gate164inter11), .b(gate164inter6), .O(gate164inter12));
  nand2 gate2030(.a(gate164inter12), .b(gate164inter1), .O(G581));
nand2 gate165( .a(G462), .b(G540), .O(G582) );

  xor2  gate953(.a(G540), .b(G465), .O(gate166inter0));
  nand2 gate954(.a(gate166inter0), .b(s_58), .O(gate166inter1));
  and2  gate955(.a(G540), .b(G465), .O(gate166inter2));
  inv1  gate956(.a(s_58), .O(gate166inter3));
  inv1  gate957(.a(s_59), .O(gate166inter4));
  nand2 gate958(.a(gate166inter4), .b(gate166inter3), .O(gate166inter5));
  nor2  gate959(.a(gate166inter5), .b(gate166inter2), .O(gate166inter6));
  inv1  gate960(.a(G465), .O(gate166inter7));
  inv1  gate961(.a(G540), .O(gate166inter8));
  nand2 gate962(.a(gate166inter8), .b(gate166inter7), .O(gate166inter9));
  nand2 gate963(.a(s_59), .b(gate166inter3), .O(gate166inter10));
  nor2  gate964(.a(gate166inter10), .b(gate166inter9), .O(gate166inter11));
  nor2  gate965(.a(gate166inter11), .b(gate166inter6), .O(gate166inter12));
  nand2 gate966(.a(gate166inter12), .b(gate166inter1), .O(G583));
nand2 gate167( .a(G468), .b(G543), .O(G584) );
nand2 gate168( .a(G471), .b(G543), .O(G585) );
nand2 gate169( .a(G474), .b(G546), .O(G586) );
nand2 gate170( .a(G477), .b(G546), .O(G587) );
nand2 gate171( .a(G480), .b(G549), .O(G588) );
nand2 gate172( .a(G483), .b(G549), .O(G589) );

  xor2  gate1275(.a(G552), .b(G486), .O(gate173inter0));
  nand2 gate1276(.a(gate173inter0), .b(s_104), .O(gate173inter1));
  and2  gate1277(.a(G552), .b(G486), .O(gate173inter2));
  inv1  gate1278(.a(s_104), .O(gate173inter3));
  inv1  gate1279(.a(s_105), .O(gate173inter4));
  nand2 gate1280(.a(gate173inter4), .b(gate173inter3), .O(gate173inter5));
  nor2  gate1281(.a(gate173inter5), .b(gate173inter2), .O(gate173inter6));
  inv1  gate1282(.a(G486), .O(gate173inter7));
  inv1  gate1283(.a(G552), .O(gate173inter8));
  nand2 gate1284(.a(gate173inter8), .b(gate173inter7), .O(gate173inter9));
  nand2 gate1285(.a(s_105), .b(gate173inter3), .O(gate173inter10));
  nor2  gate1286(.a(gate173inter10), .b(gate173inter9), .O(gate173inter11));
  nor2  gate1287(.a(gate173inter11), .b(gate173inter6), .O(gate173inter12));
  nand2 gate1288(.a(gate173inter12), .b(gate173inter1), .O(G590));
nand2 gate174( .a(G489), .b(G552), .O(G591) );
nand2 gate175( .a(G492), .b(G555), .O(G592) );
nand2 gate176( .a(G495), .b(G555), .O(G593) );
nand2 gate177( .a(G498), .b(G558), .O(G594) );

  xor2  gate1835(.a(G558), .b(G501), .O(gate178inter0));
  nand2 gate1836(.a(gate178inter0), .b(s_184), .O(gate178inter1));
  and2  gate1837(.a(G558), .b(G501), .O(gate178inter2));
  inv1  gate1838(.a(s_184), .O(gate178inter3));
  inv1  gate1839(.a(s_185), .O(gate178inter4));
  nand2 gate1840(.a(gate178inter4), .b(gate178inter3), .O(gate178inter5));
  nor2  gate1841(.a(gate178inter5), .b(gate178inter2), .O(gate178inter6));
  inv1  gate1842(.a(G501), .O(gate178inter7));
  inv1  gate1843(.a(G558), .O(gate178inter8));
  nand2 gate1844(.a(gate178inter8), .b(gate178inter7), .O(gate178inter9));
  nand2 gate1845(.a(s_185), .b(gate178inter3), .O(gate178inter10));
  nor2  gate1846(.a(gate178inter10), .b(gate178inter9), .O(gate178inter11));
  nor2  gate1847(.a(gate178inter11), .b(gate178inter6), .O(gate178inter12));
  nand2 gate1848(.a(gate178inter12), .b(gate178inter1), .O(G595));

  xor2  gate981(.a(G561), .b(G504), .O(gate179inter0));
  nand2 gate982(.a(gate179inter0), .b(s_62), .O(gate179inter1));
  and2  gate983(.a(G561), .b(G504), .O(gate179inter2));
  inv1  gate984(.a(s_62), .O(gate179inter3));
  inv1  gate985(.a(s_63), .O(gate179inter4));
  nand2 gate986(.a(gate179inter4), .b(gate179inter3), .O(gate179inter5));
  nor2  gate987(.a(gate179inter5), .b(gate179inter2), .O(gate179inter6));
  inv1  gate988(.a(G504), .O(gate179inter7));
  inv1  gate989(.a(G561), .O(gate179inter8));
  nand2 gate990(.a(gate179inter8), .b(gate179inter7), .O(gate179inter9));
  nand2 gate991(.a(s_63), .b(gate179inter3), .O(gate179inter10));
  nor2  gate992(.a(gate179inter10), .b(gate179inter9), .O(gate179inter11));
  nor2  gate993(.a(gate179inter11), .b(gate179inter6), .O(gate179inter12));
  nand2 gate994(.a(gate179inter12), .b(gate179inter1), .O(G596));
nand2 gate180( .a(G507), .b(G561), .O(G597) );
nand2 gate181( .a(G510), .b(G564), .O(G598) );
nand2 gate182( .a(G513), .b(G564), .O(G599) );

  xor2  gate2101(.a(G567), .b(G516), .O(gate183inter0));
  nand2 gate2102(.a(gate183inter0), .b(s_222), .O(gate183inter1));
  and2  gate2103(.a(G567), .b(G516), .O(gate183inter2));
  inv1  gate2104(.a(s_222), .O(gate183inter3));
  inv1  gate2105(.a(s_223), .O(gate183inter4));
  nand2 gate2106(.a(gate183inter4), .b(gate183inter3), .O(gate183inter5));
  nor2  gate2107(.a(gate183inter5), .b(gate183inter2), .O(gate183inter6));
  inv1  gate2108(.a(G516), .O(gate183inter7));
  inv1  gate2109(.a(G567), .O(gate183inter8));
  nand2 gate2110(.a(gate183inter8), .b(gate183inter7), .O(gate183inter9));
  nand2 gate2111(.a(s_223), .b(gate183inter3), .O(gate183inter10));
  nor2  gate2112(.a(gate183inter10), .b(gate183inter9), .O(gate183inter11));
  nor2  gate2113(.a(gate183inter11), .b(gate183inter6), .O(gate183inter12));
  nand2 gate2114(.a(gate183inter12), .b(gate183inter1), .O(G600));
nand2 gate184( .a(G519), .b(G567), .O(G601) );
nand2 gate185( .a(G570), .b(G571), .O(G602) );
nand2 gate186( .a(G572), .b(G573), .O(G607) );
nand2 gate187( .a(G574), .b(G575), .O(G612) );
nand2 gate188( .a(G576), .b(G577), .O(G617) );
nand2 gate189( .a(G578), .b(G579), .O(G622) );
nand2 gate190( .a(G580), .b(G581), .O(G627) );
nand2 gate191( .a(G582), .b(G583), .O(G632) );
nand2 gate192( .a(G584), .b(G585), .O(G637) );

  xor2  gate2241(.a(G587), .b(G586), .O(gate193inter0));
  nand2 gate2242(.a(gate193inter0), .b(s_242), .O(gate193inter1));
  and2  gate2243(.a(G587), .b(G586), .O(gate193inter2));
  inv1  gate2244(.a(s_242), .O(gate193inter3));
  inv1  gate2245(.a(s_243), .O(gate193inter4));
  nand2 gate2246(.a(gate193inter4), .b(gate193inter3), .O(gate193inter5));
  nor2  gate2247(.a(gate193inter5), .b(gate193inter2), .O(gate193inter6));
  inv1  gate2248(.a(G586), .O(gate193inter7));
  inv1  gate2249(.a(G587), .O(gate193inter8));
  nand2 gate2250(.a(gate193inter8), .b(gate193inter7), .O(gate193inter9));
  nand2 gate2251(.a(s_243), .b(gate193inter3), .O(gate193inter10));
  nor2  gate2252(.a(gate193inter10), .b(gate193inter9), .O(gate193inter11));
  nor2  gate2253(.a(gate193inter11), .b(gate193inter6), .O(gate193inter12));
  nand2 gate2254(.a(gate193inter12), .b(gate193inter1), .O(G642));
nand2 gate194( .a(G588), .b(G589), .O(G645) );

  xor2  gate1597(.a(G591), .b(G590), .O(gate195inter0));
  nand2 gate1598(.a(gate195inter0), .b(s_150), .O(gate195inter1));
  and2  gate1599(.a(G591), .b(G590), .O(gate195inter2));
  inv1  gate1600(.a(s_150), .O(gate195inter3));
  inv1  gate1601(.a(s_151), .O(gate195inter4));
  nand2 gate1602(.a(gate195inter4), .b(gate195inter3), .O(gate195inter5));
  nor2  gate1603(.a(gate195inter5), .b(gate195inter2), .O(gate195inter6));
  inv1  gate1604(.a(G590), .O(gate195inter7));
  inv1  gate1605(.a(G591), .O(gate195inter8));
  nand2 gate1606(.a(gate195inter8), .b(gate195inter7), .O(gate195inter9));
  nand2 gate1607(.a(s_151), .b(gate195inter3), .O(gate195inter10));
  nor2  gate1608(.a(gate195inter10), .b(gate195inter9), .O(gate195inter11));
  nor2  gate1609(.a(gate195inter11), .b(gate195inter6), .O(gate195inter12));
  nand2 gate1610(.a(gate195inter12), .b(gate195inter1), .O(G648));
nand2 gate196( .a(G592), .b(G593), .O(G651) );
nand2 gate197( .a(G594), .b(G595), .O(G654) );

  xor2  gate1779(.a(G597), .b(G596), .O(gate198inter0));
  nand2 gate1780(.a(gate198inter0), .b(s_176), .O(gate198inter1));
  and2  gate1781(.a(G597), .b(G596), .O(gate198inter2));
  inv1  gate1782(.a(s_176), .O(gate198inter3));
  inv1  gate1783(.a(s_177), .O(gate198inter4));
  nand2 gate1784(.a(gate198inter4), .b(gate198inter3), .O(gate198inter5));
  nor2  gate1785(.a(gate198inter5), .b(gate198inter2), .O(gate198inter6));
  inv1  gate1786(.a(G596), .O(gate198inter7));
  inv1  gate1787(.a(G597), .O(gate198inter8));
  nand2 gate1788(.a(gate198inter8), .b(gate198inter7), .O(gate198inter9));
  nand2 gate1789(.a(s_177), .b(gate198inter3), .O(gate198inter10));
  nor2  gate1790(.a(gate198inter10), .b(gate198inter9), .O(gate198inter11));
  nor2  gate1791(.a(gate198inter11), .b(gate198inter6), .O(gate198inter12));
  nand2 gate1792(.a(gate198inter12), .b(gate198inter1), .O(G657));

  xor2  gate2227(.a(G599), .b(G598), .O(gate199inter0));
  nand2 gate2228(.a(gate199inter0), .b(s_240), .O(gate199inter1));
  and2  gate2229(.a(G599), .b(G598), .O(gate199inter2));
  inv1  gate2230(.a(s_240), .O(gate199inter3));
  inv1  gate2231(.a(s_241), .O(gate199inter4));
  nand2 gate2232(.a(gate199inter4), .b(gate199inter3), .O(gate199inter5));
  nor2  gate2233(.a(gate199inter5), .b(gate199inter2), .O(gate199inter6));
  inv1  gate2234(.a(G598), .O(gate199inter7));
  inv1  gate2235(.a(G599), .O(gate199inter8));
  nand2 gate2236(.a(gate199inter8), .b(gate199inter7), .O(gate199inter9));
  nand2 gate2237(.a(s_241), .b(gate199inter3), .O(gate199inter10));
  nor2  gate2238(.a(gate199inter10), .b(gate199inter9), .O(gate199inter11));
  nor2  gate2239(.a(gate199inter11), .b(gate199inter6), .O(gate199inter12));
  nand2 gate2240(.a(gate199inter12), .b(gate199inter1), .O(G660));

  xor2  gate631(.a(G601), .b(G600), .O(gate200inter0));
  nand2 gate632(.a(gate200inter0), .b(s_12), .O(gate200inter1));
  and2  gate633(.a(G601), .b(G600), .O(gate200inter2));
  inv1  gate634(.a(s_12), .O(gate200inter3));
  inv1  gate635(.a(s_13), .O(gate200inter4));
  nand2 gate636(.a(gate200inter4), .b(gate200inter3), .O(gate200inter5));
  nor2  gate637(.a(gate200inter5), .b(gate200inter2), .O(gate200inter6));
  inv1  gate638(.a(G600), .O(gate200inter7));
  inv1  gate639(.a(G601), .O(gate200inter8));
  nand2 gate640(.a(gate200inter8), .b(gate200inter7), .O(gate200inter9));
  nand2 gate641(.a(s_13), .b(gate200inter3), .O(gate200inter10));
  nor2  gate642(.a(gate200inter10), .b(gate200inter9), .O(gate200inter11));
  nor2  gate643(.a(gate200inter11), .b(gate200inter6), .O(gate200inter12));
  nand2 gate644(.a(gate200inter12), .b(gate200inter1), .O(G663));
nand2 gate201( .a(G602), .b(G607), .O(G666) );

  xor2  gate827(.a(G617), .b(G612), .O(gate202inter0));
  nand2 gate828(.a(gate202inter0), .b(s_40), .O(gate202inter1));
  and2  gate829(.a(G617), .b(G612), .O(gate202inter2));
  inv1  gate830(.a(s_40), .O(gate202inter3));
  inv1  gate831(.a(s_41), .O(gate202inter4));
  nand2 gate832(.a(gate202inter4), .b(gate202inter3), .O(gate202inter5));
  nor2  gate833(.a(gate202inter5), .b(gate202inter2), .O(gate202inter6));
  inv1  gate834(.a(G612), .O(gate202inter7));
  inv1  gate835(.a(G617), .O(gate202inter8));
  nand2 gate836(.a(gate202inter8), .b(gate202inter7), .O(gate202inter9));
  nand2 gate837(.a(s_41), .b(gate202inter3), .O(gate202inter10));
  nor2  gate838(.a(gate202inter10), .b(gate202inter9), .O(gate202inter11));
  nor2  gate839(.a(gate202inter11), .b(gate202inter6), .O(gate202inter12));
  nand2 gate840(.a(gate202inter12), .b(gate202inter1), .O(G669));
nand2 gate203( .a(G602), .b(G612), .O(G672) );
nand2 gate204( .a(G607), .b(G617), .O(G675) );

  xor2  gate2297(.a(G627), .b(G622), .O(gate205inter0));
  nand2 gate2298(.a(gate205inter0), .b(s_250), .O(gate205inter1));
  and2  gate2299(.a(G627), .b(G622), .O(gate205inter2));
  inv1  gate2300(.a(s_250), .O(gate205inter3));
  inv1  gate2301(.a(s_251), .O(gate205inter4));
  nand2 gate2302(.a(gate205inter4), .b(gate205inter3), .O(gate205inter5));
  nor2  gate2303(.a(gate205inter5), .b(gate205inter2), .O(gate205inter6));
  inv1  gate2304(.a(G622), .O(gate205inter7));
  inv1  gate2305(.a(G627), .O(gate205inter8));
  nand2 gate2306(.a(gate205inter8), .b(gate205inter7), .O(gate205inter9));
  nand2 gate2307(.a(s_251), .b(gate205inter3), .O(gate205inter10));
  nor2  gate2308(.a(gate205inter10), .b(gate205inter9), .O(gate205inter11));
  nor2  gate2309(.a(gate205inter11), .b(gate205inter6), .O(gate205inter12));
  nand2 gate2310(.a(gate205inter12), .b(gate205inter1), .O(G678));

  xor2  gate1205(.a(G637), .b(G632), .O(gate206inter0));
  nand2 gate1206(.a(gate206inter0), .b(s_94), .O(gate206inter1));
  and2  gate1207(.a(G637), .b(G632), .O(gate206inter2));
  inv1  gate1208(.a(s_94), .O(gate206inter3));
  inv1  gate1209(.a(s_95), .O(gate206inter4));
  nand2 gate1210(.a(gate206inter4), .b(gate206inter3), .O(gate206inter5));
  nor2  gate1211(.a(gate206inter5), .b(gate206inter2), .O(gate206inter6));
  inv1  gate1212(.a(G632), .O(gate206inter7));
  inv1  gate1213(.a(G637), .O(gate206inter8));
  nand2 gate1214(.a(gate206inter8), .b(gate206inter7), .O(gate206inter9));
  nand2 gate1215(.a(s_95), .b(gate206inter3), .O(gate206inter10));
  nor2  gate1216(.a(gate206inter10), .b(gate206inter9), .O(gate206inter11));
  nor2  gate1217(.a(gate206inter11), .b(gate206inter6), .O(gate206inter12));
  nand2 gate1218(.a(gate206inter12), .b(gate206inter1), .O(G681));
nand2 gate207( .a(G622), .b(G632), .O(G684) );
nand2 gate208( .a(G627), .b(G637), .O(G687) );
nand2 gate209( .a(G602), .b(G666), .O(G690) );

  xor2  gate785(.a(G666), .b(G607), .O(gate210inter0));
  nand2 gate786(.a(gate210inter0), .b(s_34), .O(gate210inter1));
  and2  gate787(.a(G666), .b(G607), .O(gate210inter2));
  inv1  gate788(.a(s_34), .O(gate210inter3));
  inv1  gate789(.a(s_35), .O(gate210inter4));
  nand2 gate790(.a(gate210inter4), .b(gate210inter3), .O(gate210inter5));
  nor2  gate791(.a(gate210inter5), .b(gate210inter2), .O(gate210inter6));
  inv1  gate792(.a(G607), .O(gate210inter7));
  inv1  gate793(.a(G666), .O(gate210inter8));
  nand2 gate794(.a(gate210inter8), .b(gate210inter7), .O(gate210inter9));
  nand2 gate795(.a(s_35), .b(gate210inter3), .O(gate210inter10));
  nor2  gate796(.a(gate210inter10), .b(gate210inter9), .O(gate210inter11));
  nor2  gate797(.a(gate210inter11), .b(gate210inter6), .O(gate210inter12));
  nand2 gate798(.a(gate210inter12), .b(gate210inter1), .O(G691));
nand2 gate211( .a(G612), .b(G669), .O(G692) );
nand2 gate212( .a(G617), .b(G669), .O(G693) );
nand2 gate213( .a(G602), .b(G672), .O(G694) );
nand2 gate214( .a(G612), .b(G672), .O(G695) );
nand2 gate215( .a(G607), .b(G675), .O(G696) );
nand2 gate216( .a(G617), .b(G675), .O(G697) );
nand2 gate217( .a(G622), .b(G678), .O(G698) );
nand2 gate218( .a(G627), .b(G678), .O(G699) );
nand2 gate219( .a(G632), .b(G681), .O(G700) );

  xor2  gate1303(.a(G681), .b(G637), .O(gate220inter0));
  nand2 gate1304(.a(gate220inter0), .b(s_108), .O(gate220inter1));
  and2  gate1305(.a(G681), .b(G637), .O(gate220inter2));
  inv1  gate1306(.a(s_108), .O(gate220inter3));
  inv1  gate1307(.a(s_109), .O(gate220inter4));
  nand2 gate1308(.a(gate220inter4), .b(gate220inter3), .O(gate220inter5));
  nor2  gate1309(.a(gate220inter5), .b(gate220inter2), .O(gate220inter6));
  inv1  gate1310(.a(G637), .O(gate220inter7));
  inv1  gate1311(.a(G681), .O(gate220inter8));
  nand2 gate1312(.a(gate220inter8), .b(gate220inter7), .O(gate220inter9));
  nand2 gate1313(.a(s_109), .b(gate220inter3), .O(gate220inter10));
  nor2  gate1314(.a(gate220inter10), .b(gate220inter9), .O(gate220inter11));
  nor2  gate1315(.a(gate220inter11), .b(gate220inter6), .O(gate220inter12));
  nand2 gate1316(.a(gate220inter12), .b(gate220inter1), .O(G701));
nand2 gate221( .a(G622), .b(G684), .O(G702) );
nand2 gate222( .a(G632), .b(G684), .O(G703) );
nand2 gate223( .a(G627), .b(G687), .O(G704) );

  xor2  gate1163(.a(G687), .b(G637), .O(gate224inter0));
  nand2 gate1164(.a(gate224inter0), .b(s_88), .O(gate224inter1));
  and2  gate1165(.a(G687), .b(G637), .O(gate224inter2));
  inv1  gate1166(.a(s_88), .O(gate224inter3));
  inv1  gate1167(.a(s_89), .O(gate224inter4));
  nand2 gate1168(.a(gate224inter4), .b(gate224inter3), .O(gate224inter5));
  nor2  gate1169(.a(gate224inter5), .b(gate224inter2), .O(gate224inter6));
  inv1  gate1170(.a(G637), .O(gate224inter7));
  inv1  gate1171(.a(G687), .O(gate224inter8));
  nand2 gate1172(.a(gate224inter8), .b(gate224inter7), .O(gate224inter9));
  nand2 gate1173(.a(s_89), .b(gate224inter3), .O(gate224inter10));
  nor2  gate1174(.a(gate224inter10), .b(gate224inter9), .O(gate224inter11));
  nor2  gate1175(.a(gate224inter11), .b(gate224inter6), .O(gate224inter12));
  nand2 gate1176(.a(gate224inter12), .b(gate224inter1), .O(G705));
nand2 gate225( .a(G690), .b(G691), .O(G706) );
nand2 gate226( .a(G692), .b(G693), .O(G709) );

  xor2  gate1191(.a(G695), .b(G694), .O(gate227inter0));
  nand2 gate1192(.a(gate227inter0), .b(s_92), .O(gate227inter1));
  and2  gate1193(.a(G695), .b(G694), .O(gate227inter2));
  inv1  gate1194(.a(s_92), .O(gate227inter3));
  inv1  gate1195(.a(s_93), .O(gate227inter4));
  nand2 gate1196(.a(gate227inter4), .b(gate227inter3), .O(gate227inter5));
  nor2  gate1197(.a(gate227inter5), .b(gate227inter2), .O(gate227inter6));
  inv1  gate1198(.a(G694), .O(gate227inter7));
  inv1  gate1199(.a(G695), .O(gate227inter8));
  nand2 gate1200(.a(gate227inter8), .b(gate227inter7), .O(gate227inter9));
  nand2 gate1201(.a(s_93), .b(gate227inter3), .O(gate227inter10));
  nor2  gate1202(.a(gate227inter10), .b(gate227inter9), .O(gate227inter11));
  nor2  gate1203(.a(gate227inter11), .b(gate227inter6), .O(gate227inter12));
  nand2 gate1204(.a(gate227inter12), .b(gate227inter1), .O(G712));
nand2 gate228( .a(G696), .b(G697), .O(G715) );
nand2 gate229( .a(G698), .b(G699), .O(G718) );
nand2 gate230( .a(G700), .b(G701), .O(G721) );

  xor2  gate1121(.a(G703), .b(G702), .O(gate231inter0));
  nand2 gate1122(.a(gate231inter0), .b(s_82), .O(gate231inter1));
  and2  gate1123(.a(G703), .b(G702), .O(gate231inter2));
  inv1  gate1124(.a(s_82), .O(gate231inter3));
  inv1  gate1125(.a(s_83), .O(gate231inter4));
  nand2 gate1126(.a(gate231inter4), .b(gate231inter3), .O(gate231inter5));
  nor2  gate1127(.a(gate231inter5), .b(gate231inter2), .O(gate231inter6));
  inv1  gate1128(.a(G702), .O(gate231inter7));
  inv1  gate1129(.a(G703), .O(gate231inter8));
  nand2 gate1130(.a(gate231inter8), .b(gate231inter7), .O(gate231inter9));
  nand2 gate1131(.a(s_83), .b(gate231inter3), .O(gate231inter10));
  nor2  gate1132(.a(gate231inter10), .b(gate231inter9), .O(gate231inter11));
  nor2  gate1133(.a(gate231inter11), .b(gate231inter6), .O(gate231inter12));
  nand2 gate1134(.a(gate231inter12), .b(gate231inter1), .O(G724));

  xor2  gate1975(.a(G705), .b(G704), .O(gate232inter0));
  nand2 gate1976(.a(gate232inter0), .b(s_204), .O(gate232inter1));
  and2  gate1977(.a(G705), .b(G704), .O(gate232inter2));
  inv1  gate1978(.a(s_204), .O(gate232inter3));
  inv1  gate1979(.a(s_205), .O(gate232inter4));
  nand2 gate1980(.a(gate232inter4), .b(gate232inter3), .O(gate232inter5));
  nor2  gate1981(.a(gate232inter5), .b(gate232inter2), .O(gate232inter6));
  inv1  gate1982(.a(G704), .O(gate232inter7));
  inv1  gate1983(.a(G705), .O(gate232inter8));
  nand2 gate1984(.a(gate232inter8), .b(gate232inter7), .O(gate232inter9));
  nand2 gate1985(.a(s_205), .b(gate232inter3), .O(gate232inter10));
  nor2  gate1986(.a(gate232inter10), .b(gate232inter9), .O(gate232inter11));
  nor2  gate1987(.a(gate232inter11), .b(gate232inter6), .O(gate232inter12));
  nand2 gate1988(.a(gate232inter12), .b(gate232inter1), .O(G727));
nand2 gate233( .a(G242), .b(G718), .O(G730) );
nand2 gate234( .a(G245), .b(G721), .O(G733) );
nand2 gate235( .a(G248), .b(G724), .O(G736) );

  xor2  gate1611(.a(G727), .b(G251), .O(gate236inter0));
  nand2 gate1612(.a(gate236inter0), .b(s_152), .O(gate236inter1));
  and2  gate1613(.a(G727), .b(G251), .O(gate236inter2));
  inv1  gate1614(.a(s_152), .O(gate236inter3));
  inv1  gate1615(.a(s_153), .O(gate236inter4));
  nand2 gate1616(.a(gate236inter4), .b(gate236inter3), .O(gate236inter5));
  nor2  gate1617(.a(gate236inter5), .b(gate236inter2), .O(gate236inter6));
  inv1  gate1618(.a(G251), .O(gate236inter7));
  inv1  gate1619(.a(G727), .O(gate236inter8));
  nand2 gate1620(.a(gate236inter8), .b(gate236inter7), .O(gate236inter9));
  nand2 gate1621(.a(s_153), .b(gate236inter3), .O(gate236inter10));
  nor2  gate1622(.a(gate236inter10), .b(gate236inter9), .O(gate236inter11));
  nor2  gate1623(.a(gate236inter11), .b(gate236inter6), .O(gate236inter12));
  nand2 gate1624(.a(gate236inter12), .b(gate236inter1), .O(G739));

  xor2  gate743(.a(G706), .b(G254), .O(gate237inter0));
  nand2 gate744(.a(gate237inter0), .b(s_28), .O(gate237inter1));
  and2  gate745(.a(G706), .b(G254), .O(gate237inter2));
  inv1  gate746(.a(s_28), .O(gate237inter3));
  inv1  gate747(.a(s_29), .O(gate237inter4));
  nand2 gate748(.a(gate237inter4), .b(gate237inter3), .O(gate237inter5));
  nor2  gate749(.a(gate237inter5), .b(gate237inter2), .O(gate237inter6));
  inv1  gate750(.a(G254), .O(gate237inter7));
  inv1  gate751(.a(G706), .O(gate237inter8));
  nand2 gate752(.a(gate237inter8), .b(gate237inter7), .O(gate237inter9));
  nand2 gate753(.a(s_29), .b(gate237inter3), .O(gate237inter10));
  nor2  gate754(.a(gate237inter10), .b(gate237inter9), .O(gate237inter11));
  nor2  gate755(.a(gate237inter11), .b(gate237inter6), .O(gate237inter12));
  nand2 gate756(.a(gate237inter12), .b(gate237inter1), .O(G742));
nand2 gate238( .a(G257), .b(G709), .O(G745) );
nand2 gate239( .a(G260), .b(G712), .O(G748) );

  xor2  gate1359(.a(G715), .b(G263), .O(gate240inter0));
  nand2 gate1360(.a(gate240inter0), .b(s_116), .O(gate240inter1));
  and2  gate1361(.a(G715), .b(G263), .O(gate240inter2));
  inv1  gate1362(.a(s_116), .O(gate240inter3));
  inv1  gate1363(.a(s_117), .O(gate240inter4));
  nand2 gate1364(.a(gate240inter4), .b(gate240inter3), .O(gate240inter5));
  nor2  gate1365(.a(gate240inter5), .b(gate240inter2), .O(gate240inter6));
  inv1  gate1366(.a(G263), .O(gate240inter7));
  inv1  gate1367(.a(G715), .O(gate240inter8));
  nand2 gate1368(.a(gate240inter8), .b(gate240inter7), .O(gate240inter9));
  nand2 gate1369(.a(s_117), .b(gate240inter3), .O(gate240inter10));
  nor2  gate1370(.a(gate240inter10), .b(gate240inter9), .O(gate240inter11));
  nor2  gate1371(.a(gate240inter11), .b(gate240inter6), .O(gate240inter12));
  nand2 gate1372(.a(gate240inter12), .b(gate240inter1), .O(G751));
nand2 gate241( .a(G242), .b(G730), .O(G754) );

  xor2  gate1919(.a(G730), .b(G718), .O(gate242inter0));
  nand2 gate1920(.a(gate242inter0), .b(s_196), .O(gate242inter1));
  and2  gate1921(.a(G730), .b(G718), .O(gate242inter2));
  inv1  gate1922(.a(s_196), .O(gate242inter3));
  inv1  gate1923(.a(s_197), .O(gate242inter4));
  nand2 gate1924(.a(gate242inter4), .b(gate242inter3), .O(gate242inter5));
  nor2  gate1925(.a(gate242inter5), .b(gate242inter2), .O(gate242inter6));
  inv1  gate1926(.a(G718), .O(gate242inter7));
  inv1  gate1927(.a(G730), .O(gate242inter8));
  nand2 gate1928(.a(gate242inter8), .b(gate242inter7), .O(gate242inter9));
  nand2 gate1929(.a(s_197), .b(gate242inter3), .O(gate242inter10));
  nor2  gate1930(.a(gate242inter10), .b(gate242inter9), .O(gate242inter11));
  nor2  gate1931(.a(gate242inter11), .b(gate242inter6), .O(gate242inter12));
  nand2 gate1932(.a(gate242inter12), .b(gate242inter1), .O(G755));

  xor2  gate1583(.a(G733), .b(G245), .O(gate243inter0));
  nand2 gate1584(.a(gate243inter0), .b(s_148), .O(gate243inter1));
  and2  gate1585(.a(G733), .b(G245), .O(gate243inter2));
  inv1  gate1586(.a(s_148), .O(gate243inter3));
  inv1  gate1587(.a(s_149), .O(gate243inter4));
  nand2 gate1588(.a(gate243inter4), .b(gate243inter3), .O(gate243inter5));
  nor2  gate1589(.a(gate243inter5), .b(gate243inter2), .O(gate243inter6));
  inv1  gate1590(.a(G245), .O(gate243inter7));
  inv1  gate1591(.a(G733), .O(gate243inter8));
  nand2 gate1592(.a(gate243inter8), .b(gate243inter7), .O(gate243inter9));
  nand2 gate1593(.a(s_149), .b(gate243inter3), .O(gate243inter10));
  nor2  gate1594(.a(gate243inter10), .b(gate243inter9), .O(gate243inter11));
  nor2  gate1595(.a(gate243inter11), .b(gate243inter6), .O(gate243inter12));
  nand2 gate1596(.a(gate243inter12), .b(gate243inter1), .O(G756));
nand2 gate244( .a(G721), .b(G733), .O(G757) );
nand2 gate245( .a(G248), .b(G736), .O(G758) );
nand2 gate246( .a(G724), .b(G736), .O(G759) );

  xor2  gate1751(.a(G739), .b(G251), .O(gate247inter0));
  nand2 gate1752(.a(gate247inter0), .b(s_172), .O(gate247inter1));
  and2  gate1753(.a(G739), .b(G251), .O(gate247inter2));
  inv1  gate1754(.a(s_172), .O(gate247inter3));
  inv1  gate1755(.a(s_173), .O(gate247inter4));
  nand2 gate1756(.a(gate247inter4), .b(gate247inter3), .O(gate247inter5));
  nor2  gate1757(.a(gate247inter5), .b(gate247inter2), .O(gate247inter6));
  inv1  gate1758(.a(G251), .O(gate247inter7));
  inv1  gate1759(.a(G739), .O(gate247inter8));
  nand2 gate1760(.a(gate247inter8), .b(gate247inter7), .O(gate247inter9));
  nand2 gate1761(.a(s_173), .b(gate247inter3), .O(gate247inter10));
  nor2  gate1762(.a(gate247inter10), .b(gate247inter9), .O(gate247inter11));
  nor2  gate1763(.a(gate247inter11), .b(gate247inter6), .O(gate247inter12));
  nand2 gate1764(.a(gate247inter12), .b(gate247inter1), .O(G760));
nand2 gate248( .a(G727), .b(G739), .O(G761) );
nand2 gate249( .a(G254), .b(G742), .O(G762) );
nand2 gate250( .a(G706), .b(G742), .O(G763) );
nand2 gate251( .a(G257), .b(G745), .O(G764) );

  xor2  gate1765(.a(G745), .b(G709), .O(gate252inter0));
  nand2 gate1766(.a(gate252inter0), .b(s_174), .O(gate252inter1));
  and2  gate1767(.a(G745), .b(G709), .O(gate252inter2));
  inv1  gate1768(.a(s_174), .O(gate252inter3));
  inv1  gate1769(.a(s_175), .O(gate252inter4));
  nand2 gate1770(.a(gate252inter4), .b(gate252inter3), .O(gate252inter5));
  nor2  gate1771(.a(gate252inter5), .b(gate252inter2), .O(gate252inter6));
  inv1  gate1772(.a(G709), .O(gate252inter7));
  inv1  gate1773(.a(G745), .O(gate252inter8));
  nand2 gate1774(.a(gate252inter8), .b(gate252inter7), .O(gate252inter9));
  nand2 gate1775(.a(s_175), .b(gate252inter3), .O(gate252inter10));
  nor2  gate1776(.a(gate252inter10), .b(gate252inter9), .O(gate252inter11));
  nor2  gate1777(.a(gate252inter11), .b(gate252inter6), .O(gate252inter12));
  nand2 gate1778(.a(gate252inter12), .b(gate252inter1), .O(G765));
nand2 gate253( .a(G260), .b(G748), .O(G766) );
nand2 gate254( .a(G712), .b(G748), .O(G767) );
nand2 gate255( .a(G263), .b(G751), .O(G768) );
nand2 gate256( .a(G715), .b(G751), .O(G769) );
nand2 gate257( .a(G754), .b(G755), .O(G770) );
nand2 gate258( .a(G756), .b(G757), .O(G773) );
nand2 gate259( .a(G758), .b(G759), .O(G776) );

  xor2  gate1037(.a(G761), .b(G760), .O(gate260inter0));
  nand2 gate1038(.a(gate260inter0), .b(s_70), .O(gate260inter1));
  and2  gate1039(.a(G761), .b(G760), .O(gate260inter2));
  inv1  gate1040(.a(s_70), .O(gate260inter3));
  inv1  gate1041(.a(s_71), .O(gate260inter4));
  nand2 gate1042(.a(gate260inter4), .b(gate260inter3), .O(gate260inter5));
  nor2  gate1043(.a(gate260inter5), .b(gate260inter2), .O(gate260inter6));
  inv1  gate1044(.a(G760), .O(gate260inter7));
  inv1  gate1045(.a(G761), .O(gate260inter8));
  nand2 gate1046(.a(gate260inter8), .b(gate260inter7), .O(gate260inter9));
  nand2 gate1047(.a(s_71), .b(gate260inter3), .O(gate260inter10));
  nor2  gate1048(.a(gate260inter10), .b(gate260inter9), .O(gate260inter11));
  nor2  gate1049(.a(gate260inter11), .b(gate260inter6), .O(gate260inter12));
  nand2 gate1050(.a(gate260inter12), .b(gate260inter1), .O(G779));

  xor2  gate1821(.a(G763), .b(G762), .O(gate261inter0));
  nand2 gate1822(.a(gate261inter0), .b(s_182), .O(gate261inter1));
  and2  gate1823(.a(G763), .b(G762), .O(gate261inter2));
  inv1  gate1824(.a(s_182), .O(gate261inter3));
  inv1  gate1825(.a(s_183), .O(gate261inter4));
  nand2 gate1826(.a(gate261inter4), .b(gate261inter3), .O(gate261inter5));
  nor2  gate1827(.a(gate261inter5), .b(gate261inter2), .O(gate261inter6));
  inv1  gate1828(.a(G762), .O(gate261inter7));
  inv1  gate1829(.a(G763), .O(gate261inter8));
  nand2 gate1830(.a(gate261inter8), .b(gate261inter7), .O(gate261inter9));
  nand2 gate1831(.a(s_183), .b(gate261inter3), .O(gate261inter10));
  nor2  gate1832(.a(gate261inter10), .b(gate261inter9), .O(gate261inter11));
  nor2  gate1833(.a(gate261inter11), .b(gate261inter6), .O(gate261inter12));
  nand2 gate1834(.a(gate261inter12), .b(gate261inter1), .O(G782));
nand2 gate262( .a(G764), .b(G765), .O(G785) );
nand2 gate263( .a(G766), .b(G767), .O(G788) );
nand2 gate264( .a(G768), .b(G769), .O(G791) );
nand2 gate265( .a(G642), .b(G770), .O(G794) );
nand2 gate266( .a(G645), .b(G773), .O(G797) );
nand2 gate267( .a(G648), .b(G776), .O(G800) );

  xor2  gate1079(.a(G779), .b(G651), .O(gate268inter0));
  nand2 gate1080(.a(gate268inter0), .b(s_76), .O(gate268inter1));
  and2  gate1081(.a(G779), .b(G651), .O(gate268inter2));
  inv1  gate1082(.a(s_76), .O(gate268inter3));
  inv1  gate1083(.a(s_77), .O(gate268inter4));
  nand2 gate1084(.a(gate268inter4), .b(gate268inter3), .O(gate268inter5));
  nor2  gate1085(.a(gate268inter5), .b(gate268inter2), .O(gate268inter6));
  inv1  gate1086(.a(G651), .O(gate268inter7));
  inv1  gate1087(.a(G779), .O(gate268inter8));
  nand2 gate1088(.a(gate268inter8), .b(gate268inter7), .O(gate268inter9));
  nand2 gate1089(.a(s_77), .b(gate268inter3), .O(gate268inter10));
  nor2  gate1090(.a(gate268inter10), .b(gate268inter9), .O(gate268inter11));
  nor2  gate1091(.a(gate268inter11), .b(gate268inter6), .O(gate268inter12));
  nand2 gate1092(.a(gate268inter12), .b(gate268inter1), .O(G803));
nand2 gate269( .a(G654), .b(G782), .O(G806) );
nand2 gate270( .a(G657), .b(G785), .O(G809) );
nand2 gate271( .a(G660), .b(G788), .O(G812) );

  xor2  gate1317(.a(G791), .b(G663), .O(gate272inter0));
  nand2 gate1318(.a(gate272inter0), .b(s_110), .O(gate272inter1));
  and2  gate1319(.a(G791), .b(G663), .O(gate272inter2));
  inv1  gate1320(.a(s_110), .O(gate272inter3));
  inv1  gate1321(.a(s_111), .O(gate272inter4));
  nand2 gate1322(.a(gate272inter4), .b(gate272inter3), .O(gate272inter5));
  nor2  gate1323(.a(gate272inter5), .b(gate272inter2), .O(gate272inter6));
  inv1  gate1324(.a(G663), .O(gate272inter7));
  inv1  gate1325(.a(G791), .O(gate272inter8));
  nand2 gate1326(.a(gate272inter8), .b(gate272inter7), .O(gate272inter9));
  nand2 gate1327(.a(s_111), .b(gate272inter3), .O(gate272inter10));
  nor2  gate1328(.a(gate272inter10), .b(gate272inter9), .O(gate272inter11));
  nor2  gate1329(.a(gate272inter11), .b(gate272inter6), .O(gate272inter12));
  nand2 gate1330(.a(gate272inter12), .b(gate272inter1), .O(G815));

  xor2  gate869(.a(G794), .b(G642), .O(gate273inter0));
  nand2 gate870(.a(gate273inter0), .b(s_46), .O(gate273inter1));
  and2  gate871(.a(G794), .b(G642), .O(gate273inter2));
  inv1  gate872(.a(s_46), .O(gate273inter3));
  inv1  gate873(.a(s_47), .O(gate273inter4));
  nand2 gate874(.a(gate273inter4), .b(gate273inter3), .O(gate273inter5));
  nor2  gate875(.a(gate273inter5), .b(gate273inter2), .O(gate273inter6));
  inv1  gate876(.a(G642), .O(gate273inter7));
  inv1  gate877(.a(G794), .O(gate273inter8));
  nand2 gate878(.a(gate273inter8), .b(gate273inter7), .O(gate273inter9));
  nand2 gate879(.a(s_47), .b(gate273inter3), .O(gate273inter10));
  nor2  gate880(.a(gate273inter10), .b(gate273inter9), .O(gate273inter11));
  nor2  gate881(.a(gate273inter11), .b(gate273inter6), .O(gate273inter12));
  nand2 gate882(.a(gate273inter12), .b(gate273inter1), .O(G818));

  xor2  gate2045(.a(G794), .b(G770), .O(gate274inter0));
  nand2 gate2046(.a(gate274inter0), .b(s_214), .O(gate274inter1));
  and2  gate2047(.a(G794), .b(G770), .O(gate274inter2));
  inv1  gate2048(.a(s_214), .O(gate274inter3));
  inv1  gate2049(.a(s_215), .O(gate274inter4));
  nand2 gate2050(.a(gate274inter4), .b(gate274inter3), .O(gate274inter5));
  nor2  gate2051(.a(gate274inter5), .b(gate274inter2), .O(gate274inter6));
  inv1  gate2052(.a(G770), .O(gate274inter7));
  inv1  gate2053(.a(G794), .O(gate274inter8));
  nand2 gate2054(.a(gate274inter8), .b(gate274inter7), .O(gate274inter9));
  nand2 gate2055(.a(s_215), .b(gate274inter3), .O(gate274inter10));
  nor2  gate2056(.a(gate274inter10), .b(gate274inter9), .O(gate274inter11));
  nor2  gate2057(.a(gate274inter11), .b(gate274inter6), .O(gate274inter12));
  nand2 gate2058(.a(gate274inter12), .b(gate274inter1), .O(G819));

  xor2  gate967(.a(G797), .b(G645), .O(gate275inter0));
  nand2 gate968(.a(gate275inter0), .b(s_60), .O(gate275inter1));
  and2  gate969(.a(G797), .b(G645), .O(gate275inter2));
  inv1  gate970(.a(s_60), .O(gate275inter3));
  inv1  gate971(.a(s_61), .O(gate275inter4));
  nand2 gate972(.a(gate275inter4), .b(gate275inter3), .O(gate275inter5));
  nor2  gate973(.a(gate275inter5), .b(gate275inter2), .O(gate275inter6));
  inv1  gate974(.a(G645), .O(gate275inter7));
  inv1  gate975(.a(G797), .O(gate275inter8));
  nand2 gate976(.a(gate275inter8), .b(gate275inter7), .O(gate275inter9));
  nand2 gate977(.a(s_61), .b(gate275inter3), .O(gate275inter10));
  nor2  gate978(.a(gate275inter10), .b(gate275inter9), .O(gate275inter11));
  nor2  gate979(.a(gate275inter11), .b(gate275inter6), .O(gate275inter12));
  nand2 gate980(.a(gate275inter12), .b(gate275inter1), .O(G820));

  xor2  gate1345(.a(G797), .b(G773), .O(gate276inter0));
  nand2 gate1346(.a(gate276inter0), .b(s_114), .O(gate276inter1));
  and2  gate1347(.a(G797), .b(G773), .O(gate276inter2));
  inv1  gate1348(.a(s_114), .O(gate276inter3));
  inv1  gate1349(.a(s_115), .O(gate276inter4));
  nand2 gate1350(.a(gate276inter4), .b(gate276inter3), .O(gate276inter5));
  nor2  gate1351(.a(gate276inter5), .b(gate276inter2), .O(gate276inter6));
  inv1  gate1352(.a(G773), .O(gate276inter7));
  inv1  gate1353(.a(G797), .O(gate276inter8));
  nand2 gate1354(.a(gate276inter8), .b(gate276inter7), .O(gate276inter9));
  nand2 gate1355(.a(s_115), .b(gate276inter3), .O(gate276inter10));
  nor2  gate1356(.a(gate276inter10), .b(gate276inter9), .O(gate276inter11));
  nor2  gate1357(.a(gate276inter11), .b(gate276inter6), .O(gate276inter12));
  nand2 gate1358(.a(gate276inter12), .b(gate276inter1), .O(G821));
nand2 gate277( .a(G648), .b(G800), .O(G822) );
nand2 gate278( .a(G776), .b(G800), .O(G823) );

  xor2  gate1947(.a(G803), .b(G651), .O(gate279inter0));
  nand2 gate1948(.a(gate279inter0), .b(s_200), .O(gate279inter1));
  and2  gate1949(.a(G803), .b(G651), .O(gate279inter2));
  inv1  gate1950(.a(s_200), .O(gate279inter3));
  inv1  gate1951(.a(s_201), .O(gate279inter4));
  nand2 gate1952(.a(gate279inter4), .b(gate279inter3), .O(gate279inter5));
  nor2  gate1953(.a(gate279inter5), .b(gate279inter2), .O(gate279inter6));
  inv1  gate1954(.a(G651), .O(gate279inter7));
  inv1  gate1955(.a(G803), .O(gate279inter8));
  nand2 gate1956(.a(gate279inter8), .b(gate279inter7), .O(gate279inter9));
  nand2 gate1957(.a(s_201), .b(gate279inter3), .O(gate279inter10));
  nor2  gate1958(.a(gate279inter10), .b(gate279inter9), .O(gate279inter11));
  nor2  gate1959(.a(gate279inter11), .b(gate279inter6), .O(gate279inter12));
  nand2 gate1960(.a(gate279inter12), .b(gate279inter1), .O(G824));

  xor2  gate2199(.a(G803), .b(G779), .O(gate280inter0));
  nand2 gate2200(.a(gate280inter0), .b(s_236), .O(gate280inter1));
  and2  gate2201(.a(G803), .b(G779), .O(gate280inter2));
  inv1  gate2202(.a(s_236), .O(gate280inter3));
  inv1  gate2203(.a(s_237), .O(gate280inter4));
  nand2 gate2204(.a(gate280inter4), .b(gate280inter3), .O(gate280inter5));
  nor2  gate2205(.a(gate280inter5), .b(gate280inter2), .O(gate280inter6));
  inv1  gate2206(.a(G779), .O(gate280inter7));
  inv1  gate2207(.a(G803), .O(gate280inter8));
  nand2 gate2208(.a(gate280inter8), .b(gate280inter7), .O(gate280inter9));
  nand2 gate2209(.a(s_237), .b(gate280inter3), .O(gate280inter10));
  nor2  gate2210(.a(gate280inter10), .b(gate280inter9), .O(gate280inter11));
  nor2  gate2211(.a(gate280inter11), .b(gate280inter6), .O(gate280inter12));
  nand2 gate2212(.a(gate280inter12), .b(gate280inter1), .O(G825));

  xor2  gate995(.a(G806), .b(G654), .O(gate281inter0));
  nand2 gate996(.a(gate281inter0), .b(s_64), .O(gate281inter1));
  and2  gate997(.a(G806), .b(G654), .O(gate281inter2));
  inv1  gate998(.a(s_64), .O(gate281inter3));
  inv1  gate999(.a(s_65), .O(gate281inter4));
  nand2 gate1000(.a(gate281inter4), .b(gate281inter3), .O(gate281inter5));
  nor2  gate1001(.a(gate281inter5), .b(gate281inter2), .O(gate281inter6));
  inv1  gate1002(.a(G654), .O(gate281inter7));
  inv1  gate1003(.a(G806), .O(gate281inter8));
  nand2 gate1004(.a(gate281inter8), .b(gate281inter7), .O(gate281inter9));
  nand2 gate1005(.a(s_65), .b(gate281inter3), .O(gate281inter10));
  nor2  gate1006(.a(gate281inter10), .b(gate281inter9), .O(gate281inter11));
  nor2  gate1007(.a(gate281inter11), .b(gate281inter6), .O(gate281inter12));
  nand2 gate1008(.a(gate281inter12), .b(gate281inter1), .O(G826));

  xor2  gate1541(.a(G806), .b(G782), .O(gate282inter0));
  nand2 gate1542(.a(gate282inter0), .b(s_142), .O(gate282inter1));
  and2  gate1543(.a(G806), .b(G782), .O(gate282inter2));
  inv1  gate1544(.a(s_142), .O(gate282inter3));
  inv1  gate1545(.a(s_143), .O(gate282inter4));
  nand2 gate1546(.a(gate282inter4), .b(gate282inter3), .O(gate282inter5));
  nor2  gate1547(.a(gate282inter5), .b(gate282inter2), .O(gate282inter6));
  inv1  gate1548(.a(G782), .O(gate282inter7));
  inv1  gate1549(.a(G806), .O(gate282inter8));
  nand2 gate1550(.a(gate282inter8), .b(gate282inter7), .O(gate282inter9));
  nand2 gate1551(.a(s_143), .b(gate282inter3), .O(gate282inter10));
  nor2  gate1552(.a(gate282inter10), .b(gate282inter9), .O(gate282inter11));
  nor2  gate1553(.a(gate282inter11), .b(gate282inter6), .O(gate282inter12));
  nand2 gate1554(.a(gate282inter12), .b(gate282inter1), .O(G827));
nand2 gate283( .a(G657), .b(G809), .O(G828) );

  xor2  gate2003(.a(G809), .b(G785), .O(gate284inter0));
  nand2 gate2004(.a(gate284inter0), .b(s_208), .O(gate284inter1));
  and2  gate2005(.a(G809), .b(G785), .O(gate284inter2));
  inv1  gate2006(.a(s_208), .O(gate284inter3));
  inv1  gate2007(.a(s_209), .O(gate284inter4));
  nand2 gate2008(.a(gate284inter4), .b(gate284inter3), .O(gate284inter5));
  nor2  gate2009(.a(gate284inter5), .b(gate284inter2), .O(gate284inter6));
  inv1  gate2010(.a(G785), .O(gate284inter7));
  inv1  gate2011(.a(G809), .O(gate284inter8));
  nand2 gate2012(.a(gate284inter8), .b(gate284inter7), .O(gate284inter9));
  nand2 gate2013(.a(s_209), .b(gate284inter3), .O(gate284inter10));
  nor2  gate2014(.a(gate284inter10), .b(gate284inter9), .O(gate284inter11));
  nor2  gate2015(.a(gate284inter11), .b(gate284inter6), .O(gate284inter12));
  nand2 gate2016(.a(gate284inter12), .b(gate284inter1), .O(G829));
nand2 gate285( .a(G660), .b(G812), .O(G830) );
nand2 gate286( .a(G788), .b(G812), .O(G831) );

  xor2  gate771(.a(G815), .b(G663), .O(gate287inter0));
  nand2 gate772(.a(gate287inter0), .b(s_32), .O(gate287inter1));
  and2  gate773(.a(G815), .b(G663), .O(gate287inter2));
  inv1  gate774(.a(s_32), .O(gate287inter3));
  inv1  gate775(.a(s_33), .O(gate287inter4));
  nand2 gate776(.a(gate287inter4), .b(gate287inter3), .O(gate287inter5));
  nor2  gate777(.a(gate287inter5), .b(gate287inter2), .O(gate287inter6));
  inv1  gate778(.a(G663), .O(gate287inter7));
  inv1  gate779(.a(G815), .O(gate287inter8));
  nand2 gate780(.a(gate287inter8), .b(gate287inter7), .O(gate287inter9));
  nand2 gate781(.a(s_33), .b(gate287inter3), .O(gate287inter10));
  nor2  gate782(.a(gate287inter10), .b(gate287inter9), .O(gate287inter11));
  nor2  gate783(.a(gate287inter11), .b(gate287inter6), .O(gate287inter12));
  nand2 gate784(.a(gate287inter12), .b(gate287inter1), .O(G832));

  xor2  gate1247(.a(G815), .b(G791), .O(gate288inter0));
  nand2 gate1248(.a(gate288inter0), .b(s_100), .O(gate288inter1));
  and2  gate1249(.a(G815), .b(G791), .O(gate288inter2));
  inv1  gate1250(.a(s_100), .O(gate288inter3));
  inv1  gate1251(.a(s_101), .O(gate288inter4));
  nand2 gate1252(.a(gate288inter4), .b(gate288inter3), .O(gate288inter5));
  nor2  gate1253(.a(gate288inter5), .b(gate288inter2), .O(gate288inter6));
  inv1  gate1254(.a(G791), .O(gate288inter7));
  inv1  gate1255(.a(G815), .O(gate288inter8));
  nand2 gate1256(.a(gate288inter8), .b(gate288inter7), .O(gate288inter9));
  nand2 gate1257(.a(s_101), .b(gate288inter3), .O(gate288inter10));
  nor2  gate1258(.a(gate288inter10), .b(gate288inter9), .O(gate288inter11));
  nor2  gate1259(.a(gate288inter11), .b(gate288inter6), .O(gate288inter12));
  nand2 gate1260(.a(gate288inter12), .b(gate288inter1), .O(G833));
nand2 gate289( .a(G818), .b(G819), .O(G834) );
nand2 gate290( .a(G820), .b(G821), .O(G847) );

  xor2  gate1709(.a(G823), .b(G822), .O(gate291inter0));
  nand2 gate1710(.a(gate291inter0), .b(s_166), .O(gate291inter1));
  and2  gate1711(.a(G823), .b(G822), .O(gate291inter2));
  inv1  gate1712(.a(s_166), .O(gate291inter3));
  inv1  gate1713(.a(s_167), .O(gate291inter4));
  nand2 gate1714(.a(gate291inter4), .b(gate291inter3), .O(gate291inter5));
  nor2  gate1715(.a(gate291inter5), .b(gate291inter2), .O(gate291inter6));
  inv1  gate1716(.a(G822), .O(gate291inter7));
  inv1  gate1717(.a(G823), .O(gate291inter8));
  nand2 gate1718(.a(gate291inter8), .b(gate291inter7), .O(gate291inter9));
  nand2 gate1719(.a(s_167), .b(gate291inter3), .O(gate291inter10));
  nor2  gate1720(.a(gate291inter10), .b(gate291inter9), .O(gate291inter11));
  nor2  gate1721(.a(gate291inter11), .b(gate291inter6), .O(gate291inter12));
  nand2 gate1722(.a(gate291inter12), .b(gate291inter1), .O(G860));
nand2 gate292( .a(G824), .b(G825), .O(G873) );
nand2 gate293( .a(G828), .b(G829), .O(G886) );
nand2 gate294( .a(G832), .b(G833), .O(G899) );

  xor2  gate715(.a(G831), .b(G830), .O(gate295inter0));
  nand2 gate716(.a(gate295inter0), .b(s_24), .O(gate295inter1));
  and2  gate717(.a(G831), .b(G830), .O(gate295inter2));
  inv1  gate718(.a(s_24), .O(gate295inter3));
  inv1  gate719(.a(s_25), .O(gate295inter4));
  nand2 gate720(.a(gate295inter4), .b(gate295inter3), .O(gate295inter5));
  nor2  gate721(.a(gate295inter5), .b(gate295inter2), .O(gate295inter6));
  inv1  gate722(.a(G830), .O(gate295inter7));
  inv1  gate723(.a(G831), .O(gate295inter8));
  nand2 gate724(.a(gate295inter8), .b(gate295inter7), .O(gate295inter9));
  nand2 gate725(.a(s_25), .b(gate295inter3), .O(gate295inter10));
  nor2  gate726(.a(gate295inter10), .b(gate295inter9), .O(gate295inter11));
  nor2  gate727(.a(gate295inter11), .b(gate295inter6), .O(gate295inter12));
  nand2 gate728(.a(gate295inter12), .b(gate295inter1), .O(G912));
nand2 gate296( .a(G826), .b(G827), .O(G925) );
inv1 gate297( .a(G834), .O(G938) );
inv1 gate298( .a(G847), .O(G939) );
inv1 gate299( .a(G860), .O(G940) );
inv1 gate300( .a(G834), .O(G941) );
inv1 gate301( .a(G847), .O(G942) );
inv1 gate302( .a(G873), .O(G943) );
inv1 gate303( .a(G834), .O(G944) );
inv1 gate304( .a(G860), .O(G945) );
inv1 gate305( .a(G873), .O(G946) );
inv1 gate306( .a(G847), .O(G947) );
inv1 gate307( .a(G860), .O(G948) );
inv1 gate308( .a(G873), .O(G949) );
inv1 gate309( .a(G886), .O(G950) );
inv1 gate310( .a(G899), .O(G951) );
inv1 gate311( .a(G886), .O(G952) );
inv1 gate312( .a(G912), .O(G953) );
inv1 gate313( .a(G925), .O(G954) );
inv1 gate314( .a(G899), .O(G955) );
inv1 gate315( .a(G925), .O(G956) );
inv1 gate316( .a(G912), .O(G957) );
inv1 gate317( .a(G925), .O(G958) );
inv1 gate318( .a(G886), .O(G959) );
inv1 gate319( .a(G912), .O(G960) );
inv1 gate320( .a(G925), .O(G961) );
inv1 gate321( .a(G886), .O(G962) );
inv1 gate322( .a(G899), .O(G963) );
inv1 gate323( .a(G925), .O(G964) );
inv1 gate324( .a(G912), .O(G965) );
inv1 gate325( .a(G899), .O(G966) );
inv1 gate326( .a(G886), .O(G967) );
inv1 gate327( .a(G912), .O(G968) );
inv1 gate328( .a(G899), .O(G969) );
inv1 gate329( .a(G847), .O(G970) );
inv1 gate330( .a(G873), .O(G971) );
inv1 gate331( .a(G847), .O(G972) );
inv1 gate332( .a(G860), .O(G973) );
inv1 gate333( .a(G834), .O(G974) );
inv1 gate334( .a(G873), .O(G975) );
inv1 gate335( .a(G834), .O(G976) );
inv1 gate336( .a(G860), .O(G977) );
and4 gate337( .a(G938), .b(G939), .c(G940), .d(G873), .O(G978) );
and4 gate338( .a(G941), .b(G942), .c(G860), .d(G943), .O(G979) );
and4 gate339( .a(G944), .b(G847), .c(G945), .d(G946), .O(G980) );
and4 gate340( .a(G834), .b(G947), .c(G948), .d(G949), .O(G981) );
and4 gate341( .a(G958), .b(G959), .c(G960), .d(G899), .O(G982) );
and4 gate342( .a(G961), .b(G962), .c(G912), .d(G963), .O(G983) );
and4 gate343( .a(G964), .b(G886), .c(G965), .d(G966), .O(G984) );
and4 gate344( .a(G925), .b(G967), .c(G968), .d(G969), .O(G985) );
or4 gate345( .a(G978), .b(G979), .c(G980), .d(G981), .O(G986) );
or4 gate346( .a(G982), .b(G983), .c(G984), .d(G985), .O(G991) );
and5 gate347( .a(G925), .b(G950), .c(G912), .d(G951), .e(G986), .O(G996) );
and5 gate348( .a(G925), .b(G952), .c(G953), .d(G899), .e(G986), .O(G1001) );
and5 gate349( .a(G954), .b(G886), .c(G912), .d(G955), .e(G986), .O(G1006) );
and5 gate350( .a(G956), .b(G886), .c(G957), .d(G899), .e(G986), .O(G1011) );
and5 gate351( .a(G834), .b(G970), .c(G860), .d(G971), .e(G991), .O(G1016) );
and5 gate352( .a(G834), .b(G972), .c(G973), .d(G873), .e(G991), .O(G1021) );
and5 gate353( .a(G974), .b(G847), .c(G860), .d(G975), .e(G991), .O(G1026) );
and5 gate354( .a(G976), .b(G847), .c(G977), .d(G873), .e(G991), .O(G1031) );
and2 gate355( .a(G834), .b(G996), .O(G1036) );
and2 gate356( .a(G847), .b(G996), .O(G1039) );
and2 gate357( .a(G860), .b(G996), .O(G1042) );
and2 gate358( .a(G873), .b(G996), .O(G1045) );
and2 gate359( .a(G834), .b(G1001), .O(G1048) );
and2 gate360( .a(G847), .b(G1001), .O(G1051) );
and2 gate361( .a(G860), .b(G1001), .O(G1054) );
and2 gate362( .a(G873), .b(G1001), .O(G1057) );
and2 gate363( .a(G834), .b(G1006), .O(G1060) );
and2 gate364( .a(G847), .b(G1006), .O(G1063) );
and2 gate365( .a(G860), .b(G1006), .O(G1066) );
and2 gate366( .a(G873), .b(G1006), .O(G1069) );
and2 gate367( .a(G834), .b(G1011), .O(G1072) );
and2 gate368( .a(G847), .b(G1011), .O(G1075) );
and2 gate369( .a(G860), .b(G1011), .O(G1078) );
and2 gate370( .a(G873), .b(G1011), .O(G1081) );
and2 gate371( .a(G925), .b(G1016), .O(G1084) );
and2 gate372( .a(G886), .b(G1016), .O(G1087) );
and2 gate373( .a(G912), .b(G1016), .O(G1090) );
and2 gate374( .a(G899), .b(G1016), .O(G1093) );
and2 gate375( .a(G925), .b(G1021), .O(G1096) );
and2 gate376( .a(G886), .b(G1021), .O(G1099) );
and2 gate377( .a(G912), .b(G1021), .O(G1102) );
and2 gate378( .a(G899), .b(G1021), .O(G1105) );
and2 gate379( .a(G925), .b(G1026), .O(G1108) );
and2 gate380( .a(G886), .b(G1026), .O(G1111) );
and2 gate381( .a(G912), .b(G1026), .O(G1114) );
and2 gate382( .a(G899), .b(G1026), .O(G1117) );
and2 gate383( .a(G925), .b(G1031), .O(G1120) );
and2 gate384( .a(G886), .b(G1031), .O(G1123) );
and2 gate385( .a(G912), .b(G1031), .O(G1126) );
and2 gate386( .a(G899), .b(G1031), .O(G1129) );

  xor2  gate2031(.a(G1036), .b(G1), .O(gate387inter0));
  nand2 gate2032(.a(gate387inter0), .b(s_212), .O(gate387inter1));
  and2  gate2033(.a(G1036), .b(G1), .O(gate387inter2));
  inv1  gate2034(.a(s_212), .O(gate387inter3));
  inv1  gate2035(.a(s_213), .O(gate387inter4));
  nand2 gate2036(.a(gate387inter4), .b(gate387inter3), .O(gate387inter5));
  nor2  gate2037(.a(gate387inter5), .b(gate387inter2), .O(gate387inter6));
  inv1  gate2038(.a(G1), .O(gate387inter7));
  inv1  gate2039(.a(G1036), .O(gate387inter8));
  nand2 gate2040(.a(gate387inter8), .b(gate387inter7), .O(gate387inter9));
  nand2 gate2041(.a(s_213), .b(gate387inter3), .O(gate387inter10));
  nor2  gate2042(.a(gate387inter10), .b(gate387inter9), .O(gate387inter11));
  nor2  gate2043(.a(gate387inter11), .b(gate387inter6), .O(gate387inter12));
  nand2 gate2044(.a(gate387inter12), .b(gate387inter1), .O(G1132));
nand2 gate388( .a(G2), .b(G1039), .O(G1135) );
nand2 gate389( .a(G3), .b(G1042), .O(G1138) );
nand2 gate390( .a(G4), .b(G1045), .O(G1141) );
nand2 gate391( .a(G5), .b(G1048), .O(G1144) );
nand2 gate392( .a(G6), .b(G1051), .O(G1147) );

  xor2  gate1457(.a(G1054), .b(G7), .O(gate393inter0));
  nand2 gate1458(.a(gate393inter0), .b(s_130), .O(gate393inter1));
  and2  gate1459(.a(G1054), .b(G7), .O(gate393inter2));
  inv1  gate1460(.a(s_130), .O(gate393inter3));
  inv1  gate1461(.a(s_131), .O(gate393inter4));
  nand2 gate1462(.a(gate393inter4), .b(gate393inter3), .O(gate393inter5));
  nor2  gate1463(.a(gate393inter5), .b(gate393inter2), .O(gate393inter6));
  inv1  gate1464(.a(G7), .O(gate393inter7));
  inv1  gate1465(.a(G1054), .O(gate393inter8));
  nand2 gate1466(.a(gate393inter8), .b(gate393inter7), .O(gate393inter9));
  nand2 gate1467(.a(s_131), .b(gate393inter3), .O(gate393inter10));
  nor2  gate1468(.a(gate393inter10), .b(gate393inter9), .O(gate393inter11));
  nor2  gate1469(.a(gate393inter11), .b(gate393inter6), .O(gate393inter12));
  nand2 gate1470(.a(gate393inter12), .b(gate393inter1), .O(G1150));
nand2 gate394( .a(G8), .b(G1057), .O(G1153) );
nand2 gate395( .a(G9), .b(G1060), .O(G1156) );
nand2 gate396( .a(G10), .b(G1063), .O(G1159) );
nand2 gate397( .a(G11), .b(G1066), .O(G1162) );
nand2 gate398( .a(G12), .b(G1069), .O(G1165) );
nand2 gate399( .a(G13), .b(G1072), .O(G1168) );
nand2 gate400( .a(G14), .b(G1075), .O(G1171) );

  xor2  gate1135(.a(G1078), .b(G15), .O(gate401inter0));
  nand2 gate1136(.a(gate401inter0), .b(s_84), .O(gate401inter1));
  and2  gate1137(.a(G1078), .b(G15), .O(gate401inter2));
  inv1  gate1138(.a(s_84), .O(gate401inter3));
  inv1  gate1139(.a(s_85), .O(gate401inter4));
  nand2 gate1140(.a(gate401inter4), .b(gate401inter3), .O(gate401inter5));
  nor2  gate1141(.a(gate401inter5), .b(gate401inter2), .O(gate401inter6));
  inv1  gate1142(.a(G15), .O(gate401inter7));
  inv1  gate1143(.a(G1078), .O(gate401inter8));
  nand2 gate1144(.a(gate401inter8), .b(gate401inter7), .O(gate401inter9));
  nand2 gate1145(.a(s_85), .b(gate401inter3), .O(gate401inter10));
  nor2  gate1146(.a(gate401inter10), .b(gate401inter9), .O(gate401inter11));
  nor2  gate1147(.a(gate401inter11), .b(gate401inter6), .O(gate401inter12));
  nand2 gate1148(.a(gate401inter12), .b(gate401inter1), .O(G1174));

  xor2  gate2087(.a(G1081), .b(G16), .O(gate402inter0));
  nand2 gate2088(.a(gate402inter0), .b(s_220), .O(gate402inter1));
  and2  gate2089(.a(G1081), .b(G16), .O(gate402inter2));
  inv1  gate2090(.a(s_220), .O(gate402inter3));
  inv1  gate2091(.a(s_221), .O(gate402inter4));
  nand2 gate2092(.a(gate402inter4), .b(gate402inter3), .O(gate402inter5));
  nor2  gate2093(.a(gate402inter5), .b(gate402inter2), .O(gate402inter6));
  inv1  gate2094(.a(G16), .O(gate402inter7));
  inv1  gate2095(.a(G1081), .O(gate402inter8));
  nand2 gate2096(.a(gate402inter8), .b(gate402inter7), .O(gate402inter9));
  nand2 gate2097(.a(s_221), .b(gate402inter3), .O(gate402inter10));
  nor2  gate2098(.a(gate402inter10), .b(gate402inter9), .O(gate402inter11));
  nor2  gate2099(.a(gate402inter11), .b(gate402inter6), .O(gate402inter12));
  nand2 gate2100(.a(gate402inter12), .b(gate402inter1), .O(G1177));
nand2 gate403( .a(G17), .b(G1084), .O(G1180) );

  xor2  gate2073(.a(G1087), .b(G18), .O(gate404inter0));
  nand2 gate2074(.a(gate404inter0), .b(s_218), .O(gate404inter1));
  and2  gate2075(.a(G1087), .b(G18), .O(gate404inter2));
  inv1  gate2076(.a(s_218), .O(gate404inter3));
  inv1  gate2077(.a(s_219), .O(gate404inter4));
  nand2 gate2078(.a(gate404inter4), .b(gate404inter3), .O(gate404inter5));
  nor2  gate2079(.a(gate404inter5), .b(gate404inter2), .O(gate404inter6));
  inv1  gate2080(.a(G18), .O(gate404inter7));
  inv1  gate2081(.a(G1087), .O(gate404inter8));
  nand2 gate2082(.a(gate404inter8), .b(gate404inter7), .O(gate404inter9));
  nand2 gate2083(.a(s_219), .b(gate404inter3), .O(gate404inter10));
  nor2  gate2084(.a(gate404inter10), .b(gate404inter9), .O(gate404inter11));
  nor2  gate2085(.a(gate404inter11), .b(gate404inter6), .O(gate404inter12));
  nand2 gate2086(.a(gate404inter12), .b(gate404inter1), .O(G1183));
nand2 gate405( .a(G19), .b(G1090), .O(G1186) );
nand2 gate406( .a(G20), .b(G1093), .O(G1189) );
nand2 gate407( .a(G21), .b(G1096), .O(G1192) );

  xor2  gate2059(.a(G1099), .b(G22), .O(gate408inter0));
  nand2 gate2060(.a(gate408inter0), .b(s_216), .O(gate408inter1));
  and2  gate2061(.a(G1099), .b(G22), .O(gate408inter2));
  inv1  gate2062(.a(s_216), .O(gate408inter3));
  inv1  gate2063(.a(s_217), .O(gate408inter4));
  nand2 gate2064(.a(gate408inter4), .b(gate408inter3), .O(gate408inter5));
  nor2  gate2065(.a(gate408inter5), .b(gate408inter2), .O(gate408inter6));
  inv1  gate2066(.a(G22), .O(gate408inter7));
  inv1  gate2067(.a(G1099), .O(gate408inter8));
  nand2 gate2068(.a(gate408inter8), .b(gate408inter7), .O(gate408inter9));
  nand2 gate2069(.a(s_217), .b(gate408inter3), .O(gate408inter10));
  nor2  gate2070(.a(gate408inter10), .b(gate408inter9), .O(gate408inter11));
  nor2  gate2071(.a(gate408inter11), .b(gate408inter6), .O(gate408inter12));
  nand2 gate2072(.a(gate408inter12), .b(gate408inter1), .O(G1195));

  xor2  gate659(.a(G1102), .b(G23), .O(gate409inter0));
  nand2 gate660(.a(gate409inter0), .b(s_16), .O(gate409inter1));
  and2  gate661(.a(G1102), .b(G23), .O(gate409inter2));
  inv1  gate662(.a(s_16), .O(gate409inter3));
  inv1  gate663(.a(s_17), .O(gate409inter4));
  nand2 gate664(.a(gate409inter4), .b(gate409inter3), .O(gate409inter5));
  nor2  gate665(.a(gate409inter5), .b(gate409inter2), .O(gate409inter6));
  inv1  gate666(.a(G23), .O(gate409inter7));
  inv1  gate667(.a(G1102), .O(gate409inter8));
  nand2 gate668(.a(gate409inter8), .b(gate409inter7), .O(gate409inter9));
  nand2 gate669(.a(s_17), .b(gate409inter3), .O(gate409inter10));
  nor2  gate670(.a(gate409inter10), .b(gate409inter9), .O(gate409inter11));
  nor2  gate671(.a(gate409inter11), .b(gate409inter6), .O(gate409inter12));
  nand2 gate672(.a(gate409inter12), .b(gate409inter1), .O(G1198));

  xor2  gate1415(.a(G1105), .b(G24), .O(gate410inter0));
  nand2 gate1416(.a(gate410inter0), .b(s_124), .O(gate410inter1));
  and2  gate1417(.a(G1105), .b(G24), .O(gate410inter2));
  inv1  gate1418(.a(s_124), .O(gate410inter3));
  inv1  gate1419(.a(s_125), .O(gate410inter4));
  nand2 gate1420(.a(gate410inter4), .b(gate410inter3), .O(gate410inter5));
  nor2  gate1421(.a(gate410inter5), .b(gate410inter2), .O(gate410inter6));
  inv1  gate1422(.a(G24), .O(gate410inter7));
  inv1  gate1423(.a(G1105), .O(gate410inter8));
  nand2 gate1424(.a(gate410inter8), .b(gate410inter7), .O(gate410inter9));
  nand2 gate1425(.a(s_125), .b(gate410inter3), .O(gate410inter10));
  nor2  gate1426(.a(gate410inter10), .b(gate410inter9), .O(gate410inter11));
  nor2  gate1427(.a(gate410inter11), .b(gate410inter6), .O(gate410inter12));
  nand2 gate1428(.a(gate410inter12), .b(gate410inter1), .O(G1201));
nand2 gate411( .a(G25), .b(G1108), .O(G1204) );

  xor2  gate2115(.a(G1111), .b(G26), .O(gate412inter0));
  nand2 gate2116(.a(gate412inter0), .b(s_224), .O(gate412inter1));
  and2  gate2117(.a(G1111), .b(G26), .O(gate412inter2));
  inv1  gate2118(.a(s_224), .O(gate412inter3));
  inv1  gate2119(.a(s_225), .O(gate412inter4));
  nand2 gate2120(.a(gate412inter4), .b(gate412inter3), .O(gate412inter5));
  nor2  gate2121(.a(gate412inter5), .b(gate412inter2), .O(gate412inter6));
  inv1  gate2122(.a(G26), .O(gate412inter7));
  inv1  gate2123(.a(G1111), .O(gate412inter8));
  nand2 gate2124(.a(gate412inter8), .b(gate412inter7), .O(gate412inter9));
  nand2 gate2125(.a(s_225), .b(gate412inter3), .O(gate412inter10));
  nor2  gate2126(.a(gate412inter10), .b(gate412inter9), .O(gate412inter11));
  nor2  gate2127(.a(gate412inter11), .b(gate412inter6), .O(gate412inter12));
  nand2 gate2128(.a(gate412inter12), .b(gate412inter1), .O(G1207));
nand2 gate413( .a(G27), .b(G1114), .O(G1210) );
nand2 gate414( .a(G28), .b(G1117), .O(G1213) );

  xor2  gate1807(.a(G1120), .b(G29), .O(gate415inter0));
  nand2 gate1808(.a(gate415inter0), .b(s_180), .O(gate415inter1));
  and2  gate1809(.a(G1120), .b(G29), .O(gate415inter2));
  inv1  gate1810(.a(s_180), .O(gate415inter3));
  inv1  gate1811(.a(s_181), .O(gate415inter4));
  nand2 gate1812(.a(gate415inter4), .b(gate415inter3), .O(gate415inter5));
  nor2  gate1813(.a(gate415inter5), .b(gate415inter2), .O(gate415inter6));
  inv1  gate1814(.a(G29), .O(gate415inter7));
  inv1  gate1815(.a(G1120), .O(gate415inter8));
  nand2 gate1816(.a(gate415inter8), .b(gate415inter7), .O(gate415inter9));
  nand2 gate1817(.a(s_181), .b(gate415inter3), .O(gate415inter10));
  nor2  gate1818(.a(gate415inter10), .b(gate415inter9), .O(gate415inter11));
  nor2  gate1819(.a(gate415inter11), .b(gate415inter6), .O(gate415inter12));
  nand2 gate1820(.a(gate415inter12), .b(gate415inter1), .O(G1216));
nand2 gate416( .a(G30), .b(G1123), .O(G1219) );

  xor2  gate1149(.a(G1126), .b(G31), .O(gate417inter0));
  nand2 gate1150(.a(gate417inter0), .b(s_86), .O(gate417inter1));
  and2  gate1151(.a(G1126), .b(G31), .O(gate417inter2));
  inv1  gate1152(.a(s_86), .O(gate417inter3));
  inv1  gate1153(.a(s_87), .O(gate417inter4));
  nand2 gate1154(.a(gate417inter4), .b(gate417inter3), .O(gate417inter5));
  nor2  gate1155(.a(gate417inter5), .b(gate417inter2), .O(gate417inter6));
  inv1  gate1156(.a(G31), .O(gate417inter7));
  inv1  gate1157(.a(G1126), .O(gate417inter8));
  nand2 gate1158(.a(gate417inter8), .b(gate417inter7), .O(gate417inter9));
  nand2 gate1159(.a(s_87), .b(gate417inter3), .O(gate417inter10));
  nor2  gate1160(.a(gate417inter10), .b(gate417inter9), .O(gate417inter11));
  nor2  gate1161(.a(gate417inter11), .b(gate417inter6), .O(gate417inter12));
  nand2 gate1162(.a(gate417inter12), .b(gate417inter1), .O(G1222));

  xor2  gate729(.a(G1129), .b(G32), .O(gate418inter0));
  nand2 gate730(.a(gate418inter0), .b(s_26), .O(gate418inter1));
  and2  gate731(.a(G1129), .b(G32), .O(gate418inter2));
  inv1  gate732(.a(s_26), .O(gate418inter3));
  inv1  gate733(.a(s_27), .O(gate418inter4));
  nand2 gate734(.a(gate418inter4), .b(gate418inter3), .O(gate418inter5));
  nor2  gate735(.a(gate418inter5), .b(gate418inter2), .O(gate418inter6));
  inv1  gate736(.a(G32), .O(gate418inter7));
  inv1  gate737(.a(G1129), .O(gate418inter8));
  nand2 gate738(.a(gate418inter8), .b(gate418inter7), .O(gate418inter9));
  nand2 gate739(.a(s_27), .b(gate418inter3), .O(gate418inter10));
  nor2  gate740(.a(gate418inter10), .b(gate418inter9), .O(gate418inter11));
  nor2  gate741(.a(gate418inter11), .b(gate418inter6), .O(gate418inter12));
  nand2 gate742(.a(gate418inter12), .b(gate418inter1), .O(G1225));

  xor2  gate589(.a(G1132), .b(G1), .O(gate419inter0));
  nand2 gate590(.a(gate419inter0), .b(s_6), .O(gate419inter1));
  and2  gate591(.a(G1132), .b(G1), .O(gate419inter2));
  inv1  gate592(.a(s_6), .O(gate419inter3));
  inv1  gate593(.a(s_7), .O(gate419inter4));
  nand2 gate594(.a(gate419inter4), .b(gate419inter3), .O(gate419inter5));
  nor2  gate595(.a(gate419inter5), .b(gate419inter2), .O(gate419inter6));
  inv1  gate596(.a(G1), .O(gate419inter7));
  inv1  gate597(.a(G1132), .O(gate419inter8));
  nand2 gate598(.a(gate419inter8), .b(gate419inter7), .O(gate419inter9));
  nand2 gate599(.a(s_7), .b(gate419inter3), .O(gate419inter10));
  nor2  gate600(.a(gate419inter10), .b(gate419inter9), .O(gate419inter11));
  nor2  gate601(.a(gate419inter11), .b(gate419inter6), .O(gate419inter12));
  nand2 gate602(.a(gate419inter12), .b(gate419inter1), .O(G1228));

  xor2  gate1849(.a(G1132), .b(G1036), .O(gate420inter0));
  nand2 gate1850(.a(gate420inter0), .b(s_186), .O(gate420inter1));
  and2  gate1851(.a(G1132), .b(G1036), .O(gate420inter2));
  inv1  gate1852(.a(s_186), .O(gate420inter3));
  inv1  gate1853(.a(s_187), .O(gate420inter4));
  nand2 gate1854(.a(gate420inter4), .b(gate420inter3), .O(gate420inter5));
  nor2  gate1855(.a(gate420inter5), .b(gate420inter2), .O(gate420inter6));
  inv1  gate1856(.a(G1036), .O(gate420inter7));
  inv1  gate1857(.a(G1132), .O(gate420inter8));
  nand2 gate1858(.a(gate420inter8), .b(gate420inter7), .O(gate420inter9));
  nand2 gate1859(.a(s_187), .b(gate420inter3), .O(gate420inter10));
  nor2  gate1860(.a(gate420inter10), .b(gate420inter9), .O(gate420inter11));
  nor2  gate1861(.a(gate420inter11), .b(gate420inter6), .O(gate420inter12));
  nand2 gate1862(.a(gate420inter12), .b(gate420inter1), .O(G1229));
nand2 gate421( .a(G2), .b(G1135), .O(G1230) );
nand2 gate422( .a(G1039), .b(G1135), .O(G1231) );

  xor2  gate1555(.a(G1138), .b(G3), .O(gate423inter0));
  nand2 gate1556(.a(gate423inter0), .b(s_144), .O(gate423inter1));
  and2  gate1557(.a(G1138), .b(G3), .O(gate423inter2));
  inv1  gate1558(.a(s_144), .O(gate423inter3));
  inv1  gate1559(.a(s_145), .O(gate423inter4));
  nand2 gate1560(.a(gate423inter4), .b(gate423inter3), .O(gate423inter5));
  nor2  gate1561(.a(gate423inter5), .b(gate423inter2), .O(gate423inter6));
  inv1  gate1562(.a(G3), .O(gate423inter7));
  inv1  gate1563(.a(G1138), .O(gate423inter8));
  nand2 gate1564(.a(gate423inter8), .b(gate423inter7), .O(gate423inter9));
  nand2 gate1565(.a(s_145), .b(gate423inter3), .O(gate423inter10));
  nor2  gate1566(.a(gate423inter10), .b(gate423inter9), .O(gate423inter11));
  nor2  gate1567(.a(gate423inter11), .b(gate423inter6), .O(gate423inter12));
  nand2 gate1568(.a(gate423inter12), .b(gate423inter1), .O(G1232));

  xor2  gate1989(.a(G1138), .b(G1042), .O(gate424inter0));
  nand2 gate1990(.a(gate424inter0), .b(s_206), .O(gate424inter1));
  and2  gate1991(.a(G1138), .b(G1042), .O(gate424inter2));
  inv1  gate1992(.a(s_206), .O(gate424inter3));
  inv1  gate1993(.a(s_207), .O(gate424inter4));
  nand2 gate1994(.a(gate424inter4), .b(gate424inter3), .O(gate424inter5));
  nor2  gate1995(.a(gate424inter5), .b(gate424inter2), .O(gate424inter6));
  inv1  gate1996(.a(G1042), .O(gate424inter7));
  inv1  gate1997(.a(G1138), .O(gate424inter8));
  nand2 gate1998(.a(gate424inter8), .b(gate424inter7), .O(gate424inter9));
  nand2 gate1999(.a(s_207), .b(gate424inter3), .O(gate424inter10));
  nor2  gate2000(.a(gate424inter10), .b(gate424inter9), .O(gate424inter11));
  nor2  gate2001(.a(gate424inter11), .b(gate424inter6), .O(gate424inter12));
  nand2 gate2002(.a(gate424inter12), .b(gate424inter1), .O(G1233));

  xor2  gate911(.a(G1141), .b(G4), .O(gate425inter0));
  nand2 gate912(.a(gate425inter0), .b(s_52), .O(gate425inter1));
  and2  gate913(.a(G1141), .b(G4), .O(gate425inter2));
  inv1  gate914(.a(s_52), .O(gate425inter3));
  inv1  gate915(.a(s_53), .O(gate425inter4));
  nand2 gate916(.a(gate425inter4), .b(gate425inter3), .O(gate425inter5));
  nor2  gate917(.a(gate425inter5), .b(gate425inter2), .O(gate425inter6));
  inv1  gate918(.a(G4), .O(gate425inter7));
  inv1  gate919(.a(G1141), .O(gate425inter8));
  nand2 gate920(.a(gate425inter8), .b(gate425inter7), .O(gate425inter9));
  nand2 gate921(.a(s_53), .b(gate425inter3), .O(gate425inter10));
  nor2  gate922(.a(gate425inter10), .b(gate425inter9), .O(gate425inter11));
  nor2  gate923(.a(gate425inter11), .b(gate425inter6), .O(gate425inter12));
  nand2 gate924(.a(gate425inter12), .b(gate425inter1), .O(G1234));

  xor2  gate1023(.a(G1141), .b(G1045), .O(gate426inter0));
  nand2 gate1024(.a(gate426inter0), .b(s_68), .O(gate426inter1));
  and2  gate1025(.a(G1141), .b(G1045), .O(gate426inter2));
  inv1  gate1026(.a(s_68), .O(gate426inter3));
  inv1  gate1027(.a(s_69), .O(gate426inter4));
  nand2 gate1028(.a(gate426inter4), .b(gate426inter3), .O(gate426inter5));
  nor2  gate1029(.a(gate426inter5), .b(gate426inter2), .O(gate426inter6));
  inv1  gate1030(.a(G1045), .O(gate426inter7));
  inv1  gate1031(.a(G1141), .O(gate426inter8));
  nand2 gate1032(.a(gate426inter8), .b(gate426inter7), .O(gate426inter9));
  nand2 gate1033(.a(s_69), .b(gate426inter3), .O(gate426inter10));
  nor2  gate1034(.a(gate426inter10), .b(gate426inter9), .O(gate426inter11));
  nor2  gate1035(.a(gate426inter11), .b(gate426inter6), .O(gate426inter12));
  nand2 gate1036(.a(gate426inter12), .b(gate426inter1), .O(G1235));
nand2 gate427( .a(G5), .b(G1144), .O(G1236) );
nand2 gate428( .a(G1048), .b(G1144), .O(G1237) );
nand2 gate429( .a(G6), .b(G1147), .O(G1238) );
nand2 gate430( .a(G1051), .b(G1147), .O(G1239) );
nand2 gate431( .a(G7), .b(G1150), .O(G1240) );
nand2 gate432( .a(G1054), .b(G1150), .O(G1241) );

  xor2  gate1429(.a(G1153), .b(G8), .O(gate433inter0));
  nand2 gate1430(.a(gate433inter0), .b(s_126), .O(gate433inter1));
  and2  gate1431(.a(G1153), .b(G8), .O(gate433inter2));
  inv1  gate1432(.a(s_126), .O(gate433inter3));
  inv1  gate1433(.a(s_127), .O(gate433inter4));
  nand2 gate1434(.a(gate433inter4), .b(gate433inter3), .O(gate433inter5));
  nor2  gate1435(.a(gate433inter5), .b(gate433inter2), .O(gate433inter6));
  inv1  gate1436(.a(G8), .O(gate433inter7));
  inv1  gate1437(.a(G1153), .O(gate433inter8));
  nand2 gate1438(.a(gate433inter8), .b(gate433inter7), .O(gate433inter9));
  nand2 gate1439(.a(s_127), .b(gate433inter3), .O(gate433inter10));
  nor2  gate1440(.a(gate433inter10), .b(gate433inter9), .O(gate433inter11));
  nor2  gate1441(.a(gate433inter11), .b(gate433inter6), .O(gate433inter12));
  nand2 gate1442(.a(gate433inter12), .b(gate433inter1), .O(G1242));
nand2 gate434( .a(G1057), .b(G1153), .O(G1243) );
nand2 gate435( .a(G9), .b(G1156), .O(G1244) );
nand2 gate436( .a(G1060), .b(G1156), .O(G1245) );
nand2 gate437( .a(G10), .b(G1159), .O(G1246) );
nand2 gate438( .a(G1063), .b(G1159), .O(G1247) );
nand2 gate439( .a(G11), .b(G1162), .O(G1248) );
nand2 gate440( .a(G1066), .b(G1162), .O(G1249) );
nand2 gate441( .a(G12), .b(G1165), .O(G1250) );

  xor2  gate897(.a(G1165), .b(G1069), .O(gate442inter0));
  nand2 gate898(.a(gate442inter0), .b(s_50), .O(gate442inter1));
  and2  gate899(.a(G1165), .b(G1069), .O(gate442inter2));
  inv1  gate900(.a(s_50), .O(gate442inter3));
  inv1  gate901(.a(s_51), .O(gate442inter4));
  nand2 gate902(.a(gate442inter4), .b(gate442inter3), .O(gate442inter5));
  nor2  gate903(.a(gate442inter5), .b(gate442inter2), .O(gate442inter6));
  inv1  gate904(.a(G1069), .O(gate442inter7));
  inv1  gate905(.a(G1165), .O(gate442inter8));
  nand2 gate906(.a(gate442inter8), .b(gate442inter7), .O(gate442inter9));
  nand2 gate907(.a(s_51), .b(gate442inter3), .O(gate442inter10));
  nor2  gate908(.a(gate442inter10), .b(gate442inter9), .O(gate442inter11));
  nor2  gate909(.a(gate442inter11), .b(gate442inter6), .O(gate442inter12));
  nand2 gate910(.a(gate442inter12), .b(gate442inter1), .O(G1251));
nand2 gate443( .a(G13), .b(G1168), .O(G1252) );
nand2 gate444( .a(G1072), .b(G1168), .O(G1253) );
nand2 gate445( .a(G14), .b(G1171), .O(G1254) );
nand2 gate446( .a(G1075), .b(G1171), .O(G1255) );
nand2 gate447( .a(G15), .b(G1174), .O(G1256) );
nand2 gate448( .a(G1078), .b(G1174), .O(G1257) );

  xor2  gate1485(.a(G1177), .b(G16), .O(gate449inter0));
  nand2 gate1486(.a(gate449inter0), .b(s_134), .O(gate449inter1));
  and2  gate1487(.a(G1177), .b(G16), .O(gate449inter2));
  inv1  gate1488(.a(s_134), .O(gate449inter3));
  inv1  gate1489(.a(s_135), .O(gate449inter4));
  nand2 gate1490(.a(gate449inter4), .b(gate449inter3), .O(gate449inter5));
  nor2  gate1491(.a(gate449inter5), .b(gate449inter2), .O(gate449inter6));
  inv1  gate1492(.a(G16), .O(gate449inter7));
  inv1  gate1493(.a(G1177), .O(gate449inter8));
  nand2 gate1494(.a(gate449inter8), .b(gate449inter7), .O(gate449inter9));
  nand2 gate1495(.a(s_135), .b(gate449inter3), .O(gate449inter10));
  nor2  gate1496(.a(gate449inter10), .b(gate449inter9), .O(gate449inter11));
  nor2  gate1497(.a(gate449inter11), .b(gate449inter6), .O(gate449inter12));
  nand2 gate1498(.a(gate449inter12), .b(gate449inter1), .O(G1258));
nand2 gate450( .a(G1081), .b(G1177), .O(G1259) );
nand2 gate451( .a(G17), .b(G1180), .O(G1260) );
nand2 gate452( .a(G1084), .b(G1180), .O(G1261) );
nand2 gate453( .a(G18), .b(G1183), .O(G1262) );
nand2 gate454( .a(G1087), .b(G1183), .O(G1263) );

  xor2  gate1933(.a(G1186), .b(G19), .O(gate455inter0));
  nand2 gate1934(.a(gate455inter0), .b(s_198), .O(gate455inter1));
  and2  gate1935(.a(G1186), .b(G19), .O(gate455inter2));
  inv1  gate1936(.a(s_198), .O(gate455inter3));
  inv1  gate1937(.a(s_199), .O(gate455inter4));
  nand2 gate1938(.a(gate455inter4), .b(gate455inter3), .O(gate455inter5));
  nor2  gate1939(.a(gate455inter5), .b(gate455inter2), .O(gate455inter6));
  inv1  gate1940(.a(G19), .O(gate455inter7));
  inv1  gate1941(.a(G1186), .O(gate455inter8));
  nand2 gate1942(.a(gate455inter8), .b(gate455inter7), .O(gate455inter9));
  nand2 gate1943(.a(s_199), .b(gate455inter3), .O(gate455inter10));
  nor2  gate1944(.a(gate455inter10), .b(gate455inter9), .O(gate455inter11));
  nor2  gate1945(.a(gate455inter11), .b(gate455inter6), .O(gate455inter12));
  nand2 gate1946(.a(gate455inter12), .b(gate455inter1), .O(G1264));
nand2 gate456( .a(G1090), .b(G1186), .O(G1265) );
nand2 gate457( .a(G20), .b(G1189), .O(G1266) );
nand2 gate458( .a(G1093), .b(G1189), .O(G1267) );

  xor2  gate1737(.a(G1192), .b(G21), .O(gate459inter0));
  nand2 gate1738(.a(gate459inter0), .b(s_170), .O(gate459inter1));
  and2  gate1739(.a(G1192), .b(G21), .O(gate459inter2));
  inv1  gate1740(.a(s_170), .O(gate459inter3));
  inv1  gate1741(.a(s_171), .O(gate459inter4));
  nand2 gate1742(.a(gate459inter4), .b(gate459inter3), .O(gate459inter5));
  nor2  gate1743(.a(gate459inter5), .b(gate459inter2), .O(gate459inter6));
  inv1  gate1744(.a(G21), .O(gate459inter7));
  inv1  gate1745(.a(G1192), .O(gate459inter8));
  nand2 gate1746(.a(gate459inter8), .b(gate459inter7), .O(gate459inter9));
  nand2 gate1747(.a(s_171), .b(gate459inter3), .O(gate459inter10));
  nor2  gate1748(.a(gate459inter10), .b(gate459inter9), .O(gate459inter11));
  nor2  gate1749(.a(gate459inter11), .b(gate459inter6), .O(gate459inter12));
  nand2 gate1750(.a(gate459inter12), .b(gate459inter1), .O(G1268));
nand2 gate460( .a(G1096), .b(G1192), .O(G1269) );

  xor2  gate1877(.a(G1195), .b(G22), .O(gate461inter0));
  nand2 gate1878(.a(gate461inter0), .b(s_190), .O(gate461inter1));
  and2  gate1879(.a(G1195), .b(G22), .O(gate461inter2));
  inv1  gate1880(.a(s_190), .O(gate461inter3));
  inv1  gate1881(.a(s_191), .O(gate461inter4));
  nand2 gate1882(.a(gate461inter4), .b(gate461inter3), .O(gate461inter5));
  nor2  gate1883(.a(gate461inter5), .b(gate461inter2), .O(gate461inter6));
  inv1  gate1884(.a(G22), .O(gate461inter7));
  inv1  gate1885(.a(G1195), .O(gate461inter8));
  nand2 gate1886(.a(gate461inter8), .b(gate461inter7), .O(gate461inter9));
  nand2 gate1887(.a(s_191), .b(gate461inter3), .O(gate461inter10));
  nor2  gate1888(.a(gate461inter10), .b(gate461inter9), .O(gate461inter11));
  nor2  gate1889(.a(gate461inter11), .b(gate461inter6), .O(gate461inter12));
  nand2 gate1890(.a(gate461inter12), .b(gate461inter1), .O(G1270));

  xor2  gate1387(.a(G1195), .b(G1099), .O(gate462inter0));
  nand2 gate1388(.a(gate462inter0), .b(s_120), .O(gate462inter1));
  and2  gate1389(.a(G1195), .b(G1099), .O(gate462inter2));
  inv1  gate1390(.a(s_120), .O(gate462inter3));
  inv1  gate1391(.a(s_121), .O(gate462inter4));
  nand2 gate1392(.a(gate462inter4), .b(gate462inter3), .O(gate462inter5));
  nor2  gate1393(.a(gate462inter5), .b(gate462inter2), .O(gate462inter6));
  inv1  gate1394(.a(G1099), .O(gate462inter7));
  inv1  gate1395(.a(G1195), .O(gate462inter8));
  nand2 gate1396(.a(gate462inter8), .b(gate462inter7), .O(gate462inter9));
  nand2 gate1397(.a(s_121), .b(gate462inter3), .O(gate462inter10));
  nor2  gate1398(.a(gate462inter10), .b(gate462inter9), .O(gate462inter11));
  nor2  gate1399(.a(gate462inter11), .b(gate462inter6), .O(gate462inter12));
  nand2 gate1400(.a(gate462inter12), .b(gate462inter1), .O(G1271));
nand2 gate463( .a(G23), .b(G1198), .O(G1272) );
nand2 gate464( .a(G1102), .b(G1198), .O(G1273) );
nand2 gate465( .a(G24), .b(G1201), .O(G1274) );

  xor2  gate813(.a(G1201), .b(G1105), .O(gate466inter0));
  nand2 gate814(.a(gate466inter0), .b(s_38), .O(gate466inter1));
  and2  gate815(.a(G1201), .b(G1105), .O(gate466inter2));
  inv1  gate816(.a(s_38), .O(gate466inter3));
  inv1  gate817(.a(s_39), .O(gate466inter4));
  nand2 gate818(.a(gate466inter4), .b(gate466inter3), .O(gate466inter5));
  nor2  gate819(.a(gate466inter5), .b(gate466inter2), .O(gate466inter6));
  inv1  gate820(.a(G1105), .O(gate466inter7));
  inv1  gate821(.a(G1201), .O(gate466inter8));
  nand2 gate822(.a(gate466inter8), .b(gate466inter7), .O(gate466inter9));
  nand2 gate823(.a(s_39), .b(gate466inter3), .O(gate466inter10));
  nor2  gate824(.a(gate466inter10), .b(gate466inter9), .O(gate466inter11));
  nor2  gate825(.a(gate466inter11), .b(gate466inter6), .O(gate466inter12));
  nand2 gate826(.a(gate466inter12), .b(gate466inter1), .O(G1275));

  xor2  gate2129(.a(G1204), .b(G25), .O(gate467inter0));
  nand2 gate2130(.a(gate467inter0), .b(s_226), .O(gate467inter1));
  and2  gate2131(.a(G1204), .b(G25), .O(gate467inter2));
  inv1  gate2132(.a(s_226), .O(gate467inter3));
  inv1  gate2133(.a(s_227), .O(gate467inter4));
  nand2 gate2134(.a(gate467inter4), .b(gate467inter3), .O(gate467inter5));
  nor2  gate2135(.a(gate467inter5), .b(gate467inter2), .O(gate467inter6));
  inv1  gate2136(.a(G25), .O(gate467inter7));
  inv1  gate2137(.a(G1204), .O(gate467inter8));
  nand2 gate2138(.a(gate467inter8), .b(gate467inter7), .O(gate467inter9));
  nand2 gate2139(.a(s_227), .b(gate467inter3), .O(gate467inter10));
  nor2  gate2140(.a(gate467inter10), .b(gate467inter9), .O(gate467inter11));
  nor2  gate2141(.a(gate467inter11), .b(gate467inter6), .O(gate467inter12));
  nand2 gate2142(.a(gate467inter12), .b(gate467inter1), .O(G1276));
nand2 gate468( .a(G1108), .b(G1204), .O(G1277) );
nand2 gate469( .a(G26), .b(G1207), .O(G1278) );
nand2 gate470( .a(G1111), .b(G1207), .O(G1279) );

  xor2  gate1093(.a(G1210), .b(G27), .O(gate471inter0));
  nand2 gate1094(.a(gate471inter0), .b(s_78), .O(gate471inter1));
  and2  gate1095(.a(G1210), .b(G27), .O(gate471inter2));
  inv1  gate1096(.a(s_78), .O(gate471inter3));
  inv1  gate1097(.a(s_79), .O(gate471inter4));
  nand2 gate1098(.a(gate471inter4), .b(gate471inter3), .O(gate471inter5));
  nor2  gate1099(.a(gate471inter5), .b(gate471inter2), .O(gate471inter6));
  inv1  gate1100(.a(G27), .O(gate471inter7));
  inv1  gate1101(.a(G1210), .O(gate471inter8));
  nand2 gate1102(.a(gate471inter8), .b(gate471inter7), .O(gate471inter9));
  nand2 gate1103(.a(s_79), .b(gate471inter3), .O(gate471inter10));
  nor2  gate1104(.a(gate471inter10), .b(gate471inter9), .O(gate471inter11));
  nor2  gate1105(.a(gate471inter11), .b(gate471inter6), .O(gate471inter12));
  nand2 gate1106(.a(gate471inter12), .b(gate471inter1), .O(G1280));

  xor2  gate701(.a(G1210), .b(G1114), .O(gate472inter0));
  nand2 gate702(.a(gate472inter0), .b(s_22), .O(gate472inter1));
  and2  gate703(.a(G1210), .b(G1114), .O(gate472inter2));
  inv1  gate704(.a(s_22), .O(gate472inter3));
  inv1  gate705(.a(s_23), .O(gate472inter4));
  nand2 gate706(.a(gate472inter4), .b(gate472inter3), .O(gate472inter5));
  nor2  gate707(.a(gate472inter5), .b(gate472inter2), .O(gate472inter6));
  inv1  gate708(.a(G1114), .O(gate472inter7));
  inv1  gate709(.a(G1210), .O(gate472inter8));
  nand2 gate710(.a(gate472inter8), .b(gate472inter7), .O(gate472inter9));
  nand2 gate711(.a(s_23), .b(gate472inter3), .O(gate472inter10));
  nor2  gate712(.a(gate472inter10), .b(gate472inter9), .O(gate472inter11));
  nor2  gate713(.a(gate472inter11), .b(gate472inter6), .O(gate472inter12));
  nand2 gate714(.a(gate472inter12), .b(gate472inter1), .O(G1281));

  xor2  gate1261(.a(G1213), .b(G28), .O(gate473inter0));
  nand2 gate1262(.a(gate473inter0), .b(s_102), .O(gate473inter1));
  and2  gate1263(.a(G1213), .b(G28), .O(gate473inter2));
  inv1  gate1264(.a(s_102), .O(gate473inter3));
  inv1  gate1265(.a(s_103), .O(gate473inter4));
  nand2 gate1266(.a(gate473inter4), .b(gate473inter3), .O(gate473inter5));
  nor2  gate1267(.a(gate473inter5), .b(gate473inter2), .O(gate473inter6));
  inv1  gate1268(.a(G28), .O(gate473inter7));
  inv1  gate1269(.a(G1213), .O(gate473inter8));
  nand2 gate1270(.a(gate473inter8), .b(gate473inter7), .O(gate473inter9));
  nand2 gate1271(.a(s_103), .b(gate473inter3), .O(gate473inter10));
  nor2  gate1272(.a(gate473inter10), .b(gate473inter9), .O(gate473inter11));
  nor2  gate1273(.a(gate473inter11), .b(gate473inter6), .O(gate473inter12));
  nand2 gate1274(.a(gate473inter12), .b(gate473inter1), .O(G1282));
nand2 gate474( .a(G1117), .b(G1213), .O(G1283) );

  xor2  gate883(.a(G1216), .b(G29), .O(gate475inter0));
  nand2 gate884(.a(gate475inter0), .b(s_48), .O(gate475inter1));
  and2  gate885(.a(G1216), .b(G29), .O(gate475inter2));
  inv1  gate886(.a(s_48), .O(gate475inter3));
  inv1  gate887(.a(s_49), .O(gate475inter4));
  nand2 gate888(.a(gate475inter4), .b(gate475inter3), .O(gate475inter5));
  nor2  gate889(.a(gate475inter5), .b(gate475inter2), .O(gate475inter6));
  inv1  gate890(.a(G29), .O(gate475inter7));
  inv1  gate891(.a(G1216), .O(gate475inter8));
  nand2 gate892(.a(gate475inter8), .b(gate475inter7), .O(gate475inter9));
  nand2 gate893(.a(s_49), .b(gate475inter3), .O(gate475inter10));
  nor2  gate894(.a(gate475inter10), .b(gate475inter9), .O(gate475inter11));
  nor2  gate895(.a(gate475inter11), .b(gate475inter6), .O(gate475inter12));
  nand2 gate896(.a(gate475inter12), .b(gate475inter1), .O(G1284));
nand2 gate476( .a(G1120), .b(G1216), .O(G1285) );

  xor2  gate1639(.a(G1219), .b(G30), .O(gate477inter0));
  nand2 gate1640(.a(gate477inter0), .b(s_156), .O(gate477inter1));
  and2  gate1641(.a(G1219), .b(G30), .O(gate477inter2));
  inv1  gate1642(.a(s_156), .O(gate477inter3));
  inv1  gate1643(.a(s_157), .O(gate477inter4));
  nand2 gate1644(.a(gate477inter4), .b(gate477inter3), .O(gate477inter5));
  nor2  gate1645(.a(gate477inter5), .b(gate477inter2), .O(gate477inter6));
  inv1  gate1646(.a(G30), .O(gate477inter7));
  inv1  gate1647(.a(G1219), .O(gate477inter8));
  nand2 gate1648(.a(gate477inter8), .b(gate477inter7), .O(gate477inter9));
  nand2 gate1649(.a(s_157), .b(gate477inter3), .O(gate477inter10));
  nor2  gate1650(.a(gate477inter10), .b(gate477inter9), .O(gate477inter11));
  nor2  gate1651(.a(gate477inter11), .b(gate477inter6), .O(gate477inter12));
  nand2 gate1652(.a(gate477inter12), .b(gate477inter1), .O(G1286));
nand2 gate478( .a(G1123), .b(G1219), .O(G1287) );
nand2 gate479( .a(G31), .b(G1222), .O(G1288) );

  xor2  gate2185(.a(G1222), .b(G1126), .O(gate480inter0));
  nand2 gate2186(.a(gate480inter0), .b(s_234), .O(gate480inter1));
  and2  gate2187(.a(G1222), .b(G1126), .O(gate480inter2));
  inv1  gate2188(.a(s_234), .O(gate480inter3));
  inv1  gate2189(.a(s_235), .O(gate480inter4));
  nand2 gate2190(.a(gate480inter4), .b(gate480inter3), .O(gate480inter5));
  nor2  gate2191(.a(gate480inter5), .b(gate480inter2), .O(gate480inter6));
  inv1  gate2192(.a(G1126), .O(gate480inter7));
  inv1  gate2193(.a(G1222), .O(gate480inter8));
  nand2 gate2194(.a(gate480inter8), .b(gate480inter7), .O(gate480inter9));
  nand2 gate2195(.a(s_235), .b(gate480inter3), .O(gate480inter10));
  nor2  gate2196(.a(gate480inter10), .b(gate480inter9), .O(gate480inter11));
  nor2  gate2197(.a(gate480inter11), .b(gate480inter6), .O(gate480inter12));
  nand2 gate2198(.a(gate480inter12), .b(gate480inter1), .O(G1289));
nand2 gate481( .a(G32), .b(G1225), .O(G1290) );

  xor2  gate1695(.a(G1225), .b(G1129), .O(gate482inter0));
  nand2 gate1696(.a(gate482inter0), .b(s_164), .O(gate482inter1));
  and2  gate1697(.a(G1225), .b(G1129), .O(gate482inter2));
  inv1  gate1698(.a(s_164), .O(gate482inter3));
  inv1  gate1699(.a(s_165), .O(gate482inter4));
  nand2 gate1700(.a(gate482inter4), .b(gate482inter3), .O(gate482inter5));
  nor2  gate1701(.a(gate482inter5), .b(gate482inter2), .O(gate482inter6));
  inv1  gate1702(.a(G1129), .O(gate482inter7));
  inv1  gate1703(.a(G1225), .O(gate482inter8));
  nand2 gate1704(.a(gate482inter8), .b(gate482inter7), .O(gate482inter9));
  nand2 gate1705(.a(s_165), .b(gate482inter3), .O(gate482inter10));
  nor2  gate1706(.a(gate482inter10), .b(gate482inter9), .O(gate482inter11));
  nor2  gate1707(.a(gate482inter11), .b(gate482inter6), .O(gate482inter12));
  nand2 gate1708(.a(gate482inter12), .b(gate482inter1), .O(G1291));

  xor2  gate1905(.a(G1229), .b(G1228), .O(gate483inter0));
  nand2 gate1906(.a(gate483inter0), .b(s_194), .O(gate483inter1));
  and2  gate1907(.a(G1229), .b(G1228), .O(gate483inter2));
  inv1  gate1908(.a(s_194), .O(gate483inter3));
  inv1  gate1909(.a(s_195), .O(gate483inter4));
  nand2 gate1910(.a(gate483inter4), .b(gate483inter3), .O(gate483inter5));
  nor2  gate1911(.a(gate483inter5), .b(gate483inter2), .O(gate483inter6));
  inv1  gate1912(.a(G1228), .O(gate483inter7));
  inv1  gate1913(.a(G1229), .O(gate483inter8));
  nand2 gate1914(.a(gate483inter8), .b(gate483inter7), .O(gate483inter9));
  nand2 gate1915(.a(s_195), .b(gate483inter3), .O(gate483inter10));
  nor2  gate1916(.a(gate483inter10), .b(gate483inter9), .O(gate483inter11));
  nor2  gate1917(.a(gate483inter11), .b(gate483inter6), .O(gate483inter12));
  nand2 gate1918(.a(gate483inter12), .b(gate483inter1), .O(G1292));
nand2 gate484( .a(G1230), .b(G1231), .O(G1293) );
nand2 gate485( .a(G1232), .b(G1233), .O(G1294) );
nand2 gate486( .a(G1234), .b(G1235), .O(G1295) );
nand2 gate487( .a(G1236), .b(G1237), .O(G1296) );
nand2 gate488( .a(G1238), .b(G1239), .O(G1297) );
nand2 gate489( .a(G1240), .b(G1241), .O(G1298) );

  xor2  gate1681(.a(G1243), .b(G1242), .O(gate490inter0));
  nand2 gate1682(.a(gate490inter0), .b(s_162), .O(gate490inter1));
  and2  gate1683(.a(G1243), .b(G1242), .O(gate490inter2));
  inv1  gate1684(.a(s_162), .O(gate490inter3));
  inv1  gate1685(.a(s_163), .O(gate490inter4));
  nand2 gate1686(.a(gate490inter4), .b(gate490inter3), .O(gate490inter5));
  nor2  gate1687(.a(gate490inter5), .b(gate490inter2), .O(gate490inter6));
  inv1  gate1688(.a(G1242), .O(gate490inter7));
  inv1  gate1689(.a(G1243), .O(gate490inter8));
  nand2 gate1690(.a(gate490inter8), .b(gate490inter7), .O(gate490inter9));
  nand2 gate1691(.a(s_163), .b(gate490inter3), .O(gate490inter10));
  nor2  gate1692(.a(gate490inter10), .b(gate490inter9), .O(gate490inter11));
  nor2  gate1693(.a(gate490inter11), .b(gate490inter6), .O(gate490inter12));
  nand2 gate1694(.a(gate490inter12), .b(gate490inter1), .O(G1299));
nand2 gate491( .a(G1244), .b(G1245), .O(G1300) );
nand2 gate492( .a(G1246), .b(G1247), .O(G1301) );
nand2 gate493( .a(G1248), .b(G1249), .O(G1302) );
nand2 gate494( .a(G1250), .b(G1251), .O(G1303) );
nand2 gate495( .a(G1252), .b(G1253), .O(G1304) );
nand2 gate496( .a(G1254), .b(G1255), .O(G1305) );
nand2 gate497( .a(G1256), .b(G1257), .O(G1306) );
nand2 gate498( .a(G1258), .b(G1259), .O(G1307) );
nand2 gate499( .a(G1260), .b(G1261), .O(G1308) );
nand2 gate500( .a(G1262), .b(G1263), .O(G1309) );

  xor2  gate1569(.a(G1265), .b(G1264), .O(gate501inter0));
  nand2 gate1570(.a(gate501inter0), .b(s_146), .O(gate501inter1));
  and2  gate1571(.a(G1265), .b(G1264), .O(gate501inter2));
  inv1  gate1572(.a(s_146), .O(gate501inter3));
  inv1  gate1573(.a(s_147), .O(gate501inter4));
  nand2 gate1574(.a(gate501inter4), .b(gate501inter3), .O(gate501inter5));
  nor2  gate1575(.a(gate501inter5), .b(gate501inter2), .O(gate501inter6));
  inv1  gate1576(.a(G1264), .O(gate501inter7));
  inv1  gate1577(.a(G1265), .O(gate501inter8));
  nand2 gate1578(.a(gate501inter8), .b(gate501inter7), .O(gate501inter9));
  nand2 gate1579(.a(s_147), .b(gate501inter3), .O(gate501inter10));
  nor2  gate1580(.a(gate501inter10), .b(gate501inter9), .O(gate501inter11));
  nor2  gate1581(.a(gate501inter11), .b(gate501inter6), .O(gate501inter12));
  nand2 gate1582(.a(gate501inter12), .b(gate501inter1), .O(G1310));
nand2 gate502( .a(G1266), .b(G1267), .O(G1311) );
nand2 gate503( .a(G1268), .b(G1269), .O(G1312) );
nand2 gate504( .a(G1270), .b(G1271), .O(G1313) );
nand2 gate505( .a(G1272), .b(G1273), .O(G1314) );
nand2 gate506( .a(G1274), .b(G1275), .O(G1315) );
nand2 gate507( .a(G1276), .b(G1277), .O(G1316) );

  xor2  gate547(.a(G1279), .b(G1278), .O(gate508inter0));
  nand2 gate548(.a(gate508inter0), .b(s_0), .O(gate508inter1));
  and2  gate549(.a(G1279), .b(G1278), .O(gate508inter2));
  inv1  gate550(.a(s_0), .O(gate508inter3));
  inv1  gate551(.a(s_1), .O(gate508inter4));
  nand2 gate552(.a(gate508inter4), .b(gate508inter3), .O(gate508inter5));
  nor2  gate553(.a(gate508inter5), .b(gate508inter2), .O(gate508inter6));
  inv1  gate554(.a(G1278), .O(gate508inter7));
  inv1  gate555(.a(G1279), .O(gate508inter8));
  nand2 gate556(.a(gate508inter8), .b(gate508inter7), .O(gate508inter9));
  nand2 gate557(.a(s_1), .b(gate508inter3), .O(gate508inter10));
  nor2  gate558(.a(gate508inter10), .b(gate508inter9), .O(gate508inter11));
  nor2  gate559(.a(gate508inter11), .b(gate508inter6), .O(gate508inter12));
  nand2 gate560(.a(gate508inter12), .b(gate508inter1), .O(G1317));
nand2 gate509( .a(G1280), .b(G1281), .O(G1318) );
nand2 gate510( .a(G1282), .b(G1283), .O(G1319) );
nand2 gate511( .a(G1284), .b(G1285), .O(G1320) );
nand2 gate512( .a(G1286), .b(G1287), .O(G1321) );
nand2 gate513( .a(G1288), .b(G1289), .O(G1322) );

  xor2  gate1065(.a(G1291), .b(G1290), .O(gate514inter0));
  nand2 gate1066(.a(gate514inter0), .b(s_74), .O(gate514inter1));
  and2  gate1067(.a(G1291), .b(G1290), .O(gate514inter2));
  inv1  gate1068(.a(s_74), .O(gate514inter3));
  inv1  gate1069(.a(s_75), .O(gate514inter4));
  nand2 gate1070(.a(gate514inter4), .b(gate514inter3), .O(gate514inter5));
  nor2  gate1071(.a(gate514inter5), .b(gate514inter2), .O(gate514inter6));
  inv1  gate1072(.a(G1290), .O(gate514inter7));
  inv1  gate1073(.a(G1291), .O(gate514inter8));
  nand2 gate1074(.a(gate514inter8), .b(gate514inter7), .O(gate514inter9));
  nand2 gate1075(.a(s_75), .b(gate514inter3), .O(gate514inter10));
  nor2  gate1076(.a(gate514inter10), .b(gate514inter9), .O(gate514inter11));
  nor2  gate1077(.a(gate514inter11), .b(gate514inter6), .O(gate514inter12));
  nand2 gate1078(.a(gate514inter12), .b(gate514inter1), .O(G1323));
inv1 gate515( .a(G1292), .O(G1324) );
inv1 gate516( .a(G1293), .O(G1325) );
inv1 gate517( .a(G1294), .O(G1326) );
inv1 gate518( .a(G1295), .O(G1327) );
inv1 gate519( .a(G1296), .O(G1328) );
inv1 gate520( .a(G1297), .O(G1329) );
inv1 gate521( .a(G1298), .O(G1330) );
inv1 gate522( .a(G1299), .O(G1331) );
inv1 gate523( .a(G1300), .O(G1332) );
inv1 gate524( .a(G1301), .O(G1333) );
inv1 gate525( .a(G1302), .O(G1334) );
inv1 gate526( .a(G1303), .O(G1335) );
inv1 gate527( .a(G1304), .O(G1336) );
inv1 gate528( .a(G1305), .O(G1337) );
inv1 gate529( .a(G1306), .O(G1338) );
inv1 gate530( .a(G1307), .O(G1339) );
inv1 gate531( .a(G1308), .O(G1340) );
inv1 gate532( .a(G1309), .O(G1341) );
inv1 gate533( .a(G1310), .O(G1342) );
inv1 gate534( .a(G1311), .O(G1343) );
inv1 gate535( .a(G1312), .O(G1344) );
inv1 gate536( .a(G1313), .O(G1345) );
inv1 gate537( .a(G1314), .O(G1346) );
inv1 gate538( .a(G1315), .O(G1347) );
inv1 gate539( .a(G1316), .O(G1348) );
inv1 gate540( .a(G1317), .O(G1349) );
inv1 gate541( .a(G1318), .O(G1350) );
inv1 gate542( .a(G1319), .O(G1351) );
inv1 gate543( .a(G1320), .O(G1352) );
inv1 gate544( .a(G1321), .O(G1353) );
inv1 gate545( .a(G1322), .O(G1354) );
inv1 gate546( .a(G1323), .O(G1355) );

endmodule